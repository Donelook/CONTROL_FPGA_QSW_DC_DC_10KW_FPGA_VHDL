// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Nov 17 2024 15:39:14

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    test,
    start_stop,
    s2_phy,
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    clock_output,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    rgb_g,
    test22,
    rgb_r,
    rgb_b,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output test;
    input start_stop;
    output s2_phy;
    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    output clock_output;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    output rgb_g;
    output test22;
    output rgb_r;
    output rgb_b;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__51921;
    wire N__51920;
    wire N__51919;
    wire N__51910;
    wire N__51909;
    wire N__51908;
    wire N__51901;
    wire N__51900;
    wire N__51899;
    wire N__51892;
    wire N__51891;
    wire N__51890;
    wire N__51883;
    wire N__51882;
    wire N__51881;
    wire N__51874;
    wire N__51873;
    wire N__51872;
    wire N__51865;
    wire N__51864;
    wire N__51863;
    wire N__51856;
    wire N__51855;
    wire N__51854;
    wire N__51847;
    wire N__51846;
    wire N__51845;
    wire N__51838;
    wire N__51837;
    wire N__51836;
    wire N__51829;
    wire N__51828;
    wire N__51827;
    wire N__51820;
    wire N__51819;
    wire N__51818;
    wire N__51811;
    wire N__51810;
    wire N__51809;
    wire N__51802;
    wire N__51801;
    wire N__51800;
    wire N__51793;
    wire N__51792;
    wire N__51791;
    wire N__51784;
    wire N__51783;
    wire N__51782;
    wire N__51765;
    wire N__51764;
    wire N__51763;
    wire N__51762;
    wire N__51759;
    wire N__51756;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51744;
    wire N__51741;
    wire N__51738;
    wire N__51735;
    wire N__51730;
    wire N__51723;
    wire N__51720;
    wire N__51717;
    wire N__51716;
    wire N__51715;
    wire N__51712;
    wire N__51709;
    wire N__51706;
    wire N__51701;
    wire N__51696;
    wire N__51695;
    wire N__51694;
    wire N__51693;
    wire N__51690;
    wire N__51687;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51672;
    wire N__51669;
    wire N__51664;
    wire N__51661;
    wire N__51654;
    wire N__51653;
    wire N__51650;
    wire N__51647;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51624;
    wire N__51623;
    wire N__51622;
    wire N__51621;
    wire N__51620;
    wire N__51619;
    wire N__51618;
    wire N__51617;
    wire N__51616;
    wire N__51613;
    wire N__51612;
    wire N__51605;
    wire N__51604;
    wire N__51603;
    wire N__51602;
    wire N__51601;
    wire N__51600;
    wire N__51597;
    wire N__51596;
    wire N__51595;
    wire N__51594;
    wire N__51593;
    wire N__51592;
    wire N__51589;
    wire N__51582;
    wire N__51581;
    wire N__51580;
    wire N__51579;
    wire N__51574;
    wire N__51571;
    wire N__51560;
    wire N__51559;
    wire N__51558;
    wire N__51557;
    wire N__51556;
    wire N__51555;
    wire N__51554;
    wire N__51553;
    wire N__51552;
    wire N__51551;
    wire N__51548;
    wire N__51543;
    wire N__51536;
    wire N__51531;
    wire N__51526;
    wire N__51523;
    wire N__51522;
    wire N__51521;
    wire N__51520;
    wire N__51519;
    wire N__51518;
    wire N__51517;
    wire N__51516;
    wire N__51515;
    wire N__51508;
    wire N__51505;
    wire N__51504;
    wire N__51503;
    wire N__51502;
    wire N__51501;
    wire N__51494;
    wire N__51491;
    wire N__51488;
    wire N__51483;
    wire N__51480;
    wire N__51469;
    wire N__51464;
    wire N__51461;
    wire N__51460;
    wire N__51457;
    wire N__51450;
    wire N__51447;
    wire N__51446;
    wire N__51445;
    wire N__51444;
    wire N__51443;
    wire N__51442;
    wire N__51441;
    wire N__51440;
    wire N__51439;
    wire N__51438;
    wire N__51437;
    wire N__51436;
    wire N__51435;
    wire N__51434;
    wire N__51433;
    wire N__51432;
    wire N__51431;
    wire N__51430;
    wire N__51427;
    wire N__51422;
    wire N__51419;
    wire N__51416;
    wire N__51415;
    wire N__51410;
    wire N__51395;
    wire N__51392;
    wire N__51391;
    wire N__51390;
    wire N__51389;
    wire N__51388;
    wire N__51387;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51374;
    wire N__51369;
    wire N__51362;
    wire N__51351;
    wire N__51346;
    wire N__51341;
    wire N__51336;
    wire N__51333;
    wire N__51326;
    wire N__51323;
    wire N__51322;
    wire N__51321;
    wire N__51320;
    wire N__51319;
    wire N__51318;
    wire N__51317;
    wire N__51316;
    wire N__51315;
    wire N__51314;
    wire N__51313;
    wire N__51310;
    wire N__51307;
    wire N__51302;
    wire N__51301;
    wire N__51300;
    wire N__51299;
    wire N__51298;
    wire N__51289;
    wire N__51288;
    wire N__51287;
    wire N__51286;
    wire N__51285;
    wire N__51284;
    wire N__51283;
    wire N__51282;
    wire N__51281;
    wire N__51280;
    wire N__51275;
    wire N__51272;
    wire N__51269;
    wire N__51264;
    wire N__51261;
    wire N__51254;
    wire N__51251;
    wire N__51242;
    wire N__51233;
    wire N__51230;
    wire N__51227;
    wire N__51218;
    wire N__51211;
    wire N__51206;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51190;
    wire N__51183;
    wire N__51176;
    wire N__51159;
    wire N__51148;
    wire N__51129;
    wire N__51128;
    wire N__51127;
    wire N__51124;
    wire N__51123;
    wire N__51120;
    wire N__51117;
    wire N__51114;
    wire N__51111;
    wire N__51108;
    wire N__51103;
    wire N__51100;
    wire N__51097;
    wire N__51092;
    wire N__51087;
    wire N__51086;
    wire N__51083;
    wire N__51082;
    wire N__51079;
    wire N__51076;
    wire N__51073;
    wire N__51066;
    wire N__51065;
    wire N__51062;
    wire N__51059;
    wire N__51054;
    wire N__51051;
    wire N__51050;
    wire N__51047;
    wire N__51044;
    wire N__51043;
    wire N__51038;
    wire N__51035;
    wire N__51032;
    wire N__51027;
    wire N__51026;
    wire N__51023;
    wire N__51020;
    wire N__51017;
    wire N__51014;
    wire N__51013;
    wire N__51008;
    wire N__51005;
    wire N__51002;
    wire N__50997;
    wire N__50996;
    wire N__50993;
    wire N__50990;
    wire N__50985;
    wire N__50982;
    wire N__50979;
    wire N__50976;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50966;
    wire N__50963;
    wire N__50960;
    wire N__50957;
    wire N__50954;
    wire N__50951;
    wire N__50946;
    wire N__50943;
    wire N__50940;
    wire N__50937;
    wire N__50934;
    wire N__50931;
    wire N__50928;
    wire N__50925;
    wire N__50922;
    wire N__50919;
    wire N__50916;
    wire N__50915;
    wire N__50914;
    wire N__50913;
    wire N__50912;
    wire N__50911;
    wire N__50910;
    wire N__50909;
    wire N__50908;
    wire N__50907;
    wire N__50906;
    wire N__50905;
    wire N__50904;
    wire N__50903;
    wire N__50902;
    wire N__50901;
    wire N__50900;
    wire N__50899;
    wire N__50898;
    wire N__50897;
    wire N__50896;
    wire N__50895;
    wire N__50894;
    wire N__50893;
    wire N__50892;
    wire N__50891;
    wire N__50890;
    wire N__50889;
    wire N__50888;
    wire N__50887;
    wire N__50886;
    wire N__50885;
    wire N__50884;
    wire N__50883;
    wire N__50882;
    wire N__50881;
    wire N__50880;
    wire N__50879;
    wire N__50878;
    wire N__50877;
    wire N__50876;
    wire N__50875;
    wire N__50874;
    wire N__50873;
    wire N__50872;
    wire N__50871;
    wire N__50870;
    wire N__50869;
    wire N__50868;
    wire N__50867;
    wire N__50866;
    wire N__50865;
    wire N__50864;
    wire N__50863;
    wire N__50862;
    wire N__50861;
    wire N__50860;
    wire N__50859;
    wire N__50858;
    wire N__50857;
    wire N__50856;
    wire N__50855;
    wire N__50854;
    wire N__50853;
    wire N__50852;
    wire N__50851;
    wire N__50850;
    wire N__50849;
    wire N__50848;
    wire N__50847;
    wire N__50846;
    wire N__50845;
    wire N__50844;
    wire N__50843;
    wire N__50842;
    wire N__50841;
    wire N__50840;
    wire N__50839;
    wire N__50838;
    wire N__50837;
    wire N__50836;
    wire N__50835;
    wire N__50834;
    wire N__50833;
    wire N__50832;
    wire N__50831;
    wire N__50830;
    wire N__50829;
    wire N__50828;
    wire N__50827;
    wire N__50826;
    wire N__50825;
    wire N__50824;
    wire N__50823;
    wire N__50822;
    wire N__50821;
    wire N__50820;
    wire N__50819;
    wire N__50818;
    wire N__50817;
    wire N__50816;
    wire N__50815;
    wire N__50814;
    wire N__50813;
    wire N__50812;
    wire N__50811;
    wire N__50810;
    wire N__50809;
    wire N__50808;
    wire N__50807;
    wire N__50806;
    wire N__50805;
    wire N__50804;
    wire N__50803;
    wire N__50802;
    wire N__50801;
    wire N__50800;
    wire N__50799;
    wire N__50798;
    wire N__50797;
    wire N__50796;
    wire N__50795;
    wire N__50794;
    wire N__50793;
    wire N__50792;
    wire N__50791;
    wire N__50790;
    wire N__50789;
    wire N__50788;
    wire N__50787;
    wire N__50786;
    wire N__50785;
    wire N__50784;
    wire N__50783;
    wire N__50782;
    wire N__50781;
    wire N__50780;
    wire N__50779;
    wire N__50778;
    wire N__50777;
    wire N__50776;
    wire N__50775;
    wire N__50774;
    wire N__50773;
    wire N__50772;
    wire N__50771;
    wire N__50770;
    wire N__50769;
    wire N__50768;
    wire N__50767;
    wire N__50766;
    wire N__50765;
    wire N__50764;
    wire N__50763;
    wire N__50762;
    wire N__50761;
    wire N__50760;
    wire N__50759;
    wire N__50758;
    wire N__50757;
    wire N__50756;
    wire N__50753;
    wire N__50752;
    wire N__50751;
    wire N__50750;
    wire N__50421;
    wire N__50418;
    wire N__50417;
    wire N__50416;
    wire N__50415;
    wire N__50412;
    wire N__50407;
    wire N__50404;
    wire N__50401;
    wire N__50398;
    wire N__50395;
    wire N__50394;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50390;
    wire N__50389;
    wire N__50388;
    wire N__50387;
    wire N__50386;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50382;
    wire N__50381;
    wire N__50380;
    wire N__50379;
    wire N__50378;
    wire N__50377;
    wire N__50376;
    wire N__50375;
    wire N__50374;
    wire N__50373;
    wire N__50372;
    wire N__50371;
    wire N__50370;
    wire N__50369;
    wire N__50368;
    wire N__50367;
    wire N__50366;
    wire N__50365;
    wire N__50364;
    wire N__50363;
    wire N__50362;
    wire N__50361;
    wire N__50360;
    wire N__50359;
    wire N__50358;
    wire N__50357;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50352;
    wire N__50351;
    wire N__50350;
    wire N__50349;
    wire N__50348;
    wire N__50347;
    wire N__50346;
    wire N__50345;
    wire N__50344;
    wire N__50343;
    wire N__50342;
    wire N__50341;
    wire N__50340;
    wire N__50339;
    wire N__50338;
    wire N__50337;
    wire N__50336;
    wire N__50335;
    wire N__50334;
    wire N__50333;
    wire N__50332;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50328;
    wire N__50327;
    wire N__50326;
    wire N__50325;
    wire N__50324;
    wire N__50323;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50313;
    wire N__50312;
    wire N__50311;
    wire N__50310;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50296;
    wire N__50295;
    wire N__50294;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50289;
    wire N__50288;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50274;
    wire N__50273;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50269;
    wire N__50268;
    wire N__50267;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50254;
    wire N__50253;
    wire N__50252;
    wire N__50251;
    wire N__50250;
    wire N__50249;
    wire N__50248;
    wire N__50247;
    wire N__50246;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50242;
    wire N__50241;
    wire N__50240;
    wire N__50239;
    wire N__50238;
    wire N__50237;
    wire N__50236;
    wire N__50235;
    wire N__50234;
    wire N__50233;
    wire N__50232;
    wire N__50231;
    wire N__50230;
    wire N__50229;
    wire N__49890;
    wire N__49887;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49879;
    wire N__49876;
    wire N__49873;
    wire N__49872;
    wire N__49871;
    wire N__49870;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49865;
    wire N__49858;
    wire N__49855;
    wire N__49848;
    wire N__49839;
    wire N__49830;
    wire N__49827;
    wire N__49826;
    wire N__49825;
    wire N__49822;
    wire N__49819;
    wire N__49818;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49811;
    wire N__49806;
    wire N__49801;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49794;
    wire N__49793;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49789;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49779;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49770;
    wire N__49769;
    wire N__49766;
    wire N__49763;
    wire N__49756;
    wire N__49753;
    wire N__49746;
    wire N__49737;
    wire N__49730;
    wire N__49727;
    wire N__49726;
    wire N__49723;
    wire N__49722;
    wire N__49719;
    wire N__49718;
    wire N__49715;
    wire N__49714;
    wire N__49711;
    wire N__49710;
    wire N__49707;
    wire N__49706;
    wire N__49703;
    wire N__49702;
    wire N__49699;
    wire N__49698;
    wire N__49695;
    wire N__49692;
    wire N__49691;
    wire N__49688;
    wire N__49687;
    wire N__49684;
    wire N__49683;
    wire N__49680;
    wire N__49679;
    wire N__49678;
    wire N__49675;
    wire N__49674;
    wire N__49671;
    wire N__49670;
    wire N__49667;
    wire N__49666;
    wire N__49661;
    wire N__49660;
    wire N__49659;
    wire N__49658;
    wire N__49649;
    wire N__49646;
    wire N__49643;
    wire N__49640;
    wire N__49625;
    wire N__49608;
    wire N__49591;
    wire N__49576;
    wire N__49573;
    wire N__49568;
    wire N__49565;
    wire N__49562;
    wire N__49559;
    wire N__49554;
    wire N__49545;
    wire N__49542;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49526;
    wire N__49523;
    wire N__49520;
    wire N__49517;
    wire N__49512;
    wire N__49507;
    wire N__49500;
    wire N__49497;
    wire N__49496;
    wire N__49493;
    wire N__49492;
    wire N__49489;
    wire N__49486;
    wire N__49483;
    wire N__49476;
    wire N__49475;
    wire N__49474;
    wire N__49473;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49458;
    wire N__49453;
    wire N__49450;
    wire N__49443;
    wire N__49440;
    wire N__49439;
    wire N__49436;
    wire N__49431;
    wire N__49428;
    wire N__49425;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49419;
    wire N__49416;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49404;
    wire N__49401;
    wire N__49396;
    wire N__49393;
    wire N__49390;
    wire N__49385;
    wire N__49380;
    wire N__49377;
    wire N__49374;
    wire N__49373;
    wire N__49372;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49357;
    wire N__49350;
    wire N__49347;
    wire N__49344;
    wire N__49341;
    wire N__49338;
    wire N__49337;
    wire N__49332;
    wire N__49329;
    wire N__49326;
    wire N__49323;
    wire N__49322;
    wire N__49319;
    wire N__49318;
    wire N__49315;
    wire N__49312;
    wire N__49309;
    wire N__49302;
    wire N__49301;
    wire N__49298;
    wire N__49297;
    wire N__49296;
    wire N__49293;
    wire N__49290;
    wire N__49285;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49271;
    wire N__49268;
    wire N__49263;
    wire N__49260;
    wire N__49257;
    wire N__49254;
    wire N__49251;
    wire N__49250;
    wire N__49249;
    wire N__49248;
    wire N__49247;
    wire N__49246;
    wire N__49245;
    wire N__49244;
    wire N__49243;
    wire N__49242;
    wire N__49241;
    wire N__49240;
    wire N__49239;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49205;
    wire N__49202;
    wire N__49201;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49171;
    wire N__49164;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49154;
    wire N__49153;
    wire N__49150;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49131;
    wire N__49130;
    wire N__49127;
    wire N__49124;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49100;
    wire N__49095;
    wire N__49094;
    wire N__49093;
    wire N__49092;
    wire N__49091;
    wire N__49090;
    wire N__49089;
    wire N__49088;
    wire N__49087;
    wire N__49086;
    wire N__49085;
    wire N__49084;
    wire N__49083;
    wire N__49082;
    wire N__49081;
    wire N__49080;
    wire N__49079;
    wire N__49078;
    wire N__49077;
    wire N__49076;
    wire N__49075;
    wire N__49074;
    wire N__49069;
    wire N__49060;
    wire N__49051;
    wire N__49042;
    wire N__49033;
    wire N__49032;
    wire N__49031;
    wire N__49030;
    wire N__49029;
    wire N__49028;
    wire N__49027;
    wire N__49026;
    wire N__49025;
    wire N__49016;
    wire N__49005;
    wire N__48996;
    wire N__48987;
    wire N__48980;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48968;
    wire N__48963;
    wire N__48962;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48939;
    wire N__48938;
    wire N__48937;
    wire N__48936;
    wire N__48933;
    wire N__48930;
    wire N__48927;
    wire N__48924;
    wire N__48921;
    wire N__48918;
    wire N__48915;
    wire N__48912;
    wire N__48909;
    wire N__48902;
    wire N__48899;
    wire N__48894;
    wire N__48893;
    wire N__48890;
    wire N__48887;
    wire N__48882;
    wire N__48879;
    wire N__48876;
    wire N__48875;
    wire N__48872;
    wire N__48869;
    wire N__48868;
    wire N__48867;
    wire N__48866;
    wire N__48863;
    wire N__48862;
    wire N__48861;
    wire N__48860;
    wire N__48857;
    wire N__48854;
    wire N__48853;
    wire N__48852;
    wire N__48851;
    wire N__48848;
    wire N__48845;
    wire N__48844;
    wire N__48843;
    wire N__48842;
    wire N__48841;
    wire N__48840;
    wire N__48839;
    wire N__48838;
    wire N__48837;
    wire N__48836;
    wire N__48835;
    wire N__48834;
    wire N__48833;
    wire N__48830;
    wire N__48827;
    wire N__48826;
    wire N__48825;
    wire N__48824;
    wire N__48821;
    wire N__48818;
    wire N__48813;
    wire N__48812;
    wire N__48811;
    wire N__48810;
    wire N__48809;
    wire N__48806;
    wire N__48803;
    wire N__48800;
    wire N__48797;
    wire N__48794;
    wire N__48787;
    wire N__48778;
    wire N__48775;
    wire N__48766;
    wire N__48761;
    wire N__48758;
    wire N__48755;
    wire N__48754;
    wire N__48753;
    wire N__48752;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48729;
    wire N__48724;
    wire N__48723;
    wire N__48722;
    wire N__48721;
    wire N__48720;
    wire N__48719;
    wire N__48718;
    wire N__48717;
    wire N__48716;
    wire N__48715;
    wire N__48714;
    wire N__48713;
    wire N__48712;
    wire N__48711;
    wire N__48708;
    wire N__48693;
    wire N__48690;
    wire N__48687;
    wire N__48678;
    wire N__48669;
    wire N__48666;
    wire N__48661;
    wire N__48652;
    wire N__48643;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48616;
    wire N__48597;
    wire N__48594;
    wire N__48593;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48578;
    wire N__48573;
    wire N__48572;
    wire N__48571;
    wire N__48568;
    wire N__48567;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48537;
    wire N__48534;
    wire N__48531;
    wire N__48528;
    wire N__48525;
    wire N__48524;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48511;
    wire N__48508;
    wire N__48501;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48493;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48471;
    wire N__48468;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48455;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48429;
    wire N__48426;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48409;
    wire N__48404;
    wire N__48399;
    wire N__48396;
    wire N__48393;
    wire N__48390;
    wire N__48387;
    wire N__48384;
    wire N__48383;
    wire N__48382;
    wire N__48381;
    wire N__48378;
    wire N__48373;
    wire N__48370;
    wire N__48367;
    wire N__48364;
    wire N__48361;
    wire N__48358;
    wire N__48355;
    wire N__48350;
    wire N__48345;
    wire N__48342;
    wire N__48339;
    wire N__48338;
    wire N__48335;
    wire N__48332;
    wire N__48327;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48312;
    wire N__48309;
    wire N__48308;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48285;
    wire N__48284;
    wire N__48283;
    wire N__48282;
    wire N__48279;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48264;
    wire N__48261;
    wire N__48258;
    wire N__48249;
    wire N__48246;
    wire N__48243;
    wire N__48240;
    wire N__48237;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48225;
    wire N__48222;
    wire N__48219;
    wire N__48216;
    wire N__48215;
    wire N__48214;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48204;
    wire N__48201;
    wire N__48196;
    wire N__48193;
    wire N__48190;
    wire N__48185;
    wire N__48182;
    wire N__48177;
    wire N__48174;
    wire N__48171;
    wire N__48170;
    wire N__48167;
    wire N__48164;
    wire N__48163;
    wire N__48162;
    wire N__48159;
    wire N__48156;
    wire N__48153;
    wire N__48150;
    wire N__48143;
    wire N__48140;
    wire N__48137;
    wire N__48134;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48120;
    wire N__48117;
    wire N__48116;
    wire N__48113;
    wire N__48110;
    wire N__48109;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48093;
    wire N__48090;
    wire N__48089;
    wire N__48088;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48074;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48054;
    wire N__48051;
    wire N__48048;
    wire N__48039;
    wire N__48038;
    wire N__48037;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48027;
    wire N__48024;
    wire N__48019;
    wire N__48016;
    wire N__48013;
    wire N__48010;
    wire N__48003;
    wire N__48000;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47992;
    wire N__47989;
    wire N__47986;
    wire N__47983;
    wire N__47978;
    wire N__47973;
    wire N__47970;
    wire N__47969;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47943;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47889;
    wire N__47888;
    wire N__47887;
    wire N__47884;
    wire N__47881;
    wire N__47878;
    wire N__47875;
    wire N__47872;
    wire N__47869;
    wire N__47866;
    wire N__47861;
    wire N__47856;
    wire N__47855;
    wire N__47854;
    wire N__47853;
    wire N__47850;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47836;
    wire N__47833;
    wire N__47830;
    wire N__47825;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47808;
    wire N__47805;
    wire N__47802;
    wire N__47799;
    wire N__47794;
    wire N__47789;
    wire N__47784;
    wire N__47781;
    wire N__47778;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47739;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47718;
    wire N__47715;
    wire N__47712;
    wire N__47709;
    wire N__47706;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47685;
    wire N__47682;
    wire N__47679;
    wire N__47676;
    wire N__47673;
    wire N__47670;
    wire N__47667;
    wire N__47664;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47652;
    wire N__47649;
    wire N__47646;
    wire N__47643;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47619;
    wire N__47616;
    wire N__47613;
    wire N__47612;
    wire N__47611;
    wire N__47610;
    wire N__47609;
    wire N__47608;
    wire N__47607;
    wire N__47606;
    wire N__47603;
    wire N__47602;
    wire N__47599;
    wire N__47598;
    wire N__47595;
    wire N__47594;
    wire N__47591;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47566;
    wire N__47563;
    wire N__47556;
    wire N__47553;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47535;
    wire N__47532;
    wire N__47529;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47508;
    wire N__47505;
    wire N__47502;
    wire N__47499;
    wire N__47496;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47466;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47427;
    wire N__47424;
    wire N__47421;
    wire N__47418;
    wire N__47415;
    wire N__47412;
    wire N__47409;
    wire N__47406;
    wire N__47403;
    wire N__47400;
    wire N__47397;
    wire N__47394;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47382;
    wire N__47379;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47367;
    wire N__47364;
    wire N__47361;
    wire N__47358;
    wire N__47355;
    wire N__47352;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47238;
    wire N__47235;
    wire N__47232;
    wire N__47229;
    wire N__47226;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47208;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47181;
    wire N__47178;
    wire N__47175;
    wire N__47174;
    wire N__47169;
    wire N__47166;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47162;
    wire N__47161;
    wire N__47160;
    wire N__47159;
    wire N__47158;
    wire N__47157;
    wire N__47156;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47152;
    wire N__47151;
    wire N__47150;
    wire N__47149;
    wire N__47148;
    wire N__47147;
    wire N__47146;
    wire N__47145;
    wire N__47144;
    wire N__47143;
    wire N__47142;
    wire N__47141;
    wire N__47140;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47134;
    wire N__47133;
    wire N__47124;
    wire N__47117;
    wire N__47108;
    wire N__47107;
    wire N__47098;
    wire N__47089;
    wire N__47082;
    wire N__47073;
    wire N__47070;
    wire N__47061;
    wire N__47056;
    wire N__47053;
    wire N__47050;
    wire N__47047;
    wire N__47040;
    wire N__47037;
    wire N__47034;
    wire N__47029;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47000;
    wire N__46995;
    wire N__46994;
    wire N__46991;
    wire N__46988;
    wire N__46985;
    wire N__46980;
    wire N__46977;
    wire N__46976;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46966;
    wire N__46961;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46944;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46936;
    wire N__46933;
    wire N__46932;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46920;
    wire N__46915;
    wire N__46908;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46896;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46882;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46838;
    wire N__46835;
    wire N__46832;
    wire N__46829;
    wire N__46826;
    wire N__46825;
    wire N__46822;
    wire N__46819;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46806;
    wire N__46801;
    wire N__46798;
    wire N__46795;
    wire N__46792;
    wire N__46785;
    wire N__46784;
    wire N__46783;
    wire N__46782;
    wire N__46781;
    wire N__46780;
    wire N__46779;
    wire N__46778;
    wire N__46777;
    wire N__46776;
    wire N__46775;
    wire N__46774;
    wire N__46771;
    wire N__46770;
    wire N__46769;
    wire N__46768;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46764;
    wire N__46763;
    wire N__46762;
    wire N__46761;
    wire N__46758;
    wire N__46755;
    wire N__46752;
    wire N__46751;
    wire N__46750;
    wire N__46749;
    wire N__46748;
    wire N__46745;
    wire N__46742;
    wire N__46729;
    wire N__46726;
    wire N__46721;
    wire N__46720;
    wire N__46719;
    wire N__46714;
    wire N__46713;
    wire N__46712;
    wire N__46711;
    wire N__46708;
    wire N__46705;
    wire N__46702;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46676;
    wire N__46673;
    wire N__46668;
    wire N__46665;
    wire N__46660;
    wire N__46657;
    wire N__46644;
    wire N__46641;
    wire N__46634;
    wire N__46629;
    wire N__46624;
    wire N__46621;
    wire N__46608;
    wire N__46607;
    wire N__46604;
    wire N__46601;
    wire N__46598;
    wire N__46597;
    wire N__46596;
    wire N__46595;
    wire N__46594;
    wire N__46593;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46585;
    wire N__46584;
    wire N__46583;
    wire N__46582;
    wire N__46581;
    wire N__46580;
    wire N__46579;
    wire N__46576;
    wire N__46571;
    wire N__46566;
    wire N__46565;
    wire N__46564;
    wire N__46563;
    wire N__46562;
    wire N__46561;
    wire N__46560;
    wire N__46557;
    wire N__46556;
    wire N__46553;
    wire N__46550;
    wire N__46547;
    wire N__46546;
    wire N__46545;
    wire N__46544;
    wire N__46543;
    wire N__46542;
    wire N__46541;
    wire N__46540;
    wire N__46539;
    wire N__46538;
    wire N__46525;
    wire N__46522;
    wire N__46517;
    wire N__46516;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46490;
    wire N__46487;
    wire N__46482;
    wire N__46469;
    wire N__46462;
    wire N__46459;
    wire N__46452;
    wire N__46449;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46424;
    wire N__46423;
    wire N__46422;
    wire N__46421;
    wire N__46420;
    wire N__46419;
    wire N__46418;
    wire N__46417;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46404;
    wire N__46403;
    wire N__46402;
    wire N__46401;
    wire N__46398;
    wire N__46395;
    wire N__46394;
    wire N__46393;
    wire N__46392;
    wire N__46391;
    wire N__46390;
    wire N__46389;
    wire N__46388;
    wire N__46387;
    wire N__46386;
    wire N__46385;
    wire N__46384;
    wire N__46383;
    wire N__46380;
    wire N__46379;
    wire N__46378;
    wire N__46375;
    wire N__46374;
    wire N__46373;
    wire N__46372;
    wire N__46359;
    wire N__46346;
    wire N__46343;
    wire N__46330;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46320;
    wire N__46315;
    wire N__46312;
    wire N__46309;
    wire N__46306;
    wire N__46299;
    wire N__46294;
    wire N__46289;
    wire N__46284;
    wire N__46279;
    wire N__46276;
    wire N__46263;
    wire N__46256;
    wire N__46253;
    wire N__46248;
    wire N__46245;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46235;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46220;
    wire N__46219;
    wire N__46214;
    wire N__46211;
    wire N__46208;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46182;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46140;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46110;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46020;
    wire N__46017;
    wire N__46014;
    wire N__46011;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45995;
    wire N__45992;
    wire N__45989;
    wire N__45986;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45947;
    wire N__45944;
    wire N__45941;
    wire N__45938;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45923;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45900;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45888;
    wire N__45887;
    wire N__45884;
    wire N__45881;
    wire N__45878;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45864;
    wire N__45861;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45783;
    wire N__45780;
    wire N__45779;
    wire N__45776;
    wire N__45773;
    wire N__45770;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45749;
    wire N__45746;
    wire N__45743;
    wire N__45740;
    wire N__45735;
    wire N__45732;
    wire N__45729;
    wire N__45726;
    wire N__45723;
    wire N__45722;
    wire N__45719;
    wire N__45716;
    wire N__45713;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45692;
    wire N__45689;
    wire N__45686;
    wire N__45683;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45669;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45654;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45617;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45567;
    wire N__45564;
    wire N__45561;
    wire N__45558;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45546;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45540;
    wire N__45537;
    wire N__45532;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45513;
    wire N__45510;
    wire N__45509;
    wire N__45504;
    wire N__45501;
    wire N__45500;
    wire N__45497;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45487;
    wire N__45484;
    wire N__45481;
    wire N__45478;
    wire N__45471;
    wire N__45470;
    wire N__45467;
    wire N__45466;
    wire N__45463;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45443;
    wire N__45440;
    wire N__45435;
    wire N__45434;
    wire N__45429;
    wire N__45426;
    wire N__45425;
    wire N__45424;
    wire N__45419;
    wire N__45416;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45398;
    wire N__45393;
    wire N__45390;
    wire N__45387;
    wire N__45384;
    wire N__45383;
    wire N__45380;
    wire N__45377;
    wire N__45372;
    wire N__45369;
    wire N__45368;
    wire N__45365;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45348;
    wire N__45347;
    wire N__45346;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45321;
    wire N__45312;
    wire N__45311;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45299;
    wire N__45294;
    wire N__45293;
    wire N__45292;
    wire N__45289;
    wire N__45284;
    wire N__45279;
    wire N__45276;
    wire N__45275;
    wire N__45274;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45262;
    wire N__45259;
    wire N__45252;
    wire N__45251;
    wire N__45248;
    wire N__45247;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45235;
    wire N__45232;
    wire N__45227;
    wire N__45222;
    wire N__45221;
    wire N__45216;
    wire N__45213;
    wire N__45210;
    wire N__45209;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45192;
    wire N__45191;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45168;
    wire N__45165;
    wire N__45162;
    wire N__45159;
    wire N__45156;
    wire N__45153;
    wire N__45148;
    wire N__45141;
    wire N__45138;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45110;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45093;
    wire N__45090;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45078;
    wire N__45075;
    wire N__45074;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45057;
    wire N__45056;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45046;
    wire N__45045;
    wire N__45042;
    wire N__45037;
    wire N__45034;
    wire N__45027;
    wire N__45024;
    wire N__45021;
    wire N__45018;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45006;
    wire N__45003;
    wire N__45002;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44985;
    wire N__44984;
    wire N__44983;
    wire N__44982;
    wire N__44979;
    wire N__44976;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44936;
    wire N__44933;
    wire N__44930;
    wire N__44929;
    wire N__44926;
    wire N__44923;
    wire N__44920;
    wire N__44913;
    wire N__44912;
    wire N__44911;
    wire N__44908;
    wire N__44903;
    wire N__44898;
    wire N__44895;
    wire N__44894;
    wire N__44893;
    wire N__44888;
    wire N__44885;
    wire N__44882;
    wire N__44877;
    wire N__44874;
    wire N__44873;
    wire N__44872;
    wire N__44869;
    wire N__44866;
    wire N__44863;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44849;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44825;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44808;
    wire N__44807;
    wire N__44806;
    wire N__44805;
    wire N__44802;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44781;
    wire N__44778;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44768;
    wire N__44767;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44744;
    wire N__44743;
    wire N__44740;
    wire N__44737;
    wire N__44734;
    wire N__44727;
    wire N__44724;
    wire N__44721;
    wire N__44720;
    wire N__44719;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44696;
    wire N__44695;
    wire N__44692;
    wire N__44689;
    wire N__44686;
    wire N__44679;
    wire N__44678;
    wire N__44675;
    wire N__44672;
    wire N__44671;
    wire N__44670;
    wire N__44665;
    wire N__44662;
    wire N__44659;
    wire N__44654;
    wire N__44651;
    wire N__44648;
    wire N__44643;
    wire N__44640;
    wire N__44637;
    wire N__44636;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44619;
    wire N__44618;
    wire N__44617;
    wire N__44614;
    wire N__44613;
    wire N__44610;
    wire N__44607;
    wire N__44604;
    wire N__44601;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44577;
    wire N__44574;
    wire N__44571;
    wire N__44570;
    wire N__44569;
    wire N__44566;
    wire N__44563;
    wire N__44560;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44546;
    wire N__44545;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44529;
    wire N__44526;
    wire N__44523;
    wire N__44522;
    wire N__44521;
    wire N__44518;
    wire N__44515;
    wire N__44512;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44498;
    wire N__44497;
    wire N__44494;
    wire N__44491;
    wire N__44488;
    wire N__44481;
    wire N__44480;
    wire N__44479;
    wire N__44476;
    wire N__44475;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44459;
    wire N__44456;
    wire N__44453;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44441;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44424;
    wire N__44421;
    wire N__44418;
    wire N__44417;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44407;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44393;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44383;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44369;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44352;
    wire N__44349;
    wire N__44346;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44334;
    wire N__44331;
    wire N__44328;
    wire N__44325;
    wire N__44324;
    wire N__44323;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44300;
    wire N__44299;
    wire N__44296;
    wire N__44293;
    wire N__44290;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44276;
    wire N__44275;
    wire N__44272;
    wire N__44269;
    wire N__44266;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44252;
    wire N__44251;
    wire N__44248;
    wire N__44245;
    wire N__44242;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44228;
    wire N__44227;
    wire N__44224;
    wire N__44221;
    wire N__44218;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44204;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44180;
    wire N__44177;
    wire N__44174;
    wire N__44169;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44144;
    wire N__44141;
    wire N__44138;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44127;
    wire N__44126;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44107;
    wire N__44104;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44082;
    wire N__44081;
    wire N__44078;
    wire N__44075;
    wire N__44074;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44058;
    wire N__44057;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44036;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43979;
    wire N__43978;
    wire N__43977;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43932;
    wire N__43929;
    wire N__43926;
    wire N__43923;
    wire N__43922;
    wire N__43919;
    wire N__43916;
    wire N__43915;
    wire N__43912;
    wire N__43909;
    wire N__43906;
    wire N__43905;
    wire N__43902;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43881;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43843;
    wire N__43842;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43824;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43802;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43765;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43734;
    wire N__43731;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43716;
    wire N__43713;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43689;
    wire N__43688;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43676;
    wire N__43673;
    wire N__43670;
    wire N__43669;
    wire N__43664;
    wire N__43663;
    wire N__43660;
    wire N__43659;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43647;
    wire N__43642;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43628;
    wire N__43627;
    wire N__43626;
    wire N__43625;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43611;
    wire N__43608;
    wire N__43607;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43599;
    wire N__43596;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43574;
    wire N__43571;
    wire N__43566;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43542;
    wire N__43539;
    wire N__43536;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43514;
    wire N__43513;
    wire N__43512;
    wire N__43509;
    wire N__43506;
    wire N__43503;
    wire N__43500;
    wire N__43495;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43467;
    wire N__43466;
    wire N__43463;
    wire N__43462;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43443;
    wire N__43440;
    wire N__43437;
    wire N__43434;
    wire N__43425;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43403;
    wire N__43402;
    wire N__43399;
    wire N__43396;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43386;
    wire N__43383;
    wire N__43380;
    wire N__43371;
    wire N__43368;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43349;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43335;
    wire N__43332;
    wire N__43329;
    wire N__43326;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43305;
    wire N__43302;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43286;
    wire N__43283;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43272;
    wire N__43269;
    wire N__43264;
    wire N__43261;
    wire N__43256;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43232;
    wire N__43231;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43190;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43166;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43156;
    wire N__43155;
    wire N__43152;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43131;
    wire N__43128;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43096;
    wire N__43093;
    wire N__43092;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43074;
    wire N__43071;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42987;
    wire N__42984;
    wire N__42981;
    wire N__42978;
    wire N__42977;
    wire N__42974;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42960;
    wire N__42959;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42894;
    wire N__42893;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42836;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42789;
    wire N__42786;
    wire N__42783;
    wire N__42780;
    wire N__42777;
    wire N__42776;
    wire N__42773;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42762;
    wire N__42759;
    wire N__42754;
    wire N__42751;
    wire N__42746;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42719;
    wire N__42718;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42700;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42659;
    wire N__42656;
    wire N__42655;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42623;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42569;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42524;
    wire N__42519;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42489;
    wire N__42486;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42458;
    wire N__42457;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42441;
    wire N__42438;
    wire N__42433;
    wire N__42430;
    wire N__42425;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42411;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42374;
    wire N__42373;
    wire N__42370;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42308;
    wire N__42305;
    wire N__42302;
    wire N__42301;
    wire N__42296;
    wire N__42293;
    wire N__42292;
    wire N__42289;
    wire N__42286;
    wire N__42283;
    wire N__42280;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42226;
    wire N__42223;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42207;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42191;
    wire N__42188;
    wire N__42187;
    wire N__42184;
    wire N__42181;
    wire N__42178;
    wire N__42171;
    wire N__42170;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42152;
    wire N__42149;
    wire N__42146;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42132;
    wire N__42129;
    wire N__42128;
    wire N__42125;
    wire N__42122;
    wire N__42119;
    wire N__42116;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42106;
    wire N__42103;
    wire N__42098;
    wire N__42093;
    wire N__42090;
    wire N__42089;
    wire N__42084;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42074;
    wire N__42069;
    wire N__42068;
    wire N__42065;
    wire N__42064;
    wire N__42061;
    wire N__42058;
    wire N__42053;
    wire N__42050;
    wire N__42049;
    wire N__42046;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42025;
    wire N__42018;
    wire N__42017;
    wire N__42014;
    wire N__42011;
    wire N__42006;
    wire N__42005;
    wire N__42004;
    wire N__42003;
    wire N__42000;
    wire N__41993;
    wire N__41988;
    wire N__41985;
    wire N__41984;
    wire N__41981;
    wire N__41978;
    wire N__41975;
    wire N__41972;
    wire N__41969;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41924;
    wire N__41919;
    wire N__41918;
    wire N__41915;
    wire N__41912;
    wire N__41909;
    wire N__41908;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41892;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41879;
    wire N__41876;
    wire N__41873;
    wire N__41862;
    wire N__41859;
    wire N__41858;
    wire N__41857;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41832;
    wire N__41829;
    wire N__41820;
    wire N__41819;
    wire N__41816;
    wire N__41813;
    wire N__41810;
    wire N__41805;
    wire N__41802;
    wire N__41799;
    wire N__41796;
    wire N__41795;
    wire N__41794;
    wire N__41791;
    wire N__41790;
    wire N__41787;
    wire N__41784;
    wire N__41781;
    wire N__41778;
    wire N__41777;
    wire N__41774;
    wire N__41771;
    wire N__41768;
    wire N__41765;
    wire N__41762;
    wire N__41759;
    wire N__41756;
    wire N__41751;
    wire N__41742;
    wire N__41739;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41720;
    wire N__41717;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41693;
    wire N__41692;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41672;
    wire N__41669;
    wire N__41664;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41627;
    wire N__41624;
    wire N__41621;
    wire N__41618;
    wire N__41615;
    wire N__41614;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41596;
    wire N__41591;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41562;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41552;
    wire N__41549;
    wire N__41544;
    wire N__41541;
    wire N__41540;
    wire N__41537;
    wire N__41534;
    wire N__41531;
    wire N__41526;
    wire N__41523;
    wire N__41520;
    wire N__41517;
    wire N__41516;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41504;
    wire N__41499;
    wire N__41498;
    wire N__41497;
    wire N__41494;
    wire N__41489;
    wire N__41484;
    wire N__41483;
    wire N__41480;
    wire N__41477;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41454;
    wire N__41453;
    wire N__41448;
    wire N__41445;
    wire N__41444;
    wire N__41441;
    wire N__41440;
    wire N__41437;
    wire N__41432;
    wire N__41427;
    wire N__41424;
    wire N__41423;
    wire N__41418;
    wire N__41415;
    wire N__41414;
    wire N__41413;
    wire N__41410;
    wire N__41405;
    wire N__41400;
    wire N__41397;
    wire N__41396;
    wire N__41391;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41376;
    wire N__41373;
    wire N__41372;
    wire N__41371;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41355;
    wire N__41352;
    wire N__41349;
    wire N__41346;
    wire N__41345;
    wire N__41344;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41328;
    wire N__41325;
    wire N__41324;
    wire N__41323;
    wire N__41320;
    wire N__41315;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41300;
    wire N__41295;
    wire N__41292;
    wire N__41291;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41232;
    wire N__41229;
    wire N__41226;
    wire N__41223;
    wire N__41220;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41187;
    wire N__41184;
    wire N__41183;
    wire N__41182;
    wire N__41181;
    wire N__41180;
    wire N__41179;
    wire N__41178;
    wire N__41177;
    wire N__41168;
    wire N__41167;
    wire N__41166;
    wire N__41165;
    wire N__41164;
    wire N__41163;
    wire N__41162;
    wire N__41161;
    wire N__41160;
    wire N__41159;
    wire N__41158;
    wire N__41157;
    wire N__41156;
    wire N__41155;
    wire N__41154;
    wire N__41153;
    wire N__41152;
    wire N__41143;
    wire N__41142;
    wire N__41141;
    wire N__41140;
    wire N__41139;
    wire N__41138;
    wire N__41137;
    wire N__41134;
    wire N__41125;
    wire N__41116;
    wire N__41107;
    wire N__41098;
    wire N__41095;
    wire N__41090;
    wire N__41081;
    wire N__41078;
    wire N__41069;
    wire N__41066;
    wire N__41057;
    wire N__41052;
    wire N__41049;
    wire N__41048;
    wire N__41045;
    wire N__41042;
    wire N__41041;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40983;
    wire N__40980;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40940;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40928;
    wire N__40925;
    wire N__40924;
    wire N__40921;
    wire N__40918;
    wire N__40915;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40895;
    wire N__40890;
    wire N__40887;
    wire N__40886;
    wire N__40881;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40866;
    wire N__40865;
    wire N__40860;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40817;
    wire N__40812;
    wire N__40811;
    wire N__40808;
    wire N__40805;
    wire N__40802;
    wire N__40797;
    wire N__40796;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40760;
    wire N__40755;
    wire N__40752;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40736;
    wire N__40733;
    wire N__40730;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40701;
    wire N__40698;
    wire N__40695;
    wire N__40692;
    wire N__40691;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40679;
    wire N__40674;
    wire N__40671;
    wire N__40670;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40658;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40643;
    wire N__40642;
    wire N__40639;
    wire N__40636;
    wire N__40635;
    wire N__40632;
    wire N__40631;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40615;
    wire N__40610;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40587;
    wire N__40586;
    wire N__40583;
    wire N__40580;
    wire N__40575;
    wire N__40574;
    wire N__40571;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40554;
    wire N__40553;
    wire N__40552;
    wire N__40551;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40518;
    wire N__40517;
    wire N__40516;
    wire N__40513;
    wire N__40512;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40497;
    wire N__40488;
    wire N__40487;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40464;
    wire N__40463;
    wire N__40460;
    wire N__40457;
    wire N__40454;
    wire N__40451;
    wire N__40446;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40410;
    wire N__40407;
    wire N__40406;
    wire N__40405;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40391;
    wire N__40386;
    wire N__40383;
    wire N__40382;
    wire N__40381;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40365;
    wire N__40362;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40337;
    wire N__40334;
    wire N__40331;
    wire N__40328;
    wire N__40323;
    wire N__40322;
    wire N__40319;
    wire N__40316;
    wire N__40315;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40291;
    wire N__40284;
    wire N__40281;
    wire N__40280;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40265;
    wire N__40262;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40238;
    wire N__40237;
    wire N__40232;
    wire N__40229;
    wire N__40226;
    wire N__40221;
    wire N__40218;
    wire N__40217;
    wire N__40216;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40193;
    wire N__40190;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40175;
    wire N__40170;
    wire N__40167;
    wire N__40166;
    wire N__40163;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40148;
    wire N__40143;
    wire N__40140;
    wire N__40139;
    wire N__40136;
    wire N__40133;
    wire N__40132;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40105;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40082;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40067;
    wire N__40062;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40045;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40029;
    wire N__40026;
    wire N__40025;
    wire N__40022;
    wire N__40019;
    wire N__40016;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39993;
    wire N__39990;
    wire N__39989;
    wire N__39988;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39972;
    wire N__39969;
    wire N__39968;
    wire N__39967;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39951;
    wire N__39948;
    wire N__39947;
    wire N__39944;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39929;
    wire N__39924;
    wire N__39921;
    wire N__39920;
    wire N__39917;
    wire N__39914;
    wire N__39913;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39897;
    wire N__39894;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39886;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39870;
    wire N__39867;
    wire N__39866;
    wire N__39865;
    wire N__39860;
    wire N__39857;
    wire N__39854;
    wire N__39849;
    wire N__39846;
    wire N__39843;
    wire N__39842;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39827;
    wire N__39822;
    wire N__39819;
    wire N__39816;
    wire N__39815;
    wire N__39812;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39802;
    wire N__39799;
    wire N__39796;
    wire N__39793;
    wire N__39788;
    wire N__39783;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39772;
    wire N__39769;
    wire N__39766;
    wire N__39763;
    wire N__39760;
    wire N__39753;
    wire N__39750;
    wire N__39749;
    wire N__39748;
    wire N__39743;
    wire N__39740;
    wire N__39737;
    wire N__39732;
    wire N__39729;
    wire N__39728;
    wire N__39727;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39711;
    wire N__39708;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39700;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39684;
    wire N__39681;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39673;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39657;
    wire N__39654;
    wire N__39653;
    wire N__39652;
    wire N__39647;
    wire N__39644;
    wire N__39641;
    wire N__39636;
    wire N__39633;
    wire N__39632;
    wire N__39631;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39615;
    wire N__39612;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39595;
    wire N__39590;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39578;
    wire N__39577;
    wire N__39574;
    wire N__39571;
    wire N__39568;
    wire N__39561;
    wire N__39560;
    wire N__39559;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39543;
    wire N__39540;
    wire N__39539;
    wire N__39536;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39519;
    wire N__39518;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39498;
    wire N__39497;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39485;
    wire N__39480;
    wire N__39477;
    wire N__39476;
    wire N__39473;
    wire N__39472;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39456;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39436;
    wire N__39433;
    wire N__39426;
    wire N__39423;
    wire N__39422;
    wire N__39417;
    wire N__39414;
    wire N__39413;
    wire N__39412;
    wire N__39407;
    wire N__39404;
    wire N__39401;
    wire N__39396;
    wire N__39395;
    wire N__39390;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39354;
    wire N__39353;
    wire N__39352;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39336;
    wire N__39335;
    wire N__39332;
    wire N__39331;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39296;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39264;
    wire N__39261;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39240;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39207;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39195;
    wire N__39192;
    wire N__39189;
    wire N__39188;
    wire N__39185;
    wire N__39182;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39170;
    wire N__39167;
    wire N__39164;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39138;
    wire N__39135;
    wire N__39132;
    wire N__39129;
    wire N__39128;
    wire N__39125;
    wire N__39122;
    wire N__39117;
    wire N__39114;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39102;
    wire N__39101;
    wire N__39098;
    wire N__39095;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39066;
    wire N__39063;
    wire N__39060;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39045;
    wire N__39044;
    wire N__39041;
    wire N__39038;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39024;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39012;
    wire N__39009;
    wire N__39006;
    wire N__39003;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38984;
    wire N__38981;
    wire N__38978;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38963;
    wire N__38960;
    wire N__38957;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38930;
    wire N__38927;
    wire N__38924;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38910;
    wire N__38907;
    wire N__38904;
    wire N__38901;
    wire N__38898;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38886;
    wire N__38883;
    wire N__38880;
    wire N__38877;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38845;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38834;
    wire N__38833;
    wire N__38832;
    wire N__38829;
    wire N__38824;
    wire N__38821;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38811;
    wire N__38808;
    wire N__38803;
    wire N__38800;
    wire N__38787;
    wire N__38786;
    wire N__38783;
    wire N__38780;
    wire N__38775;
    wire N__38774;
    wire N__38773;
    wire N__38772;
    wire N__38771;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38761;
    wire N__38754;
    wire N__38745;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38715;
    wire N__38714;
    wire N__38711;
    wire N__38708;
    wire N__38703;
    wire N__38702;
    wire N__38699;
    wire N__38696;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38678;
    wire N__38675;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38658;
    wire N__38655;
    wire N__38652;
    wire N__38649;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38622;
    wire N__38619;
    wire N__38616;
    wire N__38613;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38592;
    wire N__38589;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38571;
    wire N__38570;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38560;
    wire N__38555;
    wire N__38552;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38531;
    wire N__38530;
    wire N__38529;
    wire N__38528;
    wire N__38527;
    wire N__38526;
    wire N__38525;
    wire N__38524;
    wire N__38523;
    wire N__38522;
    wire N__38521;
    wire N__38520;
    wire N__38519;
    wire N__38518;
    wire N__38517;
    wire N__38510;
    wire N__38501;
    wire N__38500;
    wire N__38499;
    wire N__38498;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38486;
    wire N__38483;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38467;
    wire N__38462;
    wire N__38457;
    wire N__38452;
    wire N__38449;
    wire N__38448;
    wire N__38447;
    wire N__38440;
    wire N__38433;
    wire N__38432;
    wire N__38431;
    wire N__38430;
    wire N__38423;
    wire N__38418;
    wire N__38413;
    wire N__38410;
    wire N__38405;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38387;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38377;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38355;
    wire N__38352;
    wire N__38351;
    wire N__38348;
    wire N__38347;
    wire N__38344;
    wire N__38341;
    wire N__38338;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38296;
    wire N__38291;
    wire N__38288;
    wire N__38283;
    wire N__38280;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38272;
    wire N__38271;
    wire N__38266;
    wire N__38261;
    wire N__38258;
    wire N__38253;
    wire N__38252;
    wire N__38251;
    wire N__38250;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38222;
    wire N__38219;
    wire N__38216;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38186;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38178;
    wire N__38175;
    wire N__38170;
    wire N__38167;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38142;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38111;
    wire N__38108;
    wire N__38105;
    wire N__38102;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38085;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38060;
    wire N__38057;
    wire N__38054;
    wire N__38049;
    wire N__38048;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38031;
    wire N__38030;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37982;
    wire N__37979;
    wire N__37976;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37962;
    wire N__37961;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37944;
    wire N__37941;
    wire N__37940;
    wire N__37937;
    wire N__37934;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37924;
    wire N__37921;
    wire N__37918;
    wire N__37915;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37890;
    wire N__37889;
    wire N__37884;
    wire N__37881;
    wire N__37880;
    wire N__37879;
    wire N__37874;
    wire N__37871;
    wire N__37868;
    wire N__37863;
    wire N__37862;
    wire N__37859;
    wire N__37858;
    wire N__37853;
    wire N__37850;
    wire N__37847;
    wire N__37842;
    wire N__37841;
    wire N__37838;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37826;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37794;
    wire N__37791;
    wire N__37790;
    wire N__37789;
    wire N__37786;
    wire N__37781;
    wire N__37776;
    wire N__37775;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37763;
    wire N__37758;
    wire N__37755;
    wire N__37754;
    wire N__37749;
    wire N__37746;
    wire N__37745;
    wire N__37740;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37701;
    wire N__37698;
    wire N__37697;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37668;
    wire N__37665;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37647;
    wire N__37644;
    wire N__37641;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37580;
    wire N__37579;
    wire N__37576;
    wire N__37575;
    wire N__37574;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37541;
    wire N__37540;
    wire N__37535;
    wire N__37534;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37510;
    wire N__37507;
    wire N__37502;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37463;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37442;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37415;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37403;
    wire N__37402;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37388;
    wire N__37387;
    wire N__37384;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37317;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37274;
    wire N__37271;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37259;
    wire N__37256;
    wire N__37253;
    wire N__37250;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37217;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37205;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37185;
    wire N__37184;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37158;
    wire N__37155;
    wire N__37152;
    wire N__37149;
    wire N__37148;
    wire N__37145;
    wire N__37142;
    wire N__37139;
    wire N__37136;
    wire N__37133;
    wire N__37130;
    wire N__37127;
    wire N__37124;
    wire N__37119;
    wire N__37116;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37022;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__37001;
    wire N__36998;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36971;
    wire N__36968;
    wire N__36965;
    wire N__36962;
    wire N__36959;
    wire N__36956;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36900;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36885;
    wire N__36882;
    wire N__36879;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36869;
    wire N__36866;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36851;
    wire N__36848;
    wire N__36845;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36765;
    wire N__36762;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36725;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36668;
    wire N__36665;
    wire N__36662;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36648;
    wire N__36645;
    wire N__36644;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36629;
    wire N__36626;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36578;
    wire N__36575;
    wire N__36572;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36524;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36494;
    wire N__36491;
    wire N__36488;
    wire N__36485;
    wire N__36482;
    wire N__36479;
    wire N__36476;
    wire N__36473;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36443;
    wire N__36440;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36417;
    wire N__36414;
    wire N__36411;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36395;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36353;
    wire N__36350;
    wire N__36347;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36282;
    wire N__36279;
    wire N__36276;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36240;
    wire N__36237;
    wire N__36234;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36224;
    wire N__36221;
    wire N__36218;
    wire N__36215;
    wire N__36212;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36195;
    wire N__36194;
    wire N__36193;
    wire N__36192;
    wire N__36191;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36164;
    wire N__36161;
    wire N__36160;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36142;
    wire N__36139;
    wire N__36134;
    wire N__36131;
    wire N__36126;
    wire N__36125;
    wire N__36122;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36104;
    wire N__36103;
    wire N__36098;
    wire N__36095;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36067;
    wire N__36062;
    wire N__36059;
    wire N__36058;
    wire N__36053;
    wire N__36050;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36014;
    wire N__36011;
    wire N__36008;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35966;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35948;
    wire N__35945;
    wire N__35940;
    wire N__35937;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35918;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35907;
    wire N__35904;
    wire N__35899;
    wire N__35896;
    wire N__35889;
    wire N__35886;
    wire N__35883;
    wire N__35882;
    wire N__35879;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35865;
    wire N__35864;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35847;
    wire N__35844;
    wire N__35843;
    wire N__35840;
    wire N__35837;
    wire N__35834;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35823;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35805;
    wire N__35802;
    wire N__35801;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35767;
    wire N__35764;
    wire N__35761;
    wire N__35758;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35744;
    wire N__35741;
    wire N__35738;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35718;
    wire N__35715;
    wire N__35712;
    wire N__35709;
    wire N__35706;
    wire N__35697;
    wire N__35694;
    wire N__35691;
    wire N__35690;
    wire N__35687;
    wire N__35684;
    wire N__35683;
    wire N__35678;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35641;
    wire N__35636;
    wire N__35633;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35616;
    wire N__35613;
    wire N__35612;
    wire N__35609;
    wire N__35606;
    wire N__35603;
    wire N__35602;
    wire N__35597;
    wire N__35594;
    wire N__35589;
    wire N__35588;
    wire N__35585;
    wire N__35582;
    wire N__35577;
    wire N__35574;
    wire N__35573;
    wire N__35568;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35556;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35535;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35527;
    wire N__35524;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35509;
    wire N__35508;
    wire N__35505;
    wire N__35500;
    wire N__35497;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35483;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35468;
    wire N__35465;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35438;
    wire N__35435;
    wire N__35432;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35417;
    wire N__35414;
    wire N__35413;
    wire N__35408;
    wire N__35405;
    wire N__35400;
    wire N__35397;
    wire N__35394;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35376;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35358;
    wire N__35355;
    wire N__35352;
    wire N__35351;
    wire N__35348;
    wire N__35345;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35328;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35316;
    wire N__35315;
    wire N__35312;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35284;
    wire N__35277;
    wire N__35274;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35260;
    wire N__35259;
    wire N__35256;
    wire N__35253;
    wire N__35248;
    wire N__35241;
    wire N__35238;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35224;
    wire N__35219;
    wire N__35216;
    wire N__35211;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35199;
    wire N__35196;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35186;
    wire N__35183;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35165;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35138;
    wire N__35135;
    wire N__35132;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35114;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35086;
    wire N__35081;
    wire N__35078;
    wire N__35073;
    wire N__35072;
    wire N__35069;
    wire N__35066;
    wire N__35061;
    wire N__35058;
    wire N__35055;
    wire N__35052;
    wire N__35051;
    wire N__35050;
    wire N__35047;
    wire N__35042;
    wire N__35039;
    wire N__35036;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35019;
    wire N__35016;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34994;
    wire N__34991;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34974;
    wire N__34973;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34963;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34937;
    wire N__34934;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34919;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34907;
    wire N__34906;
    wire N__34905;
    wire N__34904;
    wire N__34901;
    wire N__34896;
    wire N__34893;
    wire N__34890;
    wire N__34887;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34863;
    wire N__34860;
    wire N__34859;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34839;
    wire N__34836;
    wire N__34831;
    wire N__34826;
    wire N__34823;
    wire N__34820;
    wire N__34817;
    wire N__34812;
    wire N__34809;
    wire N__34808;
    wire N__34805;
    wire N__34804;
    wire N__34803;
    wire N__34800;
    wire N__34799;
    wire N__34796;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34780;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34751;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34730;
    wire N__34729;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34723;
    wire N__34722;
    wire N__34721;
    wire N__34720;
    wire N__34719;
    wire N__34718;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34712;
    wire N__34711;
    wire N__34710;
    wire N__34709;
    wire N__34708;
    wire N__34707;
    wire N__34706;
    wire N__34705;
    wire N__34704;
    wire N__34703;
    wire N__34702;
    wire N__34701;
    wire N__34700;
    wire N__34699;
    wire N__34698;
    wire N__34697;
    wire N__34692;
    wire N__34681;
    wire N__34678;
    wire N__34667;
    wire N__34662;
    wire N__34659;
    wire N__34644;
    wire N__34635;
    wire N__34624;
    wire N__34619;
    wire N__34602;
    wire N__34599;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34587;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34341;
    wire N__34340;
    wire N__34339;
    wire N__34338;
    wire N__34337;
    wire N__34336;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34331;
    wire N__34330;
    wire N__34329;
    wire N__34328;
    wire N__34327;
    wire N__34326;
    wire N__34325;
    wire N__34324;
    wire N__34321;
    wire N__34320;
    wire N__34319;
    wire N__34318;
    wire N__34317;
    wire N__34316;
    wire N__34315;
    wire N__34314;
    wire N__34313;
    wire N__34312;
    wire N__34311;
    wire N__34308;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34290;
    wire N__34289;
    wire N__34288;
    wire N__34287;
    wire N__34286;
    wire N__34285;
    wire N__34284;
    wire N__34283;
    wire N__34282;
    wire N__34279;
    wire N__34274;
    wire N__34269;
    wire N__34262;
    wire N__34249;
    wire N__34248;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34244;
    wire N__34243;
    wire N__34242;
    wire N__34241;
    wire N__34240;
    wire N__34235;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34215;
    wire N__34214;
    wire N__34213;
    wire N__34212;
    wire N__34209;
    wire N__34204;
    wire N__34199;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34195;
    wire N__34194;
    wire N__34193;
    wire N__34192;
    wire N__34191;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34183;
    wire N__34182;
    wire N__34181;
    wire N__34180;
    wire N__34179;
    wire N__34178;
    wire N__34177;
    wire N__34176;
    wire N__34169;
    wire N__34166;
    wire N__34161;
    wire N__34154;
    wire N__34145;
    wire N__34134;
    wire N__34133;
    wire N__34132;
    wire N__34131;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34108;
    wire N__34099;
    wire N__34092;
    wire N__34087;
    wire N__34076;
    wire N__34059;
    wire N__34054;
    wire N__34049;
    wire N__34042;
    wire N__34035;
    wire N__34026;
    wire N__34017;
    wire N__33990;
    wire N__33989;
    wire N__33988;
    wire N__33987;
    wire N__33986;
    wire N__33985;
    wire N__33984;
    wire N__33983;
    wire N__33982;
    wire N__33981;
    wire N__33980;
    wire N__33979;
    wire N__33978;
    wire N__33977;
    wire N__33976;
    wire N__33975;
    wire N__33972;
    wire N__33971;
    wire N__33970;
    wire N__33969;
    wire N__33968;
    wire N__33967;
    wire N__33964;
    wire N__33963;
    wire N__33962;
    wire N__33961;
    wire N__33960;
    wire N__33959;
    wire N__33954;
    wire N__33953;
    wire N__33952;
    wire N__33949;
    wire N__33948;
    wire N__33947;
    wire N__33946;
    wire N__33945;
    wire N__33942;
    wire N__33941;
    wire N__33938;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33932;
    wire N__33931;
    wire N__33928;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33920;
    wire N__33917;
    wire N__33916;
    wire N__33915;
    wire N__33912;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33902;
    wire N__33899;
    wire N__33898;
    wire N__33897;
    wire N__33896;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33888;
    wire N__33887;
    wire N__33884;
    wire N__33883;
    wire N__33880;
    wire N__33879;
    wire N__33876;
    wire N__33875;
    wire N__33874;
    wire N__33873;
    wire N__33872;
    wire N__33871;
    wire N__33870;
    wire N__33869;
    wire N__33868;
    wire N__33867;
    wire N__33866;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33855;
    wire N__33846;
    wire N__33843;
    wire N__33838;
    wire N__33835;
    wire N__33828;
    wire N__33825;
    wire N__33814;
    wire N__33805;
    wire N__33794;
    wire N__33793;
    wire N__33790;
    wire N__33789;
    wire N__33788;
    wire N__33787;
    wire N__33786;
    wire N__33785;
    wire N__33784;
    wire N__33783;
    wire N__33782;
    wire N__33781;
    wire N__33774;
    wire N__33769;
    wire N__33766;
    wire N__33765;
    wire N__33764;
    wire N__33763;
    wire N__33762;
    wire N__33759;
    wire N__33758;
    wire N__33755;
    wire N__33754;
    wire N__33751;
    wire N__33750;
    wire N__33747;
    wire N__33746;
    wire N__33739;
    wire N__33722;
    wire N__33719;
    wire N__33718;
    wire N__33715;
    wire N__33714;
    wire N__33711;
    wire N__33710;
    wire N__33707;
    wire N__33706;
    wire N__33703;
    wire N__33702;
    wire N__33699;
    wire N__33698;
    wire N__33695;
    wire N__33694;
    wire N__33691;
    wire N__33690;
    wire N__33687;
    wire N__33686;
    wire N__33683;
    wire N__33682;
    wire N__33679;
    wire N__33678;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33667;
    wire N__33662;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33650;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33629;
    wire N__33628;
    wire N__33627;
    wire N__33626;
    wire N__33623;
    wire N__33622;
    wire N__33621;
    wire N__33618;
    wire N__33611;
    wire N__33606;
    wire N__33601;
    wire N__33594;
    wire N__33593;
    wire N__33590;
    wire N__33589;
    wire N__33586;
    wire N__33585;
    wire N__33582;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33560;
    wire N__33555;
    wire N__33538;
    wire N__33521;
    wire N__33504;
    wire N__33503;
    wire N__33502;
    wire N__33499;
    wire N__33498;
    wire N__33495;
    wire N__33494;
    wire N__33491;
    wire N__33490;
    wire N__33489;
    wire N__33488;
    wire N__33485;
    wire N__33484;
    wire N__33479;
    wire N__33474;
    wire N__33461;
    wire N__33444;
    wire N__33435;
    wire N__33418;
    wire N__33405;
    wire N__33400;
    wire N__33387;
    wire N__33378;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33331;
    wire N__33328;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33284;
    wire N__33281;
    wire N__33278;
    wire N__33273;
    wire N__33270;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33017;
    wire N__33014;
    wire N__33011;
    wire N__33006;
    wire N__33003;
    wire N__33002;
    wire N__33001;
    wire N__32998;
    wire N__32993;
    wire N__32988;
    wire N__32985;
    wire N__32982;
    wire N__32981;
    wire N__32978;
    wire N__32975;
    wire N__32972;
    wire N__32969;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32924;
    wire N__32921;
    wire N__32918;
    wire N__32917;
    wire N__32914;
    wire N__32911;
    wire N__32908;
    wire N__32901;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32856;
    wire N__32853;
    wire N__32850;
    wire N__32847;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32837;
    wire N__32834;
    wire N__32831;
    wire N__32826;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32816;
    wire N__32813;
    wire N__32812;
    wire N__32809;
    wire N__32806;
    wire N__32803;
    wire N__32800;
    wire N__32795;
    wire N__32792;
    wire N__32789;
    wire N__32784;
    wire N__32781;
    wire N__32780;
    wire N__32775;
    wire N__32772;
    wire N__32769;
    wire N__32768;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32753;
    wire N__32748;
    wire N__32747;
    wire N__32746;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32717;
    wire N__32714;
    wire N__32711;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32693;
    wire N__32692;
    wire N__32691;
    wire N__32690;
    wire N__32689;
    wire N__32688;
    wire N__32687;
    wire N__32686;
    wire N__32685;
    wire N__32684;
    wire N__32683;
    wire N__32682;
    wire N__32681;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32677;
    wire N__32676;
    wire N__32675;
    wire N__32674;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32670;
    wire N__32669;
    wire N__32668;
    wire N__32667;
    wire N__32666;
    wire N__32665;
    wire N__32664;
    wire N__32663;
    wire N__32662;
    wire N__32661;
    wire N__32660;
    wire N__32659;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32655;
    wire N__32654;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32645;
    wire N__32644;
    wire N__32641;
    wire N__32640;
    wire N__32639;
    wire N__32634;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32622;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32604;
    wire N__32603;
    wire N__32596;
    wire N__32589;
    wire N__32578;
    wire N__32571;
    wire N__32566;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32561;
    wire N__32558;
    wire N__32551;
    wire N__32542;
    wire N__32539;
    wire N__32534;
    wire N__32521;
    wire N__32510;
    wire N__32507;
    wire N__32504;
    wire N__32501;
    wire N__32498;
    wire N__32495;
    wire N__32494;
    wire N__32493;
    wire N__32492;
    wire N__32491;
    wire N__32490;
    wire N__32489;
    wire N__32488;
    wire N__32487;
    wire N__32486;
    wire N__32485;
    wire N__32478;
    wire N__32473;
    wire N__32470;
    wire N__32465;
    wire N__32460;
    wire N__32447;
    wire N__32442;
    wire N__32437;
    wire N__32434;
    wire N__32433;
    wire N__32432;
    wire N__32427;
    wire N__32422;
    wire N__32419;
    wire N__32416;
    wire N__32411;
    wire N__32400;
    wire N__32391;
    wire N__32390;
    wire N__32389;
    wire N__32388;
    wire N__32387;
    wire N__32386;
    wire N__32385;
    wire N__32384;
    wire N__32383;
    wire N__32382;
    wire N__32377;
    wire N__32374;
    wire N__32365;
    wire N__32364;
    wire N__32359;
    wire N__32356;
    wire N__32353;
    wire N__32346;
    wire N__32335;
    wire N__32330;
    wire N__32325;
    wire N__32314;
    wire N__32303;
    wire N__32294;
    wire N__32287;
    wire N__32284;
    wire N__32277;
    wire N__32272;
    wire N__32253;
    wire N__32252;
    wire N__32249;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32232;
    wire N__32231;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32214;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32200;
    wire N__32195;
    wire N__32192;
    wire N__32187;
    wire N__32186;
    wire N__32181;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32173;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32150;
    wire N__32149;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32145;
    wire N__32144;
    wire N__32143;
    wire N__32142;
    wire N__32141;
    wire N__32140;
    wire N__32139;
    wire N__32136;
    wire N__32135;
    wire N__32134;
    wire N__32133;
    wire N__32122;
    wire N__32119;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32115;
    wire N__32114;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32110;
    wire N__32109;
    wire N__32108;
    wire N__32107;
    wire N__32106;
    wire N__32105;
    wire N__32104;
    wire N__32097;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32075;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32065;
    wire N__32062;
    wire N__32059;
    wire N__32056;
    wire N__32053;
    wire N__32044;
    wire N__32035;
    wire N__32028;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31981;
    wire N__31970;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31946;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31910;
    wire N__31909;
    wire N__31906;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31894;
    wire N__31891;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31865;
    wire N__31862;
    wire N__31861;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31842;
    wire N__31839;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31811;
    wire N__31810;
    wire N__31807;
    wire N__31802;
    wire N__31801;
    wire N__31796;
    wire N__31793;
    wire N__31790;
    wire N__31787;
    wire N__31782;
    wire N__31779;
    wire N__31778;
    wire N__31775;
    wire N__31772;
    wire N__31767;
    wire N__31766;
    wire N__31763;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31746;
    wire N__31745;
    wire N__31742;
    wire N__31741;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31720;
    wire N__31715;
    wire N__31712;
    wire N__31709;
    wire N__31704;
    wire N__31703;
    wire N__31702;
    wire N__31701;
    wire N__31700;
    wire N__31699;
    wire N__31698;
    wire N__31697;
    wire N__31696;
    wire N__31695;
    wire N__31694;
    wire N__31693;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31661;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31646;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31625;
    wire N__31620;
    wire N__31617;
    wire N__31616;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31604;
    wire N__31599;
    wire N__31598;
    wire N__31595;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31585;
    wire N__31578;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31535;
    wire N__31530;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31515;
    wire N__31512;
    wire N__31511;
    wire N__31506;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31472;
    wire N__31471;
    wire N__31470;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31455;
    wire N__31448;
    wire N__31443;
    wire N__31440;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31428;
    wire N__31427;
    wire N__31422;
    wire N__31419;
    wire N__31418;
    wire N__31415;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31403;
    wire N__31402;
    wire N__31401;
    wire N__31398;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31365;
    wire N__31362;
    wire N__31359;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31347;
    wire N__31346;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31310;
    wire N__31307;
    wire N__31304;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31289;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31269;
    wire N__31268;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31223;
    wire N__31222;
    wire N__31221;
    wire N__31214;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31199;
    wire N__31196;
    wire N__31193;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30897;
    wire N__30896;
    wire N__30893;
    wire N__30890;
    wire N__30889;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30788;
    wire N__30785;
    wire N__30782;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30686;
    wire N__30683;
    wire N__30680;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30606;
    wire N__30605;
    wire N__30602;
    wire N__30599;
    wire N__30598;
    wire N__30593;
    wire N__30590;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30572;
    wire N__30569;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30420;
    wire N__30417;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30407;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30371;
    wire N__30368;
    wire N__30365;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30347;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30329;
    wire N__30326;
    wire N__30323;
    wire N__30322;
    wire N__30317;
    wire N__30314;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30287;
    wire N__30284;
    wire N__30283;
    wire N__30280;
    wire N__30275;
    wire N__30272;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30249;
    wire N__30248;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30222;
    wire N__30219;
    wire N__30218;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30182;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30167;
    wire N__30164;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30134;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30116;
    wire N__30113;
    wire N__30110;
    wire N__30105;
    wire N__30102;
    wire N__30101;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30065;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30044;
    wire N__30041;
    wire N__30038;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30016;
    wire N__30013;
    wire N__30008;
    wire N__30005;
    wire N__30002;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29990;
    wire N__29989;
    wire N__29988;
    wire N__29987;
    wire N__29986;
    wire N__29985;
    wire N__29984;
    wire N__29983;
    wire N__29982;
    wire N__29981;
    wire N__29980;
    wire N__29971;
    wire N__29962;
    wire N__29961;
    wire N__29960;
    wire N__29959;
    wire N__29958;
    wire N__29957;
    wire N__29956;
    wire N__29955;
    wire N__29954;
    wire N__29953;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29949;
    wire N__29948;
    wire N__29947;
    wire N__29946;
    wire N__29945;
    wire N__29944;
    wire N__29943;
    wire N__29934;
    wire N__29929;
    wire N__29922;
    wire N__29913;
    wire N__29912;
    wire N__29909;
    wire N__29900;
    wire N__29893;
    wire N__29884;
    wire N__29881;
    wire N__29874;
    wire N__29871;
    wire N__29858;
    wire N__29855;
    wire N__29850;
    wire N__29847;
    wire N__29846;
    wire N__29843;
    wire N__29838;
    wire N__29837;
    wire N__29834;
    wire N__29831;
    wire N__29828;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29809;
    wire N__29808;
    wire N__29803;
    wire N__29800;
    wire N__29797;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29768;
    wire N__29765;
    wire N__29762;
    wire N__29761;
    wire N__29760;
    wire N__29757;
    wire N__29750;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29702;
    wire N__29701;
    wire N__29698;
    wire N__29693;
    wire N__29688;
    wire N__29685;
    wire N__29684;
    wire N__29681;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29657;
    wire N__29654;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29642;
    wire N__29639;
    wire N__29634;
    wire N__29631;
    wire N__29630;
    wire N__29627;
    wire N__29624;
    wire N__29621;
    wire N__29616;
    wire N__29613;
    wire N__29612;
    wire N__29609;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29594;
    wire N__29589;
    wire N__29586;
    wire N__29585;
    wire N__29582;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29567;
    wire N__29562;
    wire N__29559;
    wire N__29558;
    wire N__29557;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29541;
    wire N__29538;
    wire N__29537;
    wire N__29534;
    wire N__29529;
    wire N__29528;
    wire N__29525;
    wire N__29522;
    wire N__29519;
    wire N__29514;
    wire N__29511;
    wire N__29510;
    wire N__29509;
    wire N__29504;
    wire N__29501;
    wire N__29498;
    wire N__29493;
    wire N__29490;
    wire N__29489;
    wire N__29486;
    wire N__29485;
    wire N__29480;
    wire N__29477;
    wire N__29474;
    wire N__29469;
    wire N__29466;
    wire N__29465;
    wire N__29464;
    wire N__29459;
    wire N__29456;
    wire N__29453;
    wire N__29448;
    wire N__29445;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29423;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29399;
    wire N__29396;
    wire N__29391;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29381;
    wire N__29376;
    wire N__29373;
    wire N__29372;
    wire N__29371;
    wire N__29366;
    wire N__29363;
    wire N__29360;
    wire N__29355;
    wire N__29352;
    wire N__29351;
    wire N__29346;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29324;
    wire N__29319;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29304;
    wire N__29301;
    wire N__29300;
    wire N__29295;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29273;
    wire N__29270;
    wire N__29267;
    wire N__29264;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29243;
    wire N__29238;
    wire N__29235;
    wire N__29232;
    wire N__29231;
    wire N__29228;
    wire N__29225;
    wire N__29222;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29199;
    wire N__29196;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29181;
    wire N__29178;
    wire N__29177;
    wire N__29174;
    wire N__29171;
    wire N__29168;
    wire N__29163;
    wire N__29160;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29145;
    wire N__29142;
    wire N__29139;
    wire N__29138;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29124;
    wire N__29121;
    wire N__29120;
    wire N__29117;
    wire N__29114;
    wire N__29109;
    wire N__29106;
    wire N__29103;
    wire N__29102;
    wire N__29099;
    wire N__29096;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29074;
    wire N__29073;
    wire N__29072;
    wire N__29069;
    wire N__29066;
    wire N__29059;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29036;
    wire N__29031;
    wire N__29028;
    wire N__29025;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29012;
    wire N__29009;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28992;
    wire N__28989;
    wire N__28988;
    wire N__28985;
    wire N__28982;
    wire N__28977;
    wire N__28974;
    wire N__28973;
    wire N__28970;
    wire N__28967;
    wire N__28964;
    wire N__28959;
    wire N__28956;
    wire N__28955;
    wire N__28952;
    wire N__28949;
    wire N__28944;
    wire N__28941;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28926;
    wire N__28923;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28908;
    wire N__28905;
    wire N__28904;
    wire N__28901;
    wire N__28898;
    wire N__28895;
    wire N__28890;
    wire N__28887;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28877;
    wire N__28874;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28851;
    wire N__28848;
    wire N__28847;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28806;
    wire N__28803;
    wire N__28802;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28779;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28764;
    wire N__28761;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28745;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28694;
    wire N__28691;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28674;
    wire N__28673;
    wire N__28672;
    wire N__28669;
    wire N__28664;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28628;
    wire N__28625;
    wire N__28624;
    wire N__28621;
    wire N__28616;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28581;
    wire N__28578;
    wire N__28575;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28493;
    wire N__28488;
    wire N__28487;
    wire N__28484;
    wire N__28481;
    wire N__28478;
    wire N__28473;
    wire N__28470;
    wire N__28469;
    wire N__28464;
    wire N__28463;
    wire N__28460;
    wire N__28457;
    wire N__28454;
    wire N__28449;
    wire N__28446;
    wire N__28445;
    wire N__28440;
    wire N__28439;
    wire N__28436;
    wire N__28433;
    wire N__28430;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28418;
    wire N__28417;
    wire N__28414;
    wire N__28411;
    wire N__28408;
    wire N__28403;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28349;
    wire N__28346;
    wire N__28341;
    wire N__28340;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28326;
    wire N__28323;
    wire N__28322;
    wire N__28317;
    wire N__28316;
    wire N__28313;
    wire N__28310;
    wire N__28307;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28295;
    wire N__28290;
    wire N__28289;
    wire N__28286;
    wire N__28283;
    wire N__28280;
    wire N__28275;
    wire N__28272;
    wire N__28271;
    wire N__28266;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28256;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28244;
    wire N__28241;
    wire N__28236;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28221;
    wire N__28218;
    wire N__28217;
    wire N__28212;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28197;
    wire N__28194;
    wire N__28193;
    wire N__28192;
    wire N__28187;
    wire N__28184;
    wire N__28181;
    wire N__28176;
    wire N__28173;
    wire N__28172;
    wire N__28169;
    wire N__28166;
    wire N__28163;
    wire N__28158;
    wire N__28155;
    wire N__28154;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28137;
    wire N__28136;
    wire N__28133;
    wire N__28130;
    wire N__28127;
    wire N__28122;
    wire N__28119;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28104;
    wire N__28101;
    wire N__28100;
    wire N__28097;
    wire N__28094;
    wire N__28091;
    wire N__28086;
    wire N__28083;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28068;
    wire N__28065;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28053;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28043;
    wire N__28038;
    wire N__28035;
    wire N__28034;
    wire N__28029;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28019;
    wire N__28014;
    wire N__28011;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27996;
    wire N__27993;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27981;
    wire N__27978;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27968;
    wire N__27963;
    wire N__27960;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27945;
    wire N__27942;
    wire N__27941;
    wire N__27938;
    wire N__27935;
    wire N__27932;
    wire N__27927;
    wire N__27924;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27909;
    wire N__27906;
    wire N__27905;
    wire N__27902;
    wire N__27899;
    wire N__27896;
    wire N__27891;
    wire N__27888;
    wire N__27887;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27873;
    wire N__27870;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27860;
    wire N__27855;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27732;
    wire N__27729;
    wire N__27726;
    wire N__27725;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27707;
    wire N__27704;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27398;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27365;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27321;
    wire N__27318;
    wire N__27317;
    wire N__27316;
    wire N__27313;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27298;
    wire N__27295;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27279;
    wire N__27278;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26609;
    wire N__26606;
    wire N__26605;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26574;
    wire N__26571;
    wire N__26570;
    wire N__26565;
    wire N__26562;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26550;
    wire N__26547;
    wire N__26546;
    wire N__26543;
    wire N__26540;
    wire N__26537;
    wire N__26534;
    wire N__26531;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26484;
    wire N__26481;
    wire N__26478;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26418;
    wire N__26417;
    wire N__26412;
    wire N__26409;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26397;
    wire N__26394;
    wire N__26393;
    wire N__26390;
    wire N__26389;
    wire N__26386;
    wire N__26383;
    wire N__26380;
    wire N__26373;
    wire N__26370;
    wire N__26369;
    wire N__26368;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26336;
    wire N__26331;
    wire N__26328;
    wire N__26327;
    wire N__26322;
    wire N__26319;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26307;
    wire N__26304;
    wire N__26303;
    wire N__26298;
    wire N__26295;
    wire N__26294;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26274;
    wire N__26271;
    wire N__26268;
    wire N__26267;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26246;
    wire N__26245;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26223;
    wire N__26222;
    wire N__26219;
    wire N__26216;
    wire N__26215;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26203;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26187;
    wire N__26184;
    wire N__26183;
    wire N__26180;
    wire N__26177;
    wire N__26172;
    wire N__26169;
    wire N__26168;
    wire N__26167;
    wire N__26164;
    wire N__26159;
    wire N__26158;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26144;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26132;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26120;
    wire N__26117;
    wire N__26114;
    wire N__26109;
    wire N__26108;
    wire N__26107;
    wire N__26104;
    wire N__26099;
    wire N__26096;
    wire N__26095;
    wire N__26092;
    wire N__26089;
    wire N__26086;
    wire N__26083;
    wire N__26078;
    wire N__26073;
    wire N__26070;
    wire N__26069;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26050;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26036;
    wire N__26031;
    wire N__26028;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26020;
    wire N__26015;
    wire N__26012;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25995;
    wire N__25992;
    wire N__25991;
    wire N__25988;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25971;
    wire N__25970;
    wire N__25967;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25947;
    wire N__25944;
    wire N__25937;
    wire N__25934;
    wire N__25929;
    wire N__25928;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25916;
    wire N__25911;
    wire N__25908;
    wire N__25907;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25896;
    wire N__25891;
    wire N__25888;
    wire N__25885;
    wire N__25882;
    wire N__25877;
    wire N__25872;
    wire N__25871;
    wire N__25868;
    wire N__25867;
    wire N__25864;
    wire N__25861;
    wire N__25858;
    wire N__25851;
    wire N__25850;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25838;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25791;
    wire N__25788;
    wire N__25787;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25764;
    wire N__25763;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25748;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25731;
    wire N__25728;
    wire N__25725;
    wire N__25724;
    wire N__25721;
    wire N__25718;
    wire N__25715;
    wire N__25714;
    wire N__25709;
    wire N__25706;
    wire N__25703;
    wire N__25698;
    wire N__25697;
    wire N__25696;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25556;
    wire N__25553;
    wire N__25548;
    wire N__25545;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25379;
    wire N__25374;
    wire N__25371;
    wire N__25370;
    wire N__25365;
    wire N__25362;
    wire N__25361;
    wire N__25358;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25350;
    wire N__25347;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25327;
    wire N__25320;
    wire N__25317;
    wire N__25316;
    wire N__25313;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25296;
    wire N__25293;
    wire N__25292;
    wire N__25287;
    wire N__25284;
    wire N__25283;
    wire N__25280;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25265;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25250;
    wire N__25245;
    wire N__25244;
    wire N__25241;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25231;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25213;
    wire N__25208;
    wire N__25203;
    wire N__25200;
    wire N__25199;
    wire N__25196;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25186;
    wire N__25179;
    wire N__25178;
    wire N__25175;
    wire N__25174;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25134;
    wire N__25131;
    wire N__25130;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25119;
    wire N__25114;
    wire N__25111;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25092;
    wire N__25091;
    wire N__25088;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25073;
    wire N__25068;
    wire N__25065;
    wire N__25064;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25041;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25033;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25001;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24974;
    wire N__24969;
    wire N__24966;
    wire N__24965;
    wire N__24964;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24933;
    wire N__24932;
    wire N__24929;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24900;
    wire N__24893;
    wire N__24890;
    wire N__24885;
    wire N__24882;
    wire N__24881;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24864;
    wire N__24863;
    wire N__24862;
    wire N__24859;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24835;
    wire N__24830;
    wire N__24825;
    wire N__24824;
    wire N__24821;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24804;
    wire N__24801;
    wire N__24800;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24769;
    wire N__24766;
    wire N__24759;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24737;
    wire N__24732;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24721;
    wire N__24716;
    wire N__24713;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24696;
    wire N__24693;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24685;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24669;
    wire N__24664;
    wire N__24661;
    wire N__24654;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24636;
    wire N__24635;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24617;
    wire N__24612;
    wire N__24611;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24600;
    wire N__24597;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24578;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24368;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24327;
    wire N__24324;
    wire N__24321;
    wire N__24320;
    wire N__24319;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24303;
    wire N__24300;
    wire N__24299;
    wire N__24298;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24275;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24258;
    wire N__24255;
    wire N__24254;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24239;
    wire N__24234;
    wire N__24231;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24219;
    wire N__24216;
    wire N__24215;
    wire N__24214;
    wire N__24213;
    wire N__24212;
    wire N__24211;
    wire N__24210;
    wire N__24209;
    wire N__24208;
    wire N__24207;
    wire N__24206;
    wire N__24205;
    wire N__24204;
    wire N__24203;
    wire N__24194;
    wire N__24185;
    wire N__24180;
    wire N__24179;
    wire N__24178;
    wire N__24177;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24172;
    wire N__24171;
    wire N__24170;
    wire N__24169;
    wire N__24168;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24164;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24137;
    wire N__24128;
    wire N__24119;
    wire N__24110;
    wire N__24107;
    wire N__24096;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24078;
    wire N__24075;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24063;
    wire N__24062;
    wire N__24061;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24026;
    wire N__24021;
    wire N__24018;
    wire N__24017;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24000;
    wire N__23997;
    wire N__23994;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23976;
    wire N__23973;
    wire N__23970;
    wire N__23969;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23921;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23897;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23873;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23849;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23832;
    wire N__23829;
    wire N__23826;
    wire N__23825;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23801;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23777;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23753;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23743;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23729;
    wire N__23728;
    wire N__23725;
    wire N__23722;
    wire N__23719;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23695;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23681;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23657;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23633;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23577;
    wire N__23574;
    wire N__23573;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23549;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23532;
    wire N__23529;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23513;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23442;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23284;
    wire N__23283;
    wire N__23282;
    wire N__23281;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23261;
    wire N__23256;
    wire N__23251;
    wire N__23246;
    wire N__23243;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23090;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23076;
    wire N__23073;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23054;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23038;
    wire N__23037;
    wire N__23036;
    wire N__23035;
    wire N__23034;
    wire N__23033;
    wire N__23032;
    wire N__23031;
    wire N__23028;
    wire N__23023;
    wire N__23020;
    wire N__23011;
    wire N__23006;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22896;
    wire N__22893;
    wire N__22892;
    wire N__22889;
    wire N__22886;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22838;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22802;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22779;
    wire N__22776;
    wire N__22775;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22721;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22709;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22688;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22634;
    wire N__22631;
    wire N__22628;
    wire N__22623;
    wire N__22620;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22607;
    wire N__22602;
    wire N__22599;
    wire N__22598;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22570;
    wire N__22565;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22545;
    wire N__22542;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22490;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22448;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22380;
    wire N__22377;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22365;
    wire N__22362;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22332;
    wire N__22329;
    wire N__22328;
    wire N__22327;
    wire N__22326;
    wire N__22323;
    wire N__22316;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22256;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22238;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22201;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22181;
    wire N__22178;
    wire N__22175;
    wire N__22170;
    wire N__22167;
    wire N__22166;
    wire N__22165;
    wire N__22164;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22112;
    wire N__22109;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22092;
    wire N__22089;
    wire N__22088;
    wire N__22085;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22068;
    wire N__22065;
    wire N__22064;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22044;
    wire N__22041;
    wire N__22040;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22013;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21963;
    wire N__21960;
    wire N__21957;
    wire N__21956;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21936;
    wire N__21935;
    wire N__21934;
    wire N__21933;
    wire N__21932;
    wire N__21931;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21918;
    wire N__21913;
    wire N__21904;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21827;
    wire N__21824;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21807;
    wire N__21804;
    wire N__21803;
    wire N__21800;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21783;
    wire N__21780;
    wire N__21779;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21705;
    wire N__21704;
    wire N__21703;
    wire N__21702;
    wire N__21701;
    wire N__21700;
    wire N__21699;
    wire N__21698;
    wire N__21697;
    wire N__21694;
    wire N__21677;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21662;
    wire N__21657;
    wire N__21656;
    wire N__21655;
    wire N__21654;
    wire N__21653;
    wire N__21652;
    wire N__21651;
    wire N__21650;
    wire N__21649;
    wire N__21646;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21612;
    wire N__21611;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21600;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21596;
    wire N__21595;
    wire N__21594;
    wire N__21593;
    wire N__21592;
    wire N__21591;
    wire N__21590;
    wire N__21589;
    wire N__21588;
    wire N__21583;
    wire N__21582;
    wire N__21579;
    wire N__21578;
    wire N__21575;
    wire N__21574;
    wire N__21571;
    wire N__21570;
    wire N__21567;
    wire N__21566;
    wire N__21565;
    wire N__21564;
    wire N__21563;
    wire N__21562;
    wire N__21559;
    wire N__21558;
    wire N__21541;
    wire N__21526;
    wire N__21523;
    wire N__21506;
    wire N__21501;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21477;
    wire N__21472;
    wire N__21463;
    wire N__21460;
    wire N__21455;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21254;
    wire N__21253;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21239;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21119;
    wire N__21114;
    wire N__21113;
    wire N__21112;
    wire N__21111;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21103;
    wire N__21100;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21095;
    wire N__21092;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21077;
    wire N__21070;
    wire N__21061;
    wire N__21054;
    wire N__21045;
    wire N__21044;
    wire N__21041;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21017;
    wire N__21016;
    wire N__21015;
    wire N__21014;
    wire N__21011;
    wire N__21010;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20994;
    wire N__20993;
    wire N__20988;
    wire N__20985;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20837;
    wire N__20836;
    wire N__20833;
    wire N__20828;
    wire N__20823;
    wire N__20822;
    wire N__20819;
    wire N__20816;
    wire N__20813;
    wire N__20810;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20783;
    wire N__20780;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20763;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20670;
    wire N__20667;
    wire N__20666;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20643;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20622;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20577;
    wire N__20574;
    wire N__20573;
    wire N__20570;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20546;
    wire N__20543;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20512;
    wire N__20509;
    wire N__20506;
    wire N__20503;
    wire N__20498;
    wire N__20495;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20297;
    wire N__20294;
    wire N__20291;
    wire N__20286;
    wire N__20285;
    wire N__20284;
    wire N__20283;
    wire N__20282;
    wire N__20281;
    wire N__20280;
    wire N__20277;
    wire N__20270;
    wire N__20263;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19908;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19706;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19499;
    wire N__19498;
    wire N__19493;
    wire N__19490;
    wire N__19485;
    wire N__19484;
    wire N__19483;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19464;
    wire N__19463;
    wire N__19460;
    wire N__19459;
    wire N__19456;
    wire N__19451;
    wire N__19448;
    wire N__19443;
    wire N__19442;
    wire N__19441;
    wire N__19436;
    wire N__19433;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19421;
    wire N__19420;
    wire N__19417;
    wire N__19412;
    wire N__19409;
    wire N__19404;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19392;
    wire N__19389;
    wire N__19388;
    wire N__19387;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19362;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19301;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19287;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19272;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire VCCG0;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_98_cascade_ ;
    wire bfn_1_16_0_;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire bfn_1_17_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire bfn_1_18_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_2_1_15 ;
    wire \pwm_generator_inst.un2_threshold_2_1_16 ;
    wire N_6_0;
    wire m38;
    wire pwm_duty_input_0;
    wire pwm_duty_input_1;
    wire pwm_duty_input_2;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ;
    wire pwm_duty_input_8;
    wire pwm_duty_input_9;
    wire pwm_duty_input_7;
    wire pwm_duty_input_6;
    wire \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ;
    wire pwm_duty_input_5;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_120 ;
    wire \current_shift_inst.PI_CTRL.N_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.N_97 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_306 ;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_0 ;
    wire bfn_2_12_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_8 ;
    wire bfn_2_13_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un15_threshold_1_cry_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15 ;
    wire bfn_2_14_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_4 ;
    wire bfn_2_15_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_1_20 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_1_21 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_1_22 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_1_23 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ;
    wire bfn_2_16_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_1_24 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_2_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un2_threshold_2_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un2_threshold_1_25 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15 ;
    wire \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_19_THRU_CO ;
    wire bfn_2_17_0_;
    wire \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un1_duty_inputlt3 ;
    wire pwm_duty_input_3;
    wire \pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ;
    wire bfn_3_15_0_;
    wire \pwm_generator_inst.un19_threshold_axb_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_0 ;
    wire \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_1 ;
    wire \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_2 ;
    wire \pwm_generator_inst.un19_threshold_axb_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_3 ;
    wire \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ;
    wire \pwm_generator_inst.un19_threshold_cry_4 ;
    wire \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_5 ;
    wire \pwm_generator_inst.un19_threshold_axb_7 ;
    wire \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ;
    wire \pwm_generator_inst.un19_threshold_cry_6 ;
    wire \pwm_generator_inst.un19_threshold_cry_7 ;
    wire \pwm_generator_inst.un19_threshold_axb_8 ;
    wire bfn_3_16_0_;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ;
    wire \pwm_generator_inst.un19_threshold_cry_8 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ;
    wire \pwm_generator_inst.un19_threshold_axb_6 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_5 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ;
    wire \pwm_generator_inst.un15_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ;
    wire \pwm_generator_inst.un19_threshold_axb_3 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un19_threshold_axb_0 ;
    wire \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ;
    wire \pwm_generator_inst.un15_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un19_threshold_axb_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ;
    wire bfn_3_18_0_;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire bfn_3_19_0_;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire \pwm_generator_inst.threshold_0 ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_4_13_0_;
    wire \pwm_generator_inst.un14_counter_1 ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.threshold_2 ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.threshold_3 ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.threshold_4 ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.threshold_5 ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.un14_counter_6 ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.un14_counter_7 ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_4_14_0_;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ;
    wire \pwm_generator_inst.un14_counter_8 ;
    wire \pwm_generator_inst.N_17 ;
    wire \pwm_generator_inst.N_16 ;
    wire N_19_1;
    wire \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ;
    wire \pwm_generator_inst.threshold_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire \current_shift_inst.PI_CTRL.N_118 ;
    wire bfn_5_15_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire bfn_5_16_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire bfn_5_17_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire bfn_5_18_0_;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ;
    wire bfn_7_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_7_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_7_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_7_13_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_343_i ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire bfn_8_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_8_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_8_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_8_12_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.N_344_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_8_17_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire bfn_8_18_0_;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire bfn_8_19_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire bfn_8_20_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire elapsed_time_ns_1_RNI1CPBB_0_23_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.N_43 ;
    wire \phase_controller_inst1.N_43_cascade_ ;
    wire \phase_controller_inst1.stoper_tr.N_43_0 ;
    wire \phase_controller_inst1.running ;
    wire \phase_controller_inst1.N_42_cascade_ ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire elapsed_time_ns_1_RNI4FPBB_0_26_cascade_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_1 ;
    wire bfn_11_5_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_9 ;
    wire bfn_11_6_0_;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_16 ;
    wire bfn_11_7_0_;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst2.un4_running_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt30 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_1 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_9 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_16 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_28 ;
    wire \phase_controller_inst1.un4_running_cry_30 ;
    wire \phase_controller_inst1.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.N_42 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ;
    wire bfn_11_12_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.N_42_i ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ;
    wire bfn_11_14_0_;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_11_15_0_;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ;
    wire bfn_11_16_0_;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_11_17_0_;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire bfn_11_18_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire bfn_11_19_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire s4_phy_c;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt24 ;
    wire \phase_controller_inst1.start_latched ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst2.N_38 ;
    wire bfn_12_8_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.N_38_i ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ;
    wire bfn_12_9_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ;
    wire bfn_12_10_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ;
    wire bfn_12_11_0_;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.m3_0 ;
    wire \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire bfn_12_13_0_;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire bfn_12_14_0_;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire bfn_12_15_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_12_16_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire s3_phy_c;
    wire GB_BUFFER_red_c_g_THRU_CO;
    wire \phase_controller_inst1.stoper_hc.m34_1 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_hc.m10Z0Z_1 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire \phase_controller_inst2.stoper_tr.un1_start_g ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire elapsed_time_ns_1_RNI6GOBB_0_19_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire \phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ;
    wire \phase_controller_inst1.m3 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.N_1275_i ;
    wire bfn_13_17_0_;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire bfn_13_18_0_;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire bfn_13_19_0_;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire bfn_13_20_0_;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst2.N_139_1 ;
    wire \phase_controller_inst2.stoper_hc.N_34 ;
    wire \phase_controller_inst2.stoper_hc.m20_nsZ0Z_1 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.stoper_hc.hc_time_passed ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.N_266_0 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire delay_hc_input_c_g;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.N_339_i_g ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.control_input_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire bfn_14_21_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire s2_phy_c;
    wire \phase_controller_inst1.stoper_hc.m19_ns_1 ;
    wire \phase_controller_inst1.stoper_hc.N_27 ;
    wire il_max_comp1_c;
    wire \phase_controller_inst1.N_175_1 ;
    wire \phase_controller_inst1.stoper_hc.N_8_0_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.m12_ns_1 ;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.N_14_0 ;
    wire \phase_controller_inst1.N_13_0 ;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst2.m21 ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.time_passed_er_RNI23UO1 ;
    wire s1_phy_c;
    wire bfn_15_5_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.N_45_i ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_15_6_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_15_7_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_15_8_0_;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire S1_RNI9RLH;
    wire \current_shift_inst.PI_CTRL.N_77_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_286 ;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.N_339_i ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ;
    wire \phase_controller_inst1.stateZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.N_8_0 ;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire test22_c;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_1 ;
    wire bfn_16_6_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_9 ;
    wire bfn_16_7_0_;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_16 ;
    wire bfn_16_8_0_;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire bfn_16_14_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_16_17_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.N_340_i ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12_cascade_;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_287_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ;
    wire \phase_controller_inst1.stoper_hc.hc_time_passed ;
    wire \phase_controller_inst1.stoper_hc.N_45 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.N_46 ;
    wire \phase_controller_inst1.stoper_hc.N_46_cascade_ ;
    wire \phase_controller_inst1.stoper_hc.N_46_0 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire \phase_controller_inst1.stoper_hc.un4_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.N_342_i ;
    wire bfn_17_14_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.N_265_i ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ;
    wire bfn_17_15_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ;
    wire bfn_17_16_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ;
    wire bfn_17_17_0_;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.N_47 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.mZ0Z16 ;
    wire \phase_controller_inst2.stoper_hc.m28_ns_1 ;
    wire \phase_controller_inst2.stateZ0Z_4 ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire bfn_17_21_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire bfn_17_22_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire bfn_17_23_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ;
    wire GNDG0;
    wire \phase_controller_inst1.stateZ0Z_5 ;
    wire test_c;
    wire start_stop_c;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ;
    wire \phase_controller_inst2.start_latched ;
    wire \phase_controller_inst2.running ;
    wire \phase_controller_inst2.N_39 ;
    wire \phase_controller_inst2.stoper_tr.N_39_0 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire elapsed_time_ns_1_RNI02CN9_0_13_cascade_;
    wire bfn_18_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_18_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_18_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_18_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire elapsed_time_ns_1_RNI46CN9_0_17_cascade_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_1 ;
    wire bfn_18_16_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_8 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_9 ;
    wire bfn_18_17_0_;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_time_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_15 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt18 ;
    wire bfn_18_18_0_;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_0_30 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.N_289 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.N_290 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire bfn_18_22_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire bfn_18_23_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire GB_BUFFER_clock_output_0_THRU_CO;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9_cascade_;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.N_341_i ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.un1_start_g ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.un4_running_lt22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire clock_output_0;
    wire red_c_g;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__25797),
            .RESETB(N__31242),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clock_output_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__49826),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__49816),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__37148,N__37188,N__37230,N__37274,N__37317,N__36822,N__36870,N__36906,N__36938,N__36984,N__37022,N__37059,N__36494,N__36531,N__36579,N__36612}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__49818,dangling_wire_45,N__49817}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__49872),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__49865),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__21601,N__21594,N__21599,N__21593,N__21600,N__21592,N__21602,N__21589,N__21595,N__21588,N__21596,N__21590,N__21597,N__21591,N__21598}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,N__49871,N__49868,dangling_wire_102,dangling_wire_103,dangling_wire_104,N__49866,N__49870,N__49867,N__49869}),
            .OHOLDTOP(),
            .O({dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,\pwm_generator_inst.un2_threshold_2_1_16 ,\pwm_generator_inst.un2_threshold_2_1_15 ,\pwm_generator_inst.un2_threshold_2_14 ,\pwm_generator_inst.un2_threshold_2_13 ,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__49797),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__49790),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135}),
            .ADDSUBBOT(),
            .A({dangling_wire_136,N__21562,N__21565,N__21563,N__21566,N__21564,N__19483,N__19498,N__19463,N__19441,N__19425,N__20517,N__20542,N__19272,N__19287,N__19302}),
            .C({dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152}),
            .B({dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,N__49796,N__49793,dangling_wire_160,dangling_wire_161,dangling_wire_162,N__49791,N__49795,N__49792,N__49794}),
            .OHOLDTOP(),
            .O({dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,\pwm_generator_inst.un2_threshold_1_25 ,\pwm_generator_inst.un2_threshold_1_24 ,\pwm_generator_inst.un2_threshold_1_23 ,\pwm_generator_inst.un2_threshold_1_22 ,\pwm_generator_inst.un2_threshold_1_21 ,\pwm_generator_inst.un2_threshold_1_20 ,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__49825),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__49658),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184}),
            .ADDSUBBOT(),
            .A({dangling_wire_185,N__36644,N__36680,N__36726,N__36768,N__36240,N__36282,N__38229,N__36321,N__36363,N__36395,N__50967,N__36450,N__35970,N__36015,N__30695}),
            .C({dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201}),
            .B({dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,N__49660,dangling_wire_215,N__49659}),
            .OHOLDTOP(),
            .O({dangling_wire_216,dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__51919),
            .GLOBALBUFFEROUTPUT(red_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__51921),
            .DIN(N__51920),
            .DOUT(N__51919),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__51921),
            .PADOUT(N__51920),
            .PADIN(N__51919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_output_obuf_iopad (
            .OE(N__51910),
            .DIN(N__51909),
            .DOUT(N__51908),
            .PACKAGEPIN(clock_output));
    defparam clock_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam clock_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO clock_output_obuf_preio (
            .PADOEN(N__51910),
            .PADOUT(N__51909),
            .PADIN(N__51908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__47493),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test_obuf_iopad (
            .OE(N__51901),
            .DIN(N__51900),
            .DOUT(N__51899),
            .PACKAGEPIN(test));
    defparam test_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test_obuf_preio (
            .PADOEN(N__51901),
            .PADOUT(N__51900),
            .PADIN(N__51899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__43701),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__51892),
            .DIN(N__51891),
            .DOUT(N__51890),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__51892),
            .PADOUT(N__51891),
            .PADIN(N__51890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__51883),
            .DIN(N__51882),
            .DOUT(N__51881),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__51883),
            .PADOUT(N__51882),
            .PADIN(N__51881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__51874),
            .DIN(N__51873),
            .DOUT(N__51872),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__51874),
            .PADOUT(N__51873),
            .PADIN(N__51872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21750),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__51865),
            .DIN(N__51864),
            .DOUT(N__51863),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__51865),
            .PADOUT(N__51864),
            .PADIN(N__51863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__51856),
            .DIN(N__51855),
            .DOUT(N__51854),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__51856),
            .PADOUT(N__51855),
            .PADIN(N__51854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37086),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD test22_obuf_iopad (
            .OE(N__51847),
            .DIN(N__51846),
            .DOUT(N__51845),
            .PACKAGEPIN(test22));
    defparam test22_obuf_preio.NEG_TRIGGER=1'b0;
    defparam test22_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO test22_obuf_preio (
            .PADOEN(N__51847),
            .PADOUT(N__51846),
            .PADIN(N__51845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38745),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__51838),
            .DIN(N__51837),
            .DOUT(N__51836),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__51838),
            .PADOUT(N__51837),
            .PADIN(N__51836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__51829),
            .DIN(N__51828),
            .DOUT(N__51827),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__51829),
            .PADOUT(N__51828),
            .PADIN(N__51827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37347),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__51820),
            .DIN(N__51819),
            .DOUT(N__51818),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__51820),
            .PADOUT(N__51819),
            .PADIN(N__51818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__28593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__51811),
            .DIN(N__51810),
            .DOUT(N__51809),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__51811),
            .PADOUT(N__51810),
            .PADIN(N__51809),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__51802),
            .DIN(N__51801),
            .DOUT(N__51800),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__51802),
            .PADOUT(N__51801),
            .PADIN(N__51800),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31257),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__51793),
            .DIN(N__51792),
            .DOUT(N__51791),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__51793),
            .PADOUT(N__51792),
            .PADIN(N__51791),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__51784),
            .DIN(N__51783),
            .DOUT(N__51782),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__51784),
            .PADOUT(N__51783),
            .PADIN(N__51782),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__12456 (
            .O(N__51765),
            .I(N__51759));
    InMux I__12455 (
            .O(N__51764),
            .I(N__51756));
    InMux I__12454 (
            .O(N__51763),
            .I(N__51753));
    InMux I__12453 (
            .O(N__51762),
            .I(N__51750));
    LocalMux I__12452 (
            .O(N__51759),
            .I(N__51747));
    LocalMux I__12451 (
            .O(N__51756),
            .I(N__51744));
    LocalMux I__12450 (
            .O(N__51753),
            .I(N__51741));
    LocalMux I__12449 (
            .O(N__51750),
            .I(N__51738));
    Span4Mux_h I__12448 (
            .O(N__51747),
            .I(N__51735));
    Span4Mux_h I__12447 (
            .O(N__51744),
            .I(N__51730));
    Span4Mux_h I__12446 (
            .O(N__51741),
            .I(N__51730));
    Odrv4 I__12445 (
            .O(N__51738),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__12444 (
            .O(N__51735),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    Odrv4 I__12443 (
            .O(N__51730),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    InMux I__12442 (
            .O(N__51723),
            .I(N__51720));
    LocalMux I__12441 (
            .O(N__51720),
            .I(N__51717));
    Span4Mux_v I__12440 (
            .O(N__51717),
            .I(N__51712));
    InMux I__12439 (
            .O(N__51716),
            .I(N__51709));
    InMux I__12438 (
            .O(N__51715),
            .I(N__51706));
    Span4Mux_h I__12437 (
            .O(N__51712),
            .I(N__51701));
    LocalMux I__12436 (
            .O(N__51709),
            .I(N__51701));
    LocalMux I__12435 (
            .O(N__51706),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    Odrv4 I__12434 (
            .O(N__51701),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    InMux I__12433 (
            .O(N__51696),
            .I(N__51690));
    InMux I__12432 (
            .O(N__51695),
            .I(N__51687));
    InMux I__12431 (
            .O(N__51694),
            .I(N__51684));
    InMux I__12430 (
            .O(N__51693),
            .I(N__51681));
    LocalMux I__12429 (
            .O(N__51690),
            .I(N__51678));
    LocalMux I__12428 (
            .O(N__51687),
            .I(N__51675));
    LocalMux I__12427 (
            .O(N__51684),
            .I(N__51672));
    LocalMux I__12426 (
            .O(N__51681),
            .I(N__51669));
    Span4Mux_v I__12425 (
            .O(N__51678),
            .I(N__51664));
    Span4Mux_v I__12424 (
            .O(N__51675),
            .I(N__51664));
    Span4Mux_h I__12423 (
            .O(N__51672),
            .I(N__51661));
    Odrv12 I__12422 (
            .O(N__51669),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__12421 (
            .O(N__51664),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__12420 (
            .O(N__51661),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__12419 (
            .O(N__51654),
            .I(N__51650));
    InMux I__12418 (
            .O(N__51653),
            .I(N__51647));
    LocalMux I__12417 (
            .O(N__51650),
            .I(N__51643));
    LocalMux I__12416 (
            .O(N__51647),
            .I(N__51640));
    InMux I__12415 (
            .O(N__51646),
            .I(N__51637));
    Span4Mux_h I__12414 (
            .O(N__51643),
            .I(N__51634));
    Span4Mux_v I__12413 (
            .O(N__51640),
            .I(N__51631));
    LocalMux I__12412 (
            .O(N__51637),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__12411 (
            .O(N__51634),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    Odrv4 I__12410 (
            .O(N__51631),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    CascadeMux I__12409 (
            .O(N__51624),
            .I(N__51613));
    InMux I__12408 (
            .O(N__51623),
            .I(N__51605));
    InMux I__12407 (
            .O(N__51622),
            .I(N__51605));
    InMux I__12406 (
            .O(N__51621),
            .I(N__51605));
    InMux I__12405 (
            .O(N__51620),
            .I(N__51597));
    InMux I__12404 (
            .O(N__51619),
            .I(N__51589));
    InMux I__12403 (
            .O(N__51618),
            .I(N__51582));
    InMux I__12402 (
            .O(N__51617),
            .I(N__51582));
    InMux I__12401 (
            .O(N__51616),
            .I(N__51582));
    InMux I__12400 (
            .O(N__51613),
            .I(N__51574));
    InMux I__12399 (
            .O(N__51612),
            .I(N__51574));
    LocalMux I__12398 (
            .O(N__51605),
            .I(N__51571));
    InMux I__12397 (
            .O(N__51604),
            .I(N__51560));
    InMux I__12396 (
            .O(N__51603),
            .I(N__51560));
    InMux I__12395 (
            .O(N__51602),
            .I(N__51560));
    InMux I__12394 (
            .O(N__51601),
            .I(N__51560));
    InMux I__12393 (
            .O(N__51600),
            .I(N__51560));
    LocalMux I__12392 (
            .O(N__51597),
            .I(N__51548));
    InMux I__12391 (
            .O(N__51596),
            .I(N__51543));
    InMux I__12390 (
            .O(N__51595),
            .I(N__51543));
    InMux I__12389 (
            .O(N__51594),
            .I(N__51536));
    InMux I__12388 (
            .O(N__51593),
            .I(N__51536));
    InMux I__12387 (
            .O(N__51592),
            .I(N__51536));
    LocalMux I__12386 (
            .O(N__51589),
            .I(N__51531));
    LocalMux I__12385 (
            .O(N__51582),
            .I(N__51531));
    InMux I__12384 (
            .O(N__51581),
            .I(N__51526));
    InMux I__12383 (
            .O(N__51580),
            .I(N__51526));
    CascadeMux I__12382 (
            .O(N__51579),
            .I(N__51523));
    LocalMux I__12381 (
            .O(N__51574),
            .I(N__51508));
    Span4Mux_v I__12380 (
            .O(N__51571),
            .I(N__51508));
    LocalMux I__12379 (
            .O(N__51560),
            .I(N__51508));
    InMux I__12378 (
            .O(N__51559),
            .I(N__51505));
    InMux I__12377 (
            .O(N__51558),
            .I(N__51494));
    InMux I__12376 (
            .O(N__51557),
            .I(N__51494));
    InMux I__12375 (
            .O(N__51556),
            .I(N__51494));
    InMux I__12374 (
            .O(N__51555),
            .I(N__51491));
    InMux I__12373 (
            .O(N__51554),
            .I(N__51488));
    InMux I__12372 (
            .O(N__51553),
            .I(N__51483));
    InMux I__12371 (
            .O(N__51552),
            .I(N__51483));
    InMux I__12370 (
            .O(N__51551),
            .I(N__51480));
    Span4Mux_v I__12369 (
            .O(N__51548),
            .I(N__51469));
    LocalMux I__12368 (
            .O(N__51543),
            .I(N__51469));
    LocalMux I__12367 (
            .O(N__51536),
            .I(N__51469));
    Span4Mux_v I__12366 (
            .O(N__51531),
            .I(N__51469));
    LocalMux I__12365 (
            .O(N__51526),
            .I(N__51469));
    InMux I__12364 (
            .O(N__51523),
            .I(N__51464));
    InMux I__12363 (
            .O(N__51522),
            .I(N__51464));
    InMux I__12362 (
            .O(N__51521),
            .I(N__51461));
    CascadeMux I__12361 (
            .O(N__51520),
            .I(N__51457));
    InMux I__12360 (
            .O(N__51519),
            .I(N__51450));
    InMux I__12359 (
            .O(N__51518),
            .I(N__51450));
    InMux I__12358 (
            .O(N__51517),
            .I(N__51450));
    CascadeMux I__12357 (
            .O(N__51516),
            .I(N__51447));
    InMux I__12356 (
            .O(N__51515),
            .I(N__51427));
    Span4Mux_v I__12355 (
            .O(N__51508),
            .I(N__51422));
    LocalMux I__12354 (
            .O(N__51505),
            .I(N__51422));
    InMux I__12353 (
            .O(N__51504),
            .I(N__51419));
    InMux I__12352 (
            .O(N__51503),
            .I(N__51416));
    InMux I__12351 (
            .O(N__51502),
            .I(N__51410));
    InMux I__12350 (
            .O(N__51501),
            .I(N__51410));
    LocalMux I__12349 (
            .O(N__51494),
            .I(N__51395));
    LocalMux I__12348 (
            .O(N__51491),
            .I(N__51395));
    LocalMux I__12347 (
            .O(N__51488),
            .I(N__51395));
    LocalMux I__12346 (
            .O(N__51483),
            .I(N__51395));
    LocalMux I__12345 (
            .O(N__51480),
            .I(N__51395));
    Span4Mux_v I__12344 (
            .O(N__51469),
            .I(N__51395));
    LocalMux I__12343 (
            .O(N__51464),
            .I(N__51395));
    LocalMux I__12342 (
            .O(N__51461),
            .I(N__51392));
    CascadeMux I__12341 (
            .O(N__51460),
            .I(N__51383));
    InMux I__12340 (
            .O(N__51457),
            .I(N__51380));
    LocalMux I__12339 (
            .O(N__51450),
            .I(N__51377));
    InMux I__12338 (
            .O(N__51447),
            .I(N__51374));
    InMux I__12337 (
            .O(N__51446),
            .I(N__51369));
    InMux I__12336 (
            .O(N__51445),
            .I(N__51369));
    InMux I__12335 (
            .O(N__51444),
            .I(N__51362));
    InMux I__12334 (
            .O(N__51443),
            .I(N__51362));
    InMux I__12333 (
            .O(N__51442),
            .I(N__51362));
    InMux I__12332 (
            .O(N__51441),
            .I(N__51351));
    InMux I__12331 (
            .O(N__51440),
            .I(N__51351));
    InMux I__12330 (
            .O(N__51439),
            .I(N__51351));
    InMux I__12329 (
            .O(N__51438),
            .I(N__51351));
    InMux I__12328 (
            .O(N__51437),
            .I(N__51351));
    InMux I__12327 (
            .O(N__51436),
            .I(N__51346));
    InMux I__12326 (
            .O(N__51435),
            .I(N__51346));
    InMux I__12325 (
            .O(N__51434),
            .I(N__51341));
    InMux I__12324 (
            .O(N__51433),
            .I(N__51341));
    InMux I__12323 (
            .O(N__51432),
            .I(N__51336));
    InMux I__12322 (
            .O(N__51431),
            .I(N__51336));
    InMux I__12321 (
            .O(N__51430),
            .I(N__51333));
    LocalMux I__12320 (
            .O(N__51427),
            .I(N__51326));
    Span4Mux_h I__12319 (
            .O(N__51422),
            .I(N__51326));
    LocalMux I__12318 (
            .O(N__51419),
            .I(N__51326));
    LocalMux I__12317 (
            .O(N__51416),
            .I(N__51323));
    InMux I__12316 (
            .O(N__51415),
            .I(N__51310));
    LocalMux I__12315 (
            .O(N__51410),
            .I(N__51307));
    Span4Mux_v I__12314 (
            .O(N__51395),
            .I(N__51302));
    Span4Mux_v I__12313 (
            .O(N__51392),
            .I(N__51302));
    InMux I__12312 (
            .O(N__51391),
            .I(N__51289));
    InMux I__12311 (
            .O(N__51390),
            .I(N__51289));
    InMux I__12310 (
            .O(N__51389),
            .I(N__51289));
    InMux I__12309 (
            .O(N__51388),
            .I(N__51289));
    InMux I__12308 (
            .O(N__51387),
            .I(N__51275));
    InMux I__12307 (
            .O(N__51386),
            .I(N__51275));
    InMux I__12306 (
            .O(N__51383),
            .I(N__51272));
    LocalMux I__12305 (
            .O(N__51380),
            .I(N__51269));
    Span4Mux_h I__12304 (
            .O(N__51377),
            .I(N__51264));
    LocalMux I__12303 (
            .O(N__51374),
            .I(N__51264));
    LocalMux I__12302 (
            .O(N__51369),
            .I(N__51261));
    LocalMux I__12301 (
            .O(N__51362),
            .I(N__51254));
    LocalMux I__12300 (
            .O(N__51351),
            .I(N__51254));
    LocalMux I__12299 (
            .O(N__51346),
            .I(N__51254));
    LocalMux I__12298 (
            .O(N__51341),
            .I(N__51251));
    LocalMux I__12297 (
            .O(N__51336),
            .I(N__51242));
    LocalMux I__12296 (
            .O(N__51333),
            .I(N__51242));
    Span4Mux_v I__12295 (
            .O(N__51326),
            .I(N__51242));
    Span4Mux_v I__12294 (
            .O(N__51323),
            .I(N__51242));
    InMux I__12293 (
            .O(N__51322),
            .I(N__51233));
    InMux I__12292 (
            .O(N__51321),
            .I(N__51233));
    InMux I__12291 (
            .O(N__51320),
            .I(N__51233));
    InMux I__12290 (
            .O(N__51319),
            .I(N__51233));
    InMux I__12289 (
            .O(N__51318),
            .I(N__51230));
    InMux I__12288 (
            .O(N__51317),
            .I(N__51227));
    InMux I__12287 (
            .O(N__51316),
            .I(N__51218));
    InMux I__12286 (
            .O(N__51315),
            .I(N__51218));
    InMux I__12285 (
            .O(N__51314),
            .I(N__51218));
    InMux I__12284 (
            .O(N__51313),
            .I(N__51218));
    LocalMux I__12283 (
            .O(N__51310),
            .I(N__51211));
    Span4Mux_v I__12282 (
            .O(N__51307),
            .I(N__51211));
    Span4Mux_h I__12281 (
            .O(N__51302),
            .I(N__51211));
    InMux I__12280 (
            .O(N__51301),
            .I(N__51206));
    InMux I__12279 (
            .O(N__51300),
            .I(N__51206));
    InMux I__12278 (
            .O(N__51299),
            .I(N__51203));
    InMux I__12277 (
            .O(N__51298),
            .I(N__51200));
    LocalMux I__12276 (
            .O(N__51289),
            .I(N__51197));
    InMux I__12275 (
            .O(N__51288),
            .I(N__51190));
    InMux I__12274 (
            .O(N__51287),
            .I(N__51190));
    InMux I__12273 (
            .O(N__51286),
            .I(N__51190));
    InMux I__12272 (
            .O(N__51285),
            .I(N__51183));
    InMux I__12271 (
            .O(N__51284),
            .I(N__51183));
    InMux I__12270 (
            .O(N__51283),
            .I(N__51183));
    InMux I__12269 (
            .O(N__51282),
            .I(N__51176));
    InMux I__12268 (
            .O(N__51281),
            .I(N__51176));
    InMux I__12267 (
            .O(N__51280),
            .I(N__51176));
    LocalMux I__12266 (
            .O(N__51275),
            .I(N__51159));
    LocalMux I__12265 (
            .O(N__51272),
            .I(N__51159));
    Span4Mux_v I__12264 (
            .O(N__51269),
            .I(N__51159));
    Span4Mux_v I__12263 (
            .O(N__51264),
            .I(N__51159));
    Span4Mux_v I__12262 (
            .O(N__51261),
            .I(N__51159));
    Span4Mux_v I__12261 (
            .O(N__51254),
            .I(N__51159));
    Span4Mux_h I__12260 (
            .O(N__51251),
            .I(N__51159));
    Span4Mux_h I__12259 (
            .O(N__51242),
            .I(N__51159));
    LocalMux I__12258 (
            .O(N__51233),
            .I(N__51148));
    LocalMux I__12257 (
            .O(N__51230),
            .I(N__51148));
    LocalMux I__12256 (
            .O(N__51227),
            .I(N__51148));
    LocalMux I__12255 (
            .O(N__51218),
            .I(N__51148));
    Span4Mux_v I__12254 (
            .O(N__51211),
            .I(N__51148));
    LocalMux I__12253 (
            .O(N__51206),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__12252 (
            .O(N__51203),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__12251 (
            .O(N__51200),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__12250 (
            .O(N__51197),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__12249 (
            .O(N__51190),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__12248 (
            .O(N__51183),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    LocalMux I__12247 (
            .O(N__51176),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__12246 (
            .O(N__51159),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__12245 (
            .O(N__51148),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__12244 (
            .O(N__51129),
            .I(N__51124));
    InMux I__12243 (
            .O(N__51128),
            .I(N__51120));
    InMux I__12242 (
            .O(N__51127),
            .I(N__51117));
    LocalMux I__12241 (
            .O(N__51124),
            .I(N__51114));
    InMux I__12240 (
            .O(N__51123),
            .I(N__51111));
    LocalMux I__12239 (
            .O(N__51120),
            .I(N__51108));
    LocalMux I__12238 (
            .O(N__51117),
            .I(N__51103));
    Span4Mux_v I__12237 (
            .O(N__51114),
            .I(N__51103));
    LocalMux I__12236 (
            .O(N__51111),
            .I(N__51100));
    Span4Mux_v I__12235 (
            .O(N__51108),
            .I(N__51097));
    Span4Mux_h I__12234 (
            .O(N__51103),
            .I(N__51092));
    Span4Mux_h I__12233 (
            .O(N__51100),
            .I(N__51092));
    Odrv4 I__12232 (
            .O(N__51097),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    Odrv4 I__12231 (
            .O(N__51092),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__12230 (
            .O(N__51087),
            .I(N__51083));
    InMux I__12229 (
            .O(N__51086),
            .I(N__51079));
    LocalMux I__12228 (
            .O(N__51083),
            .I(N__51076));
    InMux I__12227 (
            .O(N__51082),
            .I(N__51073));
    LocalMux I__12226 (
            .O(N__51079),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    Odrv4 I__12225 (
            .O(N__51076),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    LocalMux I__12224 (
            .O(N__51073),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__12223 (
            .O(N__51066),
            .I(N__51062));
    InMux I__12222 (
            .O(N__51065),
            .I(N__51059));
    LocalMux I__12221 (
            .O(N__51062),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    LocalMux I__12220 (
            .O(N__51059),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ));
    InMux I__12219 (
            .O(N__51054),
            .I(N__51051));
    LocalMux I__12218 (
            .O(N__51051),
            .I(N__51047));
    InMux I__12217 (
            .O(N__51050),
            .I(N__51044));
    Span4Mux_h I__12216 (
            .O(N__51047),
            .I(N__51038));
    LocalMux I__12215 (
            .O(N__51044),
            .I(N__51038));
    InMux I__12214 (
            .O(N__51043),
            .I(N__51035));
    Span4Mux_h I__12213 (
            .O(N__51038),
            .I(N__51032));
    LocalMux I__12212 (
            .O(N__51035),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__12211 (
            .O(N__51032),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ));
    CascadeMux I__12210 (
            .O(N__51027),
            .I(N__51023));
    CascadeMux I__12209 (
            .O(N__51026),
            .I(N__51020));
    InMux I__12208 (
            .O(N__51023),
            .I(N__51017));
    InMux I__12207 (
            .O(N__51020),
            .I(N__51014));
    LocalMux I__12206 (
            .O(N__51017),
            .I(N__51008));
    LocalMux I__12205 (
            .O(N__51014),
            .I(N__51008));
    InMux I__12204 (
            .O(N__51013),
            .I(N__51005));
    Span4Mux_v I__12203 (
            .O(N__51008),
            .I(N__51002));
    LocalMux I__12202 (
            .O(N__51005),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__12201 (
            .O(N__51002),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__12200 (
            .O(N__50997),
            .I(N__50993));
    InMux I__12199 (
            .O(N__50996),
            .I(N__50990));
    LocalMux I__12198 (
            .O(N__50993),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    LocalMux I__12197 (
            .O(N__50990),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ));
    CascadeMux I__12196 (
            .O(N__50985),
            .I(N__50982));
    InMux I__12195 (
            .O(N__50982),
            .I(N__50979));
    LocalMux I__12194 (
            .O(N__50979),
            .I(N__50976));
    Span4Mux_h I__12193 (
            .O(N__50976),
            .I(N__50973));
    Span4Mux_v I__12192 (
            .O(N__50973),
            .I(N__50970));
    Odrv4 I__12191 (
            .O(N__50970),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt22 ));
    InMux I__12190 (
            .O(N__50967),
            .I(N__50963));
    InMux I__12189 (
            .O(N__50966),
            .I(N__50960));
    LocalMux I__12188 (
            .O(N__50963),
            .I(N__50957));
    LocalMux I__12187 (
            .O(N__50960),
            .I(N__50954));
    Span4Mux_v I__12186 (
            .O(N__50957),
            .I(N__50951));
    Span4Mux_v I__12185 (
            .O(N__50954),
            .I(N__50946));
    Span4Mux_v I__12184 (
            .O(N__50951),
            .I(N__50946));
    Sp12to4 I__12183 (
            .O(N__50946),
            .I(N__50943));
    Odrv12 I__12182 (
            .O(N__50943),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__12181 (
            .O(N__50940),
            .I(N__50937));
    LocalMux I__12180 (
            .O(N__50937),
            .I(N__50934));
    Span4Mux_h I__12179 (
            .O(N__50934),
            .I(N__50931));
    Span4Mux_h I__12178 (
            .O(N__50931),
            .I(N__50928));
    Span4Mux_h I__12177 (
            .O(N__50928),
            .I(N__50925));
    Span4Mux_h I__12176 (
            .O(N__50925),
            .I(N__50922));
    Odrv4 I__12175 (
            .O(N__50922),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    InMux I__12174 (
            .O(N__50919),
            .I(N__50916));
    LocalMux I__12173 (
            .O(N__50916),
            .I(N__50753));
    ClkMux I__12172 (
            .O(N__50915),
            .I(N__50421));
    ClkMux I__12171 (
            .O(N__50914),
            .I(N__50421));
    ClkMux I__12170 (
            .O(N__50913),
            .I(N__50421));
    ClkMux I__12169 (
            .O(N__50912),
            .I(N__50421));
    ClkMux I__12168 (
            .O(N__50911),
            .I(N__50421));
    ClkMux I__12167 (
            .O(N__50910),
            .I(N__50421));
    ClkMux I__12166 (
            .O(N__50909),
            .I(N__50421));
    ClkMux I__12165 (
            .O(N__50908),
            .I(N__50421));
    ClkMux I__12164 (
            .O(N__50907),
            .I(N__50421));
    ClkMux I__12163 (
            .O(N__50906),
            .I(N__50421));
    ClkMux I__12162 (
            .O(N__50905),
            .I(N__50421));
    ClkMux I__12161 (
            .O(N__50904),
            .I(N__50421));
    ClkMux I__12160 (
            .O(N__50903),
            .I(N__50421));
    ClkMux I__12159 (
            .O(N__50902),
            .I(N__50421));
    ClkMux I__12158 (
            .O(N__50901),
            .I(N__50421));
    ClkMux I__12157 (
            .O(N__50900),
            .I(N__50421));
    ClkMux I__12156 (
            .O(N__50899),
            .I(N__50421));
    ClkMux I__12155 (
            .O(N__50898),
            .I(N__50421));
    ClkMux I__12154 (
            .O(N__50897),
            .I(N__50421));
    ClkMux I__12153 (
            .O(N__50896),
            .I(N__50421));
    ClkMux I__12152 (
            .O(N__50895),
            .I(N__50421));
    ClkMux I__12151 (
            .O(N__50894),
            .I(N__50421));
    ClkMux I__12150 (
            .O(N__50893),
            .I(N__50421));
    ClkMux I__12149 (
            .O(N__50892),
            .I(N__50421));
    ClkMux I__12148 (
            .O(N__50891),
            .I(N__50421));
    ClkMux I__12147 (
            .O(N__50890),
            .I(N__50421));
    ClkMux I__12146 (
            .O(N__50889),
            .I(N__50421));
    ClkMux I__12145 (
            .O(N__50888),
            .I(N__50421));
    ClkMux I__12144 (
            .O(N__50887),
            .I(N__50421));
    ClkMux I__12143 (
            .O(N__50886),
            .I(N__50421));
    ClkMux I__12142 (
            .O(N__50885),
            .I(N__50421));
    ClkMux I__12141 (
            .O(N__50884),
            .I(N__50421));
    ClkMux I__12140 (
            .O(N__50883),
            .I(N__50421));
    ClkMux I__12139 (
            .O(N__50882),
            .I(N__50421));
    ClkMux I__12138 (
            .O(N__50881),
            .I(N__50421));
    ClkMux I__12137 (
            .O(N__50880),
            .I(N__50421));
    ClkMux I__12136 (
            .O(N__50879),
            .I(N__50421));
    ClkMux I__12135 (
            .O(N__50878),
            .I(N__50421));
    ClkMux I__12134 (
            .O(N__50877),
            .I(N__50421));
    ClkMux I__12133 (
            .O(N__50876),
            .I(N__50421));
    ClkMux I__12132 (
            .O(N__50875),
            .I(N__50421));
    ClkMux I__12131 (
            .O(N__50874),
            .I(N__50421));
    ClkMux I__12130 (
            .O(N__50873),
            .I(N__50421));
    ClkMux I__12129 (
            .O(N__50872),
            .I(N__50421));
    ClkMux I__12128 (
            .O(N__50871),
            .I(N__50421));
    ClkMux I__12127 (
            .O(N__50870),
            .I(N__50421));
    ClkMux I__12126 (
            .O(N__50869),
            .I(N__50421));
    ClkMux I__12125 (
            .O(N__50868),
            .I(N__50421));
    ClkMux I__12124 (
            .O(N__50867),
            .I(N__50421));
    ClkMux I__12123 (
            .O(N__50866),
            .I(N__50421));
    ClkMux I__12122 (
            .O(N__50865),
            .I(N__50421));
    ClkMux I__12121 (
            .O(N__50864),
            .I(N__50421));
    ClkMux I__12120 (
            .O(N__50863),
            .I(N__50421));
    ClkMux I__12119 (
            .O(N__50862),
            .I(N__50421));
    ClkMux I__12118 (
            .O(N__50861),
            .I(N__50421));
    ClkMux I__12117 (
            .O(N__50860),
            .I(N__50421));
    ClkMux I__12116 (
            .O(N__50859),
            .I(N__50421));
    ClkMux I__12115 (
            .O(N__50858),
            .I(N__50421));
    ClkMux I__12114 (
            .O(N__50857),
            .I(N__50421));
    ClkMux I__12113 (
            .O(N__50856),
            .I(N__50421));
    ClkMux I__12112 (
            .O(N__50855),
            .I(N__50421));
    ClkMux I__12111 (
            .O(N__50854),
            .I(N__50421));
    ClkMux I__12110 (
            .O(N__50853),
            .I(N__50421));
    ClkMux I__12109 (
            .O(N__50852),
            .I(N__50421));
    ClkMux I__12108 (
            .O(N__50851),
            .I(N__50421));
    ClkMux I__12107 (
            .O(N__50850),
            .I(N__50421));
    ClkMux I__12106 (
            .O(N__50849),
            .I(N__50421));
    ClkMux I__12105 (
            .O(N__50848),
            .I(N__50421));
    ClkMux I__12104 (
            .O(N__50847),
            .I(N__50421));
    ClkMux I__12103 (
            .O(N__50846),
            .I(N__50421));
    ClkMux I__12102 (
            .O(N__50845),
            .I(N__50421));
    ClkMux I__12101 (
            .O(N__50844),
            .I(N__50421));
    ClkMux I__12100 (
            .O(N__50843),
            .I(N__50421));
    ClkMux I__12099 (
            .O(N__50842),
            .I(N__50421));
    ClkMux I__12098 (
            .O(N__50841),
            .I(N__50421));
    ClkMux I__12097 (
            .O(N__50840),
            .I(N__50421));
    ClkMux I__12096 (
            .O(N__50839),
            .I(N__50421));
    ClkMux I__12095 (
            .O(N__50838),
            .I(N__50421));
    ClkMux I__12094 (
            .O(N__50837),
            .I(N__50421));
    ClkMux I__12093 (
            .O(N__50836),
            .I(N__50421));
    ClkMux I__12092 (
            .O(N__50835),
            .I(N__50421));
    ClkMux I__12091 (
            .O(N__50834),
            .I(N__50421));
    ClkMux I__12090 (
            .O(N__50833),
            .I(N__50421));
    ClkMux I__12089 (
            .O(N__50832),
            .I(N__50421));
    ClkMux I__12088 (
            .O(N__50831),
            .I(N__50421));
    ClkMux I__12087 (
            .O(N__50830),
            .I(N__50421));
    ClkMux I__12086 (
            .O(N__50829),
            .I(N__50421));
    ClkMux I__12085 (
            .O(N__50828),
            .I(N__50421));
    ClkMux I__12084 (
            .O(N__50827),
            .I(N__50421));
    ClkMux I__12083 (
            .O(N__50826),
            .I(N__50421));
    ClkMux I__12082 (
            .O(N__50825),
            .I(N__50421));
    ClkMux I__12081 (
            .O(N__50824),
            .I(N__50421));
    ClkMux I__12080 (
            .O(N__50823),
            .I(N__50421));
    ClkMux I__12079 (
            .O(N__50822),
            .I(N__50421));
    ClkMux I__12078 (
            .O(N__50821),
            .I(N__50421));
    ClkMux I__12077 (
            .O(N__50820),
            .I(N__50421));
    ClkMux I__12076 (
            .O(N__50819),
            .I(N__50421));
    ClkMux I__12075 (
            .O(N__50818),
            .I(N__50421));
    ClkMux I__12074 (
            .O(N__50817),
            .I(N__50421));
    ClkMux I__12073 (
            .O(N__50816),
            .I(N__50421));
    ClkMux I__12072 (
            .O(N__50815),
            .I(N__50421));
    ClkMux I__12071 (
            .O(N__50814),
            .I(N__50421));
    ClkMux I__12070 (
            .O(N__50813),
            .I(N__50421));
    ClkMux I__12069 (
            .O(N__50812),
            .I(N__50421));
    ClkMux I__12068 (
            .O(N__50811),
            .I(N__50421));
    ClkMux I__12067 (
            .O(N__50810),
            .I(N__50421));
    ClkMux I__12066 (
            .O(N__50809),
            .I(N__50421));
    ClkMux I__12065 (
            .O(N__50808),
            .I(N__50421));
    ClkMux I__12064 (
            .O(N__50807),
            .I(N__50421));
    ClkMux I__12063 (
            .O(N__50806),
            .I(N__50421));
    ClkMux I__12062 (
            .O(N__50805),
            .I(N__50421));
    ClkMux I__12061 (
            .O(N__50804),
            .I(N__50421));
    ClkMux I__12060 (
            .O(N__50803),
            .I(N__50421));
    ClkMux I__12059 (
            .O(N__50802),
            .I(N__50421));
    ClkMux I__12058 (
            .O(N__50801),
            .I(N__50421));
    ClkMux I__12057 (
            .O(N__50800),
            .I(N__50421));
    ClkMux I__12056 (
            .O(N__50799),
            .I(N__50421));
    ClkMux I__12055 (
            .O(N__50798),
            .I(N__50421));
    ClkMux I__12054 (
            .O(N__50797),
            .I(N__50421));
    ClkMux I__12053 (
            .O(N__50796),
            .I(N__50421));
    ClkMux I__12052 (
            .O(N__50795),
            .I(N__50421));
    ClkMux I__12051 (
            .O(N__50794),
            .I(N__50421));
    ClkMux I__12050 (
            .O(N__50793),
            .I(N__50421));
    ClkMux I__12049 (
            .O(N__50792),
            .I(N__50421));
    ClkMux I__12048 (
            .O(N__50791),
            .I(N__50421));
    ClkMux I__12047 (
            .O(N__50790),
            .I(N__50421));
    ClkMux I__12046 (
            .O(N__50789),
            .I(N__50421));
    ClkMux I__12045 (
            .O(N__50788),
            .I(N__50421));
    ClkMux I__12044 (
            .O(N__50787),
            .I(N__50421));
    ClkMux I__12043 (
            .O(N__50786),
            .I(N__50421));
    ClkMux I__12042 (
            .O(N__50785),
            .I(N__50421));
    ClkMux I__12041 (
            .O(N__50784),
            .I(N__50421));
    ClkMux I__12040 (
            .O(N__50783),
            .I(N__50421));
    ClkMux I__12039 (
            .O(N__50782),
            .I(N__50421));
    ClkMux I__12038 (
            .O(N__50781),
            .I(N__50421));
    ClkMux I__12037 (
            .O(N__50780),
            .I(N__50421));
    ClkMux I__12036 (
            .O(N__50779),
            .I(N__50421));
    ClkMux I__12035 (
            .O(N__50778),
            .I(N__50421));
    ClkMux I__12034 (
            .O(N__50777),
            .I(N__50421));
    ClkMux I__12033 (
            .O(N__50776),
            .I(N__50421));
    ClkMux I__12032 (
            .O(N__50775),
            .I(N__50421));
    ClkMux I__12031 (
            .O(N__50774),
            .I(N__50421));
    ClkMux I__12030 (
            .O(N__50773),
            .I(N__50421));
    ClkMux I__12029 (
            .O(N__50772),
            .I(N__50421));
    ClkMux I__12028 (
            .O(N__50771),
            .I(N__50421));
    ClkMux I__12027 (
            .O(N__50770),
            .I(N__50421));
    ClkMux I__12026 (
            .O(N__50769),
            .I(N__50421));
    ClkMux I__12025 (
            .O(N__50768),
            .I(N__50421));
    ClkMux I__12024 (
            .O(N__50767),
            .I(N__50421));
    ClkMux I__12023 (
            .O(N__50766),
            .I(N__50421));
    ClkMux I__12022 (
            .O(N__50765),
            .I(N__50421));
    ClkMux I__12021 (
            .O(N__50764),
            .I(N__50421));
    ClkMux I__12020 (
            .O(N__50763),
            .I(N__50421));
    ClkMux I__12019 (
            .O(N__50762),
            .I(N__50421));
    ClkMux I__12018 (
            .O(N__50761),
            .I(N__50421));
    ClkMux I__12017 (
            .O(N__50760),
            .I(N__50421));
    ClkMux I__12016 (
            .O(N__50759),
            .I(N__50421));
    ClkMux I__12015 (
            .O(N__50758),
            .I(N__50421));
    ClkMux I__12014 (
            .O(N__50757),
            .I(N__50421));
    ClkMux I__12013 (
            .O(N__50756),
            .I(N__50421));
    Glb2LocalMux I__12012 (
            .O(N__50753),
            .I(N__50421));
    ClkMux I__12011 (
            .O(N__50752),
            .I(N__50421));
    ClkMux I__12010 (
            .O(N__50751),
            .I(N__50421));
    ClkMux I__12009 (
            .O(N__50750),
            .I(N__50421));
    GlobalMux I__12008 (
            .O(N__50421),
            .I(clock_output_0));
    InMux I__12007 (
            .O(N__50418),
            .I(N__50412));
    InMux I__12006 (
            .O(N__50417),
            .I(N__50407));
    InMux I__12005 (
            .O(N__50416),
            .I(N__50407));
    InMux I__12004 (
            .O(N__50415),
            .I(N__50404));
    LocalMux I__12003 (
            .O(N__50412),
            .I(N__50401));
    LocalMux I__12002 (
            .O(N__50407),
            .I(N__50398));
    LocalMux I__12001 (
            .O(N__50404),
            .I(N__50395));
    Glb2LocalMux I__12000 (
            .O(N__50401),
            .I(N__49890));
    Glb2LocalMux I__11999 (
            .O(N__50398),
            .I(N__49890));
    Glb2LocalMux I__11998 (
            .O(N__50395),
            .I(N__49890));
    SRMux I__11997 (
            .O(N__50394),
            .I(N__49890));
    SRMux I__11996 (
            .O(N__50393),
            .I(N__49890));
    SRMux I__11995 (
            .O(N__50392),
            .I(N__49890));
    SRMux I__11994 (
            .O(N__50391),
            .I(N__49890));
    SRMux I__11993 (
            .O(N__50390),
            .I(N__49890));
    SRMux I__11992 (
            .O(N__50389),
            .I(N__49890));
    SRMux I__11991 (
            .O(N__50388),
            .I(N__49890));
    SRMux I__11990 (
            .O(N__50387),
            .I(N__49890));
    SRMux I__11989 (
            .O(N__50386),
            .I(N__49890));
    SRMux I__11988 (
            .O(N__50385),
            .I(N__49890));
    SRMux I__11987 (
            .O(N__50384),
            .I(N__49890));
    SRMux I__11986 (
            .O(N__50383),
            .I(N__49890));
    SRMux I__11985 (
            .O(N__50382),
            .I(N__49890));
    SRMux I__11984 (
            .O(N__50381),
            .I(N__49890));
    SRMux I__11983 (
            .O(N__50380),
            .I(N__49890));
    SRMux I__11982 (
            .O(N__50379),
            .I(N__49890));
    SRMux I__11981 (
            .O(N__50378),
            .I(N__49890));
    SRMux I__11980 (
            .O(N__50377),
            .I(N__49890));
    SRMux I__11979 (
            .O(N__50376),
            .I(N__49890));
    SRMux I__11978 (
            .O(N__50375),
            .I(N__49890));
    SRMux I__11977 (
            .O(N__50374),
            .I(N__49890));
    SRMux I__11976 (
            .O(N__50373),
            .I(N__49890));
    SRMux I__11975 (
            .O(N__50372),
            .I(N__49890));
    SRMux I__11974 (
            .O(N__50371),
            .I(N__49890));
    SRMux I__11973 (
            .O(N__50370),
            .I(N__49890));
    SRMux I__11972 (
            .O(N__50369),
            .I(N__49890));
    SRMux I__11971 (
            .O(N__50368),
            .I(N__49890));
    SRMux I__11970 (
            .O(N__50367),
            .I(N__49890));
    SRMux I__11969 (
            .O(N__50366),
            .I(N__49890));
    SRMux I__11968 (
            .O(N__50365),
            .I(N__49890));
    SRMux I__11967 (
            .O(N__50364),
            .I(N__49890));
    SRMux I__11966 (
            .O(N__50363),
            .I(N__49890));
    SRMux I__11965 (
            .O(N__50362),
            .I(N__49890));
    SRMux I__11964 (
            .O(N__50361),
            .I(N__49890));
    SRMux I__11963 (
            .O(N__50360),
            .I(N__49890));
    SRMux I__11962 (
            .O(N__50359),
            .I(N__49890));
    SRMux I__11961 (
            .O(N__50358),
            .I(N__49890));
    SRMux I__11960 (
            .O(N__50357),
            .I(N__49890));
    SRMux I__11959 (
            .O(N__50356),
            .I(N__49890));
    SRMux I__11958 (
            .O(N__50355),
            .I(N__49890));
    SRMux I__11957 (
            .O(N__50354),
            .I(N__49890));
    SRMux I__11956 (
            .O(N__50353),
            .I(N__49890));
    SRMux I__11955 (
            .O(N__50352),
            .I(N__49890));
    SRMux I__11954 (
            .O(N__50351),
            .I(N__49890));
    SRMux I__11953 (
            .O(N__50350),
            .I(N__49890));
    SRMux I__11952 (
            .O(N__50349),
            .I(N__49890));
    SRMux I__11951 (
            .O(N__50348),
            .I(N__49890));
    SRMux I__11950 (
            .O(N__50347),
            .I(N__49890));
    SRMux I__11949 (
            .O(N__50346),
            .I(N__49890));
    SRMux I__11948 (
            .O(N__50345),
            .I(N__49890));
    SRMux I__11947 (
            .O(N__50344),
            .I(N__49890));
    SRMux I__11946 (
            .O(N__50343),
            .I(N__49890));
    SRMux I__11945 (
            .O(N__50342),
            .I(N__49890));
    SRMux I__11944 (
            .O(N__50341),
            .I(N__49890));
    SRMux I__11943 (
            .O(N__50340),
            .I(N__49890));
    SRMux I__11942 (
            .O(N__50339),
            .I(N__49890));
    SRMux I__11941 (
            .O(N__50338),
            .I(N__49890));
    SRMux I__11940 (
            .O(N__50337),
            .I(N__49890));
    SRMux I__11939 (
            .O(N__50336),
            .I(N__49890));
    SRMux I__11938 (
            .O(N__50335),
            .I(N__49890));
    SRMux I__11937 (
            .O(N__50334),
            .I(N__49890));
    SRMux I__11936 (
            .O(N__50333),
            .I(N__49890));
    SRMux I__11935 (
            .O(N__50332),
            .I(N__49890));
    SRMux I__11934 (
            .O(N__50331),
            .I(N__49890));
    SRMux I__11933 (
            .O(N__50330),
            .I(N__49890));
    SRMux I__11932 (
            .O(N__50329),
            .I(N__49890));
    SRMux I__11931 (
            .O(N__50328),
            .I(N__49890));
    SRMux I__11930 (
            .O(N__50327),
            .I(N__49890));
    SRMux I__11929 (
            .O(N__50326),
            .I(N__49890));
    SRMux I__11928 (
            .O(N__50325),
            .I(N__49890));
    SRMux I__11927 (
            .O(N__50324),
            .I(N__49890));
    SRMux I__11926 (
            .O(N__50323),
            .I(N__49890));
    SRMux I__11925 (
            .O(N__50322),
            .I(N__49890));
    SRMux I__11924 (
            .O(N__50321),
            .I(N__49890));
    SRMux I__11923 (
            .O(N__50320),
            .I(N__49890));
    SRMux I__11922 (
            .O(N__50319),
            .I(N__49890));
    SRMux I__11921 (
            .O(N__50318),
            .I(N__49890));
    SRMux I__11920 (
            .O(N__50317),
            .I(N__49890));
    SRMux I__11919 (
            .O(N__50316),
            .I(N__49890));
    SRMux I__11918 (
            .O(N__50315),
            .I(N__49890));
    SRMux I__11917 (
            .O(N__50314),
            .I(N__49890));
    SRMux I__11916 (
            .O(N__50313),
            .I(N__49890));
    SRMux I__11915 (
            .O(N__50312),
            .I(N__49890));
    SRMux I__11914 (
            .O(N__50311),
            .I(N__49890));
    SRMux I__11913 (
            .O(N__50310),
            .I(N__49890));
    SRMux I__11912 (
            .O(N__50309),
            .I(N__49890));
    SRMux I__11911 (
            .O(N__50308),
            .I(N__49890));
    SRMux I__11910 (
            .O(N__50307),
            .I(N__49890));
    SRMux I__11909 (
            .O(N__50306),
            .I(N__49890));
    SRMux I__11908 (
            .O(N__50305),
            .I(N__49890));
    SRMux I__11907 (
            .O(N__50304),
            .I(N__49890));
    SRMux I__11906 (
            .O(N__50303),
            .I(N__49890));
    SRMux I__11905 (
            .O(N__50302),
            .I(N__49890));
    SRMux I__11904 (
            .O(N__50301),
            .I(N__49890));
    SRMux I__11903 (
            .O(N__50300),
            .I(N__49890));
    SRMux I__11902 (
            .O(N__50299),
            .I(N__49890));
    SRMux I__11901 (
            .O(N__50298),
            .I(N__49890));
    SRMux I__11900 (
            .O(N__50297),
            .I(N__49890));
    SRMux I__11899 (
            .O(N__50296),
            .I(N__49890));
    SRMux I__11898 (
            .O(N__50295),
            .I(N__49890));
    SRMux I__11897 (
            .O(N__50294),
            .I(N__49890));
    SRMux I__11896 (
            .O(N__50293),
            .I(N__49890));
    SRMux I__11895 (
            .O(N__50292),
            .I(N__49890));
    SRMux I__11894 (
            .O(N__50291),
            .I(N__49890));
    SRMux I__11893 (
            .O(N__50290),
            .I(N__49890));
    SRMux I__11892 (
            .O(N__50289),
            .I(N__49890));
    SRMux I__11891 (
            .O(N__50288),
            .I(N__49890));
    SRMux I__11890 (
            .O(N__50287),
            .I(N__49890));
    SRMux I__11889 (
            .O(N__50286),
            .I(N__49890));
    SRMux I__11888 (
            .O(N__50285),
            .I(N__49890));
    SRMux I__11887 (
            .O(N__50284),
            .I(N__49890));
    SRMux I__11886 (
            .O(N__50283),
            .I(N__49890));
    SRMux I__11885 (
            .O(N__50282),
            .I(N__49890));
    SRMux I__11884 (
            .O(N__50281),
            .I(N__49890));
    SRMux I__11883 (
            .O(N__50280),
            .I(N__49890));
    SRMux I__11882 (
            .O(N__50279),
            .I(N__49890));
    SRMux I__11881 (
            .O(N__50278),
            .I(N__49890));
    SRMux I__11880 (
            .O(N__50277),
            .I(N__49890));
    SRMux I__11879 (
            .O(N__50276),
            .I(N__49890));
    SRMux I__11878 (
            .O(N__50275),
            .I(N__49890));
    SRMux I__11877 (
            .O(N__50274),
            .I(N__49890));
    SRMux I__11876 (
            .O(N__50273),
            .I(N__49890));
    SRMux I__11875 (
            .O(N__50272),
            .I(N__49890));
    SRMux I__11874 (
            .O(N__50271),
            .I(N__49890));
    SRMux I__11873 (
            .O(N__50270),
            .I(N__49890));
    SRMux I__11872 (
            .O(N__50269),
            .I(N__49890));
    SRMux I__11871 (
            .O(N__50268),
            .I(N__49890));
    SRMux I__11870 (
            .O(N__50267),
            .I(N__49890));
    SRMux I__11869 (
            .O(N__50266),
            .I(N__49890));
    SRMux I__11868 (
            .O(N__50265),
            .I(N__49890));
    SRMux I__11867 (
            .O(N__50264),
            .I(N__49890));
    SRMux I__11866 (
            .O(N__50263),
            .I(N__49890));
    SRMux I__11865 (
            .O(N__50262),
            .I(N__49890));
    SRMux I__11864 (
            .O(N__50261),
            .I(N__49890));
    SRMux I__11863 (
            .O(N__50260),
            .I(N__49890));
    SRMux I__11862 (
            .O(N__50259),
            .I(N__49890));
    SRMux I__11861 (
            .O(N__50258),
            .I(N__49890));
    SRMux I__11860 (
            .O(N__50257),
            .I(N__49890));
    SRMux I__11859 (
            .O(N__50256),
            .I(N__49890));
    SRMux I__11858 (
            .O(N__50255),
            .I(N__49890));
    SRMux I__11857 (
            .O(N__50254),
            .I(N__49890));
    SRMux I__11856 (
            .O(N__50253),
            .I(N__49890));
    SRMux I__11855 (
            .O(N__50252),
            .I(N__49890));
    SRMux I__11854 (
            .O(N__50251),
            .I(N__49890));
    SRMux I__11853 (
            .O(N__50250),
            .I(N__49890));
    SRMux I__11852 (
            .O(N__50249),
            .I(N__49890));
    SRMux I__11851 (
            .O(N__50248),
            .I(N__49890));
    SRMux I__11850 (
            .O(N__50247),
            .I(N__49890));
    SRMux I__11849 (
            .O(N__50246),
            .I(N__49890));
    SRMux I__11848 (
            .O(N__50245),
            .I(N__49890));
    SRMux I__11847 (
            .O(N__50244),
            .I(N__49890));
    SRMux I__11846 (
            .O(N__50243),
            .I(N__49890));
    SRMux I__11845 (
            .O(N__50242),
            .I(N__49890));
    SRMux I__11844 (
            .O(N__50241),
            .I(N__49890));
    SRMux I__11843 (
            .O(N__50240),
            .I(N__49890));
    SRMux I__11842 (
            .O(N__50239),
            .I(N__49890));
    SRMux I__11841 (
            .O(N__50238),
            .I(N__49890));
    SRMux I__11840 (
            .O(N__50237),
            .I(N__49890));
    SRMux I__11839 (
            .O(N__50236),
            .I(N__49890));
    SRMux I__11838 (
            .O(N__50235),
            .I(N__49890));
    SRMux I__11837 (
            .O(N__50234),
            .I(N__49890));
    SRMux I__11836 (
            .O(N__50233),
            .I(N__49890));
    SRMux I__11835 (
            .O(N__50232),
            .I(N__49890));
    SRMux I__11834 (
            .O(N__50231),
            .I(N__49890));
    SRMux I__11833 (
            .O(N__50230),
            .I(N__49890));
    SRMux I__11832 (
            .O(N__50229),
            .I(N__49890));
    GlobalMux I__11831 (
            .O(N__49890),
            .I(N__49887));
    gio2CtrlBuf I__11830 (
            .O(N__49887),
            .I(red_c_g));
    InMux I__11829 (
            .O(N__49884),
            .I(N__49879));
    InMux I__11828 (
            .O(N__49883),
            .I(N__49876));
    InMux I__11827 (
            .O(N__49882),
            .I(N__49873));
    LocalMux I__11826 (
            .O(N__49879),
            .I(N__49858));
    LocalMux I__11825 (
            .O(N__49876),
            .I(N__49858));
    LocalMux I__11824 (
            .O(N__49873),
            .I(N__49858));
    InMux I__11823 (
            .O(N__49872),
            .I(N__49855));
    InMux I__11822 (
            .O(N__49871),
            .I(N__49848));
    InMux I__11821 (
            .O(N__49870),
            .I(N__49848));
    InMux I__11820 (
            .O(N__49869),
            .I(N__49848));
    InMux I__11819 (
            .O(N__49868),
            .I(N__49839));
    InMux I__11818 (
            .O(N__49867),
            .I(N__49839));
    InMux I__11817 (
            .O(N__49866),
            .I(N__49839));
    InMux I__11816 (
            .O(N__49865),
            .I(N__49839));
    Span4Mux_s3_v I__11815 (
            .O(N__49858),
            .I(N__49830));
    LocalMux I__11814 (
            .O(N__49855),
            .I(N__49830));
    LocalMux I__11813 (
            .O(N__49848),
            .I(N__49830));
    LocalMux I__11812 (
            .O(N__49839),
            .I(N__49830));
    Span4Mux_v I__11811 (
            .O(N__49830),
            .I(N__49827));
    Span4Mux_v I__11810 (
            .O(N__49827),
            .I(N__49822));
    InMux I__11809 (
            .O(N__49826),
            .I(N__49819));
    InMux I__11808 (
            .O(N__49825),
            .I(N__49811));
    Span4Mux_v I__11807 (
            .O(N__49822),
            .I(N__49806));
    LocalMux I__11806 (
            .O(N__49819),
            .I(N__49806));
    InMux I__11805 (
            .O(N__49818),
            .I(N__49801));
    InMux I__11804 (
            .O(N__49817),
            .I(N__49801));
    InMux I__11803 (
            .O(N__49816),
            .I(N__49798));
    CascadeMux I__11802 (
            .O(N__49815),
            .I(N__49786));
    InMux I__11801 (
            .O(N__49814),
            .I(N__49766));
    LocalMux I__11800 (
            .O(N__49811),
            .I(N__49763));
    Span4Mux_v I__11799 (
            .O(N__49806),
            .I(N__49756));
    LocalMux I__11798 (
            .O(N__49801),
            .I(N__49756));
    LocalMux I__11797 (
            .O(N__49798),
            .I(N__49756));
    InMux I__11796 (
            .O(N__49797),
            .I(N__49753));
    InMux I__11795 (
            .O(N__49796),
            .I(N__49746));
    InMux I__11794 (
            .O(N__49795),
            .I(N__49746));
    InMux I__11793 (
            .O(N__49794),
            .I(N__49746));
    InMux I__11792 (
            .O(N__49793),
            .I(N__49737));
    InMux I__11791 (
            .O(N__49792),
            .I(N__49737));
    InMux I__11790 (
            .O(N__49791),
            .I(N__49737));
    InMux I__11789 (
            .O(N__49790),
            .I(N__49737));
    InMux I__11788 (
            .O(N__49789),
            .I(N__49730));
    InMux I__11787 (
            .O(N__49786),
            .I(N__49730));
    InMux I__11786 (
            .O(N__49785),
            .I(N__49730));
    InMux I__11785 (
            .O(N__49784),
            .I(N__49727));
    CascadeMux I__11784 (
            .O(N__49783),
            .I(N__49723));
    CascadeMux I__11783 (
            .O(N__49782),
            .I(N__49719));
    CascadeMux I__11782 (
            .O(N__49781),
            .I(N__49715));
    CascadeMux I__11781 (
            .O(N__49780),
            .I(N__49711));
    CascadeMux I__11780 (
            .O(N__49779),
            .I(N__49707));
    CascadeMux I__11779 (
            .O(N__49778),
            .I(N__49703));
    CascadeMux I__11778 (
            .O(N__49777),
            .I(N__49699));
    CascadeMux I__11777 (
            .O(N__49776),
            .I(N__49695));
    CascadeMux I__11776 (
            .O(N__49775),
            .I(N__49692));
    CascadeMux I__11775 (
            .O(N__49774),
            .I(N__49688));
    CascadeMux I__11774 (
            .O(N__49773),
            .I(N__49684));
    CascadeMux I__11773 (
            .O(N__49772),
            .I(N__49680));
    CascadeMux I__11772 (
            .O(N__49771),
            .I(N__49675));
    CascadeMux I__11771 (
            .O(N__49770),
            .I(N__49671));
    CascadeMux I__11770 (
            .O(N__49769),
            .I(N__49667));
    LocalMux I__11769 (
            .O(N__49766),
            .I(N__49661));
    Span4Mux_v I__11768 (
            .O(N__49763),
            .I(N__49661));
    Span4Mux_v I__11767 (
            .O(N__49756),
            .I(N__49649));
    LocalMux I__11766 (
            .O(N__49753),
            .I(N__49649));
    LocalMux I__11765 (
            .O(N__49746),
            .I(N__49649));
    LocalMux I__11764 (
            .O(N__49737),
            .I(N__49649));
    LocalMux I__11763 (
            .O(N__49730),
            .I(N__49646));
    LocalMux I__11762 (
            .O(N__49727),
            .I(N__49643));
    InMux I__11761 (
            .O(N__49726),
            .I(N__49640));
    InMux I__11760 (
            .O(N__49723),
            .I(N__49625));
    InMux I__11759 (
            .O(N__49722),
            .I(N__49625));
    InMux I__11758 (
            .O(N__49719),
            .I(N__49625));
    InMux I__11757 (
            .O(N__49718),
            .I(N__49625));
    InMux I__11756 (
            .O(N__49715),
            .I(N__49625));
    InMux I__11755 (
            .O(N__49714),
            .I(N__49625));
    InMux I__11754 (
            .O(N__49711),
            .I(N__49625));
    InMux I__11753 (
            .O(N__49710),
            .I(N__49608));
    InMux I__11752 (
            .O(N__49707),
            .I(N__49608));
    InMux I__11751 (
            .O(N__49706),
            .I(N__49608));
    InMux I__11750 (
            .O(N__49703),
            .I(N__49608));
    InMux I__11749 (
            .O(N__49702),
            .I(N__49608));
    InMux I__11748 (
            .O(N__49699),
            .I(N__49608));
    InMux I__11747 (
            .O(N__49698),
            .I(N__49608));
    InMux I__11746 (
            .O(N__49695),
            .I(N__49608));
    InMux I__11745 (
            .O(N__49692),
            .I(N__49591));
    InMux I__11744 (
            .O(N__49691),
            .I(N__49591));
    InMux I__11743 (
            .O(N__49688),
            .I(N__49591));
    InMux I__11742 (
            .O(N__49687),
            .I(N__49591));
    InMux I__11741 (
            .O(N__49684),
            .I(N__49591));
    InMux I__11740 (
            .O(N__49683),
            .I(N__49591));
    InMux I__11739 (
            .O(N__49680),
            .I(N__49591));
    InMux I__11738 (
            .O(N__49679),
            .I(N__49591));
    InMux I__11737 (
            .O(N__49678),
            .I(N__49576));
    InMux I__11736 (
            .O(N__49675),
            .I(N__49576));
    InMux I__11735 (
            .O(N__49674),
            .I(N__49576));
    InMux I__11734 (
            .O(N__49671),
            .I(N__49576));
    InMux I__11733 (
            .O(N__49670),
            .I(N__49576));
    InMux I__11732 (
            .O(N__49667),
            .I(N__49576));
    InMux I__11731 (
            .O(N__49666),
            .I(N__49576));
    IoSpan4Mux I__11730 (
            .O(N__49661),
            .I(N__49573));
    InMux I__11729 (
            .O(N__49660),
            .I(N__49568));
    InMux I__11728 (
            .O(N__49659),
            .I(N__49568));
    InMux I__11727 (
            .O(N__49658),
            .I(N__49565));
    Span4Mux_v I__11726 (
            .O(N__49649),
            .I(N__49562));
    Span4Mux_v I__11725 (
            .O(N__49646),
            .I(N__49559));
    Span4Mux_v I__11724 (
            .O(N__49643),
            .I(N__49554));
    LocalMux I__11723 (
            .O(N__49640),
            .I(N__49554));
    LocalMux I__11722 (
            .O(N__49625),
            .I(N__49545));
    LocalMux I__11721 (
            .O(N__49608),
            .I(N__49545));
    LocalMux I__11720 (
            .O(N__49591),
            .I(N__49545));
    LocalMux I__11719 (
            .O(N__49576),
            .I(N__49545));
    Span4Mux_s0_v I__11718 (
            .O(N__49573),
            .I(N__49542));
    LocalMux I__11717 (
            .O(N__49568),
            .I(N__49537));
    LocalMux I__11716 (
            .O(N__49565),
            .I(N__49537));
    Sp12to4 I__11715 (
            .O(N__49562),
            .I(N__49534));
    Sp12to4 I__11714 (
            .O(N__49559),
            .I(N__49531));
    Span4Mux_h I__11713 (
            .O(N__49554),
            .I(N__49526));
    Span4Mux_v I__11712 (
            .O(N__49545),
            .I(N__49526));
    Span4Mux_v I__11711 (
            .O(N__49542),
            .I(N__49523));
    Span4Mux_s3_h I__11710 (
            .O(N__49537),
            .I(N__49520));
    Span12Mux_s10_h I__11709 (
            .O(N__49534),
            .I(N__49517));
    Span12Mux_s10_h I__11708 (
            .O(N__49531),
            .I(N__49512));
    Sp12to4 I__11707 (
            .O(N__49526),
            .I(N__49512));
    Sp12to4 I__11706 (
            .O(N__49523),
            .I(N__49507));
    Sp12to4 I__11705 (
            .O(N__49520),
            .I(N__49507));
    Span12Mux_h I__11704 (
            .O(N__49517),
            .I(N__49500));
    Span12Mux_h I__11703 (
            .O(N__49512),
            .I(N__49500));
    Span12Mux_v I__11702 (
            .O(N__49507),
            .I(N__49500));
    Odrv12 I__11701 (
            .O(N__49500),
            .I(CONSTANT_ONE_NET));
    InMux I__11700 (
            .O(N__49497),
            .I(N__49493));
    InMux I__11699 (
            .O(N__49496),
            .I(N__49489));
    LocalMux I__11698 (
            .O(N__49493),
            .I(N__49486));
    InMux I__11697 (
            .O(N__49492),
            .I(N__49483));
    LocalMux I__11696 (
            .O(N__49489),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    Odrv4 I__11695 (
            .O(N__49486),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    LocalMux I__11694 (
            .O(N__49483),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    InMux I__11693 (
            .O(N__49476),
            .I(N__49470));
    InMux I__11692 (
            .O(N__49475),
            .I(N__49467));
    InMux I__11691 (
            .O(N__49474),
            .I(N__49464));
    InMux I__11690 (
            .O(N__49473),
            .I(N__49461));
    LocalMux I__11689 (
            .O(N__49470),
            .I(N__49458));
    LocalMux I__11688 (
            .O(N__49467),
            .I(N__49453));
    LocalMux I__11687 (
            .O(N__49464),
            .I(N__49453));
    LocalMux I__11686 (
            .O(N__49461),
            .I(N__49450));
    Span4Mux_v I__11685 (
            .O(N__49458),
            .I(N__49443));
    Span4Mux_v I__11684 (
            .O(N__49453),
            .I(N__49443));
    Span4Mux_v I__11683 (
            .O(N__49450),
            .I(N__49443));
    Odrv4 I__11682 (
            .O(N__49443),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    CascadeMux I__11681 (
            .O(N__49440),
            .I(N__49436));
    InMux I__11680 (
            .O(N__49439),
            .I(N__49431));
    InMux I__11679 (
            .O(N__49436),
            .I(N__49431));
    LocalMux I__11678 (
            .O(N__49431),
            .I(N__49428));
    Odrv4 I__11677 (
            .O(N__49428),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__11676 (
            .O(N__49425),
            .I(N__49422));
    InMux I__11675 (
            .O(N__49422),
            .I(N__49416));
    InMux I__11674 (
            .O(N__49421),
            .I(N__49413));
    InMux I__11673 (
            .O(N__49420),
            .I(N__49410));
    InMux I__11672 (
            .O(N__49419),
            .I(N__49407));
    LocalMux I__11671 (
            .O(N__49416),
            .I(N__49404));
    LocalMux I__11670 (
            .O(N__49413),
            .I(N__49401));
    LocalMux I__11669 (
            .O(N__49410),
            .I(N__49396));
    LocalMux I__11668 (
            .O(N__49407),
            .I(N__49396));
    Span4Mux_h I__11667 (
            .O(N__49404),
            .I(N__49393));
    Span4Mux_v I__11666 (
            .O(N__49401),
            .I(N__49390));
    Span4Mux_v I__11665 (
            .O(N__49396),
            .I(N__49385));
    Span4Mux_v I__11664 (
            .O(N__49393),
            .I(N__49385));
    Odrv4 I__11663 (
            .O(N__49390),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    Odrv4 I__11662 (
            .O(N__49385),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__11661 (
            .O(N__49380),
            .I(N__49377));
    LocalMux I__11660 (
            .O(N__49377),
            .I(N__49374));
    Span4Mux_h I__11659 (
            .O(N__49374),
            .I(N__49369));
    InMux I__11658 (
            .O(N__49373),
            .I(N__49366));
    InMux I__11657 (
            .O(N__49372),
            .I(N__49363));
    Span4Mux_v I__11656 (
            .O(N__49369),
            .I(N__49360));
    LocalMux I__11655 (
            .O(N__49366),
            .I(N__49357));
    LocalMux I__11654 (
            .O(N__49363),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__11653 (
            .O(N__49360),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__11652 (
            .O(N__49357),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__11651 (
            .O(N__49350),
            .I(N__49347));
    LocalMux I__11650 (
            .O(N__49347),
            .I(N__49344));
    Odrv4 I__11649 (
            .O(N__49344),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ));
    CascadeMux I__11648 (
            .O(N__49341),
            .I(N__49338));
    InMux I__11647 (
            .O(N__49338),
            .I(N__49332));
    InMux I__11646 (
            .O(N__49337),
            .I(N__49332));
    LocalMux I__11645 (
            .O(N__49332),
            .I(N__49329));
    Span4Mux_h I__11644 (
            .O(N__49329),
            .I(N__49326));
    Odrv4 I__11643 (
            .O(N__49326),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ));
    InMux I__11642 (
            .O(N__49323),
            .I(N__49319));
    InMux I__11641 (
            .O(N__49322),
            .I(N__49315));
    LocalMux I__11640 (
            .O(N__49319),
            .I(N__49312));
    InMux I__11639 (
            .O(N__49318),
            .I(N__49309));
    LocalMux I__11638 (
            .O(N__49315),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    Odrv12 I__11637 (
            .O(N__49312),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    LocalMux I__11636 (
            .O(N__49309),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    InMux I__11635 (
            .O(N__49302),
            .I(N__49298));
    InMux I__11634 (
            .O(N__49301),
            .I(N__49293));
    LocalMux I__11633 (
            .O(N__49298),
            .I(N__49290));
    InMux I__11632 (
            .O(N__49297),
            .I(N__49285));
    InMux I__11631 (
            .O(N__49296),
            .I(N__49285));
    LocalMux I__11630 (
            .O(N__49293),
            .I(N__49282));
    Span4Mux_h I__11629 (
            .O(N__49290),
            .I(N__49279));
    LocalMux I__11628 (
            .O(N__49285),
            .I(N__49276));
    Span4Mux_h I__11627 (
            .O(N__49282),
            .I(N__49271));
    Span4Mux_v I__11626 (
            .O(N__49279),
            .I(N__49271));
    Span4Mux_h I__11625 (
            .O(N__49276),
            .I(N__49268));
    Odrv4 I__11624 (
            .O(N__49271),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    Odrv4 I__11623 (
            .O(N__49268),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__11622 (
            .O(N__49263),
            .I(N__49260));
    LocalMux I__11621 (
            .O(N__49260),
            .I(N__49257));
    Span4Mux_h I__11620 (
            .O(N__49257),
            .I(N__49254));
    Odrv4 I__11619 (
            .O(N__49254),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ));
    CEMux I__11618 (
            .O(N__49251),
            .I(N__49212));
    CEMux I__11617 (
            .O(N__49250),
            .I(N__49212));
    CEMux I__11616 (
            .O(N__49249),
            .I(N__49212));
    CEMux I__11615 (
            .O(N__49248),
            .I(N__49212));
    CEMux I__11614 (
            .O(N__49247),
            .I(N__49212));
    CEMux I__11613 (
            .O(N__49246),
            .I(N__49212));
    CEMux I__11612 (
            .O(N__49245),
            .I(N__49212));
    CEMux I__11611 (
            .O(N__49244),
            .I(N__49212));
    CEMux I__11610 (
            .O(N__49243),
            .I(N__49212));
    CEMux I__11609 (
            .O(N__49242),
            .I(N__49212));
    CEMux I__11608 (
            .O(N__49241),
            .I(N__49212));
    CEMux I__11607 (
            .O(N__49240),
            .I(N__49212));
    CEMux I__11606 (
            .O(N__49239),
            .I(N__49212));
    GlobalMux I__11605 (
            .O(N__49212),
            .I(N__49209));
    gio2CtrlBuf I__11604 (
            .O(N__49209),
            .I(\phase_controller_inst2.stoper_hc.un1_start_g ));
    InMux I__11603 (
            .O(N__49206),
            .I(N__49202));
    InMux I__11602 (
            .O(N__49205),
            .I(N__49197));
    LocalMux I__11601 (
            .O(N__49202),
            .I(N__49194));
    InMux I__11600 (
            .O(N__49201),
            .I(N__49189));
    InMux I__11599 (
            .O(N__49200),
            .I(N__49189));
    LocalMux I__11598 (
            .O(N__49197),
            .I(N__49186));
    Span4Mux_v I__11597 (
            .O(N__49194),
            .I(N__49183));
    LocalMux I__11596 (
            .O(N__49189),
            .I(N__49180));
    Span4Mux_v I__11595 (
            .O(N__49186),
            .I(N__49177));
    Span4Mux_v I__11594 (
            .O(N__49183),
            .I(N__49174));
    Span4Mux_h I__11593 (
            .O(N__49180),
            .I(N__49171));
    Odrv4 I__11592 (
            .O(N__49177),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__11591 (
            .O(N__49174),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__11590 (
            .O(N__49171),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    InMux I__11589 (
            .O(N__49164),
            .I(N__49161));
    LocalMux I__11588 (
            .O(N__49161),
            .I(N__49158));
    Span4Mux_v I__11587 (
            .O(N__49158),
            .I(N__49155));
    Span4Mux_v I__11586 (
            .O(N__49155),
            .I(N__49150));
    InMux I__11585 (
            .O(N__49154),
            .I(N__49147));
    InMux I__11584 (
            .O(N__49153),
            .I(N__49144));
    Span4Mux_h I__11583 (
            .O(N__49150),
            .I(N__49141));
    LocalMux I__11582 (
            .O(N__49147),
            .I(N__49138));
    LocalMux I__11581 (
            .O(N__49144),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__11580 (
            .O(N__49141),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv4 I__11579 (
            .O(N__49138),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__11578 (
            .O(N__49131),
            .I(N__49127));
    InMux I__11577 (
            .O(N__49130),
            .I(N__49124));
    LocalMux I__11576 (
            .O(N__49127),
            .I(N__49121));
    LocalMux I__11575 (
            .O(N__49124),
            .I(N__49116));
    Span4Mux_v I__11574 (
            .O(N__49121),
            .I(N__49113));
    InMux I__11573 (
            .O(N__49120),
            .I(N__49110));
    InMux I__11572 (
            .O(N__49119),
            .I(N__49107));
    Span4Mux_v I__11571 (
            .O(N__49116),
            .I(N__49100));
    Span4Mux_h I__11570 (
            .O(N__49113),
            .I(N__49100));
    LocalMux I__11569 (
            .O(N__49110),
            .I(N__49100));
    LocalMux I__11568 (
            .O(N__49107),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__11567 (
            .O(N__49100),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__11566 (
            .O(N__49095),
            .I(N__49069));
    InMux I__11565 (
            .O(N__49094),
            .I(N__49069));
    InMux I__11564 (
            .O(N__49093),
            .I(N__49060));
    InMux I__11563 (
            .O(N__49092),
            .I(N__49060));
    InMux I__11562 (
            .O(N__49091),
            .I(N__49060));
    InMux I__11561 (
            .O(N__49090),
            .I(N__49060));
    InMux I__11560 (
            .O(N__49089),
            .I(N__49051));
    InMux I__11559 (
            .O(N__49088),
            .I(N__49051));
    InMux I__11558 (
            .O(N__49087),
            .I(N__49051));
    InMux I__11557 (
            .O(N__49086),
            .I(N__49051));
    InMux I__11556 (
            .O(N__49085),
            .I(N__49042));
    InMux I__11555 (
            .O(N__49084),
            .I(N__49042));
    InMux I__11554 (
            .O(N__49083),
            .I(N__49042));
    InMux I__11553 (
            .O(N__49082),
            .I(N__49042));
    InMux I__11552 (
            .O(N__49081),
            .I(N__49033));
    InMux I__11551 (
            .O(N__49080),
            .I(N__49033));
    InMux I__11550 (
            .O(N__49079),
            .I(N__49033));
    InMux I__11549 (
            .O(N__49078),
            .I(N__49033));
    InMux I__11548 (
            .O(N__49077),
            .I(N__49016));
    InMux I__11547 (
            .O(N__49076),
            .I(N__49016));
    InMux I__11546 (
            .O(N__49075),
            .I(N__49016));
    InMux I__11545 (
            .O(N__49074),
            .I(N__49016));
    LocalMux I__11544 (
            .O(N__49069),
            .I(N__49005));
    LocalMux I__11543 (
            .O(N__49060),
            .I(N__49005));
    LocalMux I__11542 (
            .O(N__49051),
            .I(N__49005));
    LocalMux I__11541 (
            .O(N__49042),
            .I(N__49005));
    LocalMux I__11540 (
            .O(N__49033),
            .I(N__49005));
    InMux I__11539 (
            .O(N__49032),
            .I(N__48996));
    InMux I__11538 (
            .O(N__49031),
            .I(N__48996));
    InMux I__11537 (
            .O(N__49030),
            .I(N__48996));
    InMux I__11536 (
            .O(N__49029),
            .I(N__48996));
    InMux I__11535 (
            .O(N__49028),
            .I(N__48987));
    InMux I__11534 (
            .O(N__49027),
            .I(N__48987));
    InMux I__11533 (
            .O(N__49026),
            .I(N__48987));
    InMux I__11532 (
            .O(N__49025),
            .I(N__48987));
    LocalMux I__11531 (
            .O(N__49016),
            .I(N__48980));
    Span4Mux_v I__11530 (
            .O(N__49005),
            .I(N__48980));
    LocalMux I__11529 (
            .O(N__48996),
            .I(N__48980));
    LocalMux I__11528 (
            .O(N__48987),
            .I(N__48977));
    Span4Mux_h I__11527 (
            .O(N__48980),
            .I(N__48974));
    Span4Mux_h I__11526 (
            .O(N__48977),
            .I(N__48971));
    Span4Mux_v I__11525 (
            .O(N__48974),
            .I(N__48968));
    Odrv4 I__11524 (
            .O(N__48971),
            .I(\current_shift_inst.timer_s1.running_i ));
    Odrv4 I__11523 (
            .O(N__48968),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__11522 (
            .O(N__48963),
            .I(N__48958));
    InMux I__11521 (
            .O(N__48962),
            .I(N__48955));
    InMux I__11520 (
            .O(N__48961),
            .I(N__48952));
    LocalMux I__11519 (
            .O(N__48958),
            .I(N__48949));
    LocalMux I__11518 (
            .O(N__48955),
            .I(N__48946));
    LocalMux I__11517 (
            .O(N__48952),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv12 I__11516 (
            .O(N__48949),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    Odrv4 I__11515 (
            .O(N__48946),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    CascadeMux I__11514 (
            .O(N__48939),
            .I(N__48933));
    InMux I__11513 (
            .O(N__48938),
            .I(N__48930));
    InMux I__11512 (
            .O(N__48937),
            .I(N__48927));
    InMux I__11511 (
            .O(N__48936),
            .I(N__48924));
    InMux I__11510 (
            .O(N__48933),
            .I(N__48921));
    LocalMux I__11509 (
            .O(N__48930),
            .I(N__48918));
    LocalMux I__11508 (
            .O(N__48927),
            .I(N__48915));
    LocalMux I__11507 (
            .O(N__48924),
            .I(N__48912));
    LocalMux I__11506 (
            .O(N__48921),
            .I(N__48909));
    Span4Mux_v I__11505 (
            .O(N__48918),
            .I(N__48902));
    Span4Mux_v I__11504 (
            .O(N__48915),
            .I(N__48902));
    Span4Mux_v I__11503 (
            .O(N__48912),
            .I(N__48902));
    Span4Mux_h I__11502 (
            .O(N__48909),
            .I(N__48899));
    Odrv4 I__11501 (
            .O(N__48902),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    Odrv4 I__11500 (
            .O(N__48899),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    CascadeMux I__11499 (
            .O(N__48894),
            .I(N__48890));
    CascadeMux I__11498 (
            .O(N__48893),
            .I(N__48887));
    InMux I__11497 (
            .O(N__48890),
            .I(N__48882));
    InMux I__11496 (
            .O(N__48887),
            .I(N__48882));
    LocalMux I__11495 (
            .O(N__48882),
            .I(N__48879));
    Odrv12 I__11494 (
            .O(N__48879),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ));
    CEMux I__11493 (
            .O(N__48876),
            .I(N__48872));
    CEMux I__11492 (
            .O(N__48875),
            .I(N__48869));
    LocalMux I__11491 (
            .O(N__48872),
            .I(N__48863));
    LocalMux I__11490 (
            .O(N__48869),
            .I(N__48857));
    CEMux I__11489 (
            .O(N__48868),
            .I(N__48854));
    CEMux I__11488 (
            .O(N__48867),
            .I(N__48848));
    CEMux I__11487 (
            .O(N__48866),
            .I(N__48845));
    Span4Mux_h I__11486 (
            .O(N__48863),
            .I(N__48830));
    CEMux I__11485 (
            .O(N__48862),
            .I(N__48827));
    CEMux I__11484 (
            .O(N__48861),
            .I(N__48821));
    CEMux I__11483 (
            .O(N__48860),
            .I(N__48818));
    Span4Mux_v I__11482 (
            .O(N__48857),
            .I(N__48813));
    LocalMux I__11481 (
            .O(N__48854),
            .I(N__48813));
    CEMux I__11480 (
            .O(N__48853),
            .I(N__48806));
    CEMux I__11479 (
            .O(N__48852),
            .I(N__48803));
    CEMux I__11478 (
            .O(N__48851),
            .I(N__48800));
    LocalMux I__11477 (
            .O(N__48848),
            .I(N__48797));
    LocalMux I__11476 (
            .O(N__48845),
            .I(N__48794));
    InMux I__11475 (
            .O(N__48844),
            .I(N__48787));
    InMux I__11474 (
            .O(N__48843),
            .I(N__48787));
    InMux I__11473 (
            .O(N__48842),
            .I(N__48787));
    InMux I__11472 (
            .O(N__48841),
            .I(N__48778));
    InMux I__11471 (
            .O(N__48840),
            .I(N__48778));
    InMux I__11470 (
            .O(N__48839),
            .I(N__48778));
    InMux I__11469 (
            .O(N__48838),
            .I(N__48778));
    CEMux I__11468 (
            .O(N__48837),
            .I(N__48775));
    InMux I__11467 (
            .O(N__48836),
            .I(N__48766));
    InMux I__11466 (
            .O(N__48835),
            .I(N__48766));
    InMux I__11465 (
            .O(N__48834),
            .I(N__48766));
    InMux I__11464 (
            .O(N__48833),
            .I(N__48766));
    Span4Mux_h I__11463 (
            .O(N__48830),
            .I(N__48761));
    LocalMux I__11462 (
            .O(N__48827),
            .I(N__48761));
    CEMux I__11461 (
            .O(N__48826),
            .I(N__48758));
    CEMux I__11460 (
            .O(N__48825),
            .I(N__48755));
    CEMux I__11459 (
            .O(N__48824),
            .I(N__48748));
    LocalMux I__11458 (
            .O(N__48821),
            .I(N__48745));
    LocalMux I__11457 (
            .O(N__48818),
            .I(N__48742));
    Span4Mux_v I__11456 (
            .O(N__48813),
            .I(N__48739));
    CEMux I__11455 (
            .O(N__48812),
            .I(N__48736));
    InMux I__11454 (
            .O(N__48811),
            .I(N__48729));
    InMux I__11453 (
            .O(N__48810),
            .I(N__48729));
    InMux I__11452 (
            .O(N__48809),
            .I(N__48729));
    LocalMux I__11451 (
            .O(N__48806),
            .I(N__48724));
    LocalMux I__11450 (
            .O(N__48803),
            .I(N__48724));
    LocalMux I__11449 (
            .O(N__48800),
            .I(N__48708));
    Span4Mux_h I__11448 (
            .O(N__48797),
            .I(N__48693));
    Span4Mux_h I__11447 (
            .O(N__48794),
            .I(N__48693));
    LocalMux I__11446 (
            .O(N__48787),
            .I(N__48693));
    LocalMux I__11445 (
            .O(N__48778),
            .I(N__48693));
    LocalMux I__11444 (
            .O(N__48775),
            .I(N__48693));
    LocalMux I__11443 (
            .O(N__48766),
            .I(N__48693));
    Span4Mux_h I__11442 (
            .O(N__48761),
            .I(N__48693));
    LocalMux I__11441 (
            .O(N__48758),
            .I(N__48690));
    LocalMux I__11440 (
            .O(N__48755),
            .I(N__48687));
    InMux I__11439 (
            .O(N__48754),
            .I(N__48678));
    InMux I__11438 (
            .O(N__48753),
            .I(N__48678));
    InMux I__11437 (
            .O(N__48752),
            .I(N__48678));
    InMux I__11436 (
            .O(N__48751),
            .I(N__48678));
    LocalMux I__11435 (
            .O(N__48748),
            .I(N__48669));
    Span4Mux_v I__11434 (
            .O(N__48745),
            .I(N__48669));
    Span4Mux_h I__11433 (
            .O(N__48742),
            .I(N__48669));
    Span4Mux_h I__11432 (
            .O(N__48739),
            .I(N__48669));
    LocalMux I__11431 (
            .O(N__48736),
            .I(N__48666));
    LocalMux I__11430 (
            .O(N__48729),
            .I(N__48661));
    Span4Mux_v I__11429 (
            .O(N__48724),
            .I(N__48661));
    InMux I__11428 (
            .O(N__48723),
            .I(N__48652));
    InMux I__11427 (
            .O(N__48722),
            .I(N__48652));
    InMux I__11426 (
            .O(N__48721),
            .I(N__48652));
    InMux I__11425 (
            .O(N__48720),
            .I(N__48652));
    InMux I__11424 (
            .O(N__48719),
            .I(N__48643));
    InMux I__11423 (
            .O(N__48718),
            .I(N__48643));
    InMux I__11422 (
            .O(N__48717),
            .I(N__48643));
    InMux I__11421 (
            .O(N__48716),
            .I(N__48643));
    InMux I__11420 (
            .O(N__48715),
            .I(N__48634));
    InMux I__11419 (
            .O(N__48714),
            .I(N__48634));
    InMux I__11418 (
            .O(N__48713),
            .I(N__48634));
    InMux I__11417 (
            .O(N__48712),
            .I(N__48634));
    InMux I__11416 (
            .O(N__48711),
            .I(N__48631));
    Sp12to4 I__11415 (
            .O(N__48708),
            .I(N__48628));
    Span4Mux_v I__11414 (
            .O(N__48693),
            .I(N__48625));
    Span4Mux_h I__11413 (
            .O(N__48690),
            .I(N__48616));
    Span4Mux_v I__11412 (
            .O(N__48687),
            .I(N__48616));
    LocalMux I__11411 (
            .O(N__48678),
            .I(N__48616));
    Span4Mux_h I__11410 (
            .O(N__48669),
            .I(N__48616));
    Odrv4 I__11409 (
            .O(N__48666),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11408 (
            .O(N__48661),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__11407 (
            .O(N__48652),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__11406 (
            .O(N__48643),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__11405 (
            .O(N__48634),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    LocalMux I__11404 (
            .O(N__48631),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv12 I__11403 (
            .O(N__48628),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11402 (
            .O(N__48625),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    Odrv4 I__11401 (
            .O(N__48616),
            .I(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ));
    InMux I__11400 (
            .O(N__48597),
            .I(N__48594));
    LocalMux I__11399 (
            .O(N__48594),
            .I(N__48589));
    InMux I__11398 (
            .O(N__48593),
            .I(N__48586));
    InMux I__11397 (
            .O(N__48592),
            .I(N__48583));
    Span4Mux_h I__11396 (
            .O(N__48589),
            .I(N__48578));
    LocalMux I__11395 (
            .O(N__48586),
            .I(N__48578));
    LocalMux I__11394 (
            .O(N__48583),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    Odrv4 I__11393 (
            .O(N__48578),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    InMux I__11392 (
            .O(N__48573),
            .I(N__48568));
    InMux I__11391 (
            .O(N__48572),
            .I(N__48562));
    InMux I__11390 (
            .O(N__48571),
            .I(N__48562));
    LocalMux I__11389 (
            .O(N__48568),
            .I(N__48559));
    InMux I__11388 (
            .O(N__48567),
            .I(N__48556));
    LocalMux I__11387 (
            .O(N__48562),
            .I(N__48553));
    Span4Mux_h I__11386 (
            .O(N__48559),
            .I(N__48550));
    LocalMux I__11385 (
            .O(N__48556),
            .I(N__48547));
    Span4Mux_h I__11384 (
            .O(N__48553),
            .I(N__48544));
    Odrv4 I__11383 (
            .O(N__48550),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__11382 (
            .O(N__48547),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__11381 (
            .O(N__48544),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__11380 (
            .O(N__48537),
            .I(N__48534));
    LocalMux I__11379 (
            .O(N__48534),
            .I(N__48531));
    Span4Mux_v I__11378 (
            .O(N__48531),
            .I(N__48528));
    Odrv4 I__11377 (
            .O(N__48528),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ));
    InMux I__11376 (
            .O(N__48525),
            .I(N__48520));
    InMux I__11375 (
            .O(N__48524),
            .I(N__48517));
    InMux I__11374 (
            .O(N__48523),
            .I(N__48514));
    LocalMux I__11373 (
            .O(N__48520),
            .I(N__48511));
    LocalMux I__11372 (
            .O(N__48517),
            .I(N__48508));
    LocalMux I__11371 (
            .O(N__48514),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv12 I__11370 (
            .O(N__48511),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__11369 (
            .O(N__48508),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__11368 (
            .O(N__48501),
            .I(N__48497));
    InMux I__11367 (
            .O(N__48500),
            .I(N__48494));
    LocalMux I__11366 (
            .O(N__48497),
            .I(N__48489));
    LocalMux I__11365 (
            .O(N__48494),
            .I(N__48486));
    InMux I__11364 (
            .O(N__48493),
            .I(N__48483));
    InMux I__11363 (
            .O(N__48492),
            .I(N__48480));
    Odrv12 I__11362 (
            .O(N__48489),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    Odrv4 I__11361 (
            .O(N__48486),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__11360 (
            .O(N__48483),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__11359 (
            .O(N__48480),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__11358 (
            .O(N__48471),
            .I(N__48468));
    LocalMux I__11357 (
            .O(N__48468),
            .I(N__48465));
    Span4Mux_v I__11356 (
            .O(N__48465),
            .I(N__48462));
    Odrv4 I__11355 (
            .O(N__48462),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ));
    InMux I__11354 (
            .O(N__48459),
            .I(N__48456));
    LocalMux I__11353 (
            .O(N__48456),
            .I(N__48451));
    InMux I__11352 (
            .O(N__48455),
            .I(N__48448));
    InMux I__11351 (
            .O(N__48454),
            .I(N__48445));
    Span4Mux_h I__11350 (
            .O(N__48451),
            .I(N__48442));
    LocalMux I__11349 (
            .O(N__48448),
            .I(N__48439));
    LocalMux I__11348 (
            .O(N__48445),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv4 I__11347 (
            .O(N__48442),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    Odrv12 I__11346 (
            .O(N__48439),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__11345 (
            .O(N__48432),
            .I(N__48426));
    InMux I__11344 (
            .O(N__48431),
            .I(N__48421));
    InMux I__11343 (
            .O(N__48430),
            .I(N__48421));
    InMux I__11342 (
            .O(N__48429),
            .I(N__48418));
    LocalMux I__11341 (
            .O(N__48426),
            .I(N__48415));
    LocalMux I__11340 (
            .O(N__48421),
            .I(N__48412));
    LocalMux I__11339 (
            .O(N__48418),
            .I(N__48409));
    Span4Mux_v I__11338 (
            .O(N__48415),
            .I(N__48404));
    Span4Mux_v I__11337 (
            .O(N__48412),
            .I(N__48404));
    Odrv12 I__11336 (
            .O(N__48409),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    Odrv4 I__11335 (
            .O(N__48404),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    CascadeMux I__11334 (
            .O(N__48399),
            .I(N__48396));
    InMux I__11333 (
            .O(N__48396),
            .I(N__48393));
    LocalMux I__11332 (
            .O(N__48393),
            .I(N__48390));
    Span4Mux_v I__11331 (
            .O(N__48390),
            .I(N__48387));
    Odrv4 I__11330 (
            .O(N__48387),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ));
    CascadeMux I__11329 (
            .O(N__48384),
            .I(N__48378));
    InMux I__11328 (
            .O(N__48383),
            .I(N__48373));
    InMux I__11327 (
            .O(N__48382),
            .I(N__48373));
    InMux I__11326 (
            .O(N__48381),
            .I(N__48370));
    InMux I__11325 (
            .O(N__48378),
            .I(N__48367));
    LocalMux I__11324 (
            .O(N__48373),
            .I(N__48364));
    LocalMux I__11323 (
            .O(N__48370),
            .I(N__48361));
    LocalMux I__11322 (
            .O(N__48367),
            .I(N__48358));
    Span4Mux_h I__11321 (
            .O(N__48364),
            .I(N__48355));
    Span4Mux_h I__11320 (
            .O(N__48361),
            .I(N__48350));
    Span4Mux_h I__11319 (
            .O(N__48358),
            .I(N__48350));
    Odrv4 I__11318 (
            .O(N__48355),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    Odrv4 I__11317 (
            .O(N__48350),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__11316 (
            .O(N__48345),
            .I(N__48342));
    LocalMux I__11315 (
            .O(N__48342),
            .I(N__48339));
    Span4Mux_v I__11314 (
            .O(N__48339),
            .I(N__48335));
    InMux I__11313 (
            .O(N__48338),
            .I(N__48332));
    Odrv4 I__11312 (
            .O(N__48335),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    LocalMux I__11311 (
            .O(N__48332),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    CascadeMux I__11310 (
            .O(N__48327),
            .I(N__48324));
    InMux I__11309 (
            .O(N__48324),
            .I(N__48321));
    LocalMux I__11308 (
            .O(N__48321),
            .I(N__48318));
    Span12Mux_v I__11307 (
            .O(N__48318),
            .I(N__48315));
    Odrv12 I__11306 (
            .O(N__48315),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ));
    InMux I__11305 (
            .O(N__48312),
            .I(N__48309));
    LocalMux I__11304 (
            .O(N__48309),
            .I(N__48304));
    InMux I__11303 (
            .O(N__48308),
            .I(N__48301));
    InMux I__11302 (
            .O(N__48307),
            .I(N__48298));
    Span4Mux_v I__11301 (
            .O(N__48304),
            .I(N__48295));
    LocalMux I__11300 (
            .O(N__48301),
            .I(N__48292));
    LocalMux I__11299 (
            .O(N__48298),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv4 I__11298 (
            .O(N__48295),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    Odrv12 I__11297 (
            .O(N__48292),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    InMux I__11296 (
            .O(N__48285),
            .I(N__48279));
    InMux I__11295 (
            .O(N__48284),
            .I(N__48276));
    InMux I__11294 (
            .O(N__48283),
            .I(N__48273));
    InMux I__11293 (
            .O(N__48282),
            .I(N__48270));
    LocalMux I__11292 (
            .O(N__48279),
            .I(N__48267));
    LocalMux I__11291 (
            .O(N__48276),
            .I(N__48264));
    LocalMux I__11290 (
            .O(N__48273),
            .I(N__48261));
    LocalMux I__11289 (
            .O(N__48270),
            .I(N__48258));
    Span4Mux_v I__11288 (
            .O(N__48267),
            .I(N__48249));
    Span4Mux_v I__11287 (
            .O(N__48264),
            .I(N__48249));
    Span4Mux_v I__11286 (
            .O(N__48261),
            .I(N__48249));
    Span4Mux_v I__11285 (
            .O(N__48258),
            .I(N__48249));
    Odrv4 I__11284 (
            .O(N__48249),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    CascadeMux I__11283 (
            .O(N__48246),
            .I(N__48243));
    InMux I__11282 (
            .O(N__48243),
            .I(N__48240));
    LocalMux I__11281 (
            .O(N__48240),
            .I(N__48237));
    Span4Mux_v I__11280 (
            .O(N__48237),
            .I(N__48234));
    Odrv4 I__11279 (
            .O(N__48234),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ));
    InMux I__11278 (
            .O(N__48231),
            .I(N__48228));
    LocalMux I__11277 (
            .O(N__48228),
            .I(N__48225));
    Span4Mux_h I__11276 (
            .O(N__48225),
            .I(N__48222));
    Span4Mux_v I__11275 (
            .O(N__48222),
            .I(N__48219));
    Odrv4 I__11274 (
            .O(N__48219),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ));
    InMux I__11273 (
            .O(N__48216),
            .I(N__48210));
    InMux I__11272 (
            .O(N__48215),
            .I(N__48207));
    CascadeMux I__11271 (
            .O(N__48214),
            .I(N__48204));
    InMux I__11270 (
            .O(N__48213),
            .I(N__48201));
    LocalMux I__11269 (
            .O(N__48210),
            .I(N__48196));
    LocalMux I__11268 (
            .O(N__48207),
            .I(N__48196));
    InMux I__11267 (
            .O(N__48204),
            .I(N__48193));
    LocalMux I__11266 (
            .O(N__48201),
            .I(N__48190));
    Span4Mux_v I__11265 (
            .O(N__48196),
            .I(N__48185));
    LocalMux I__11264 (
            .O(N__48193),
            .I(N__48185));
    Span4Mux_h I__11263 (
            .O(N__48190),
            .I(N__48182));
    Odrv4 I__11262 (
            .O(N__48185),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__11261 (
            .O(N__48182),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__11260 (
            .O(N__48177),
            .I(N__48174));
    LocalMux I__11259 (
            .O(N__48174),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    InMux I__11258 (
            .O(N__48171),
            .I(N__48167));
    InMux I__11257 (
            .O(N__48170),
            .I(N__48164));
    LocalMux I__11256 (
            .O(N__48167),
            .I(N__48159));
    LocalMux I__11255 (
            .O(N__48164),
            .I(N__48156));
    InMux I__11254 (
            .O(N__48163),
            .I(N__48153));
    InMux I__11253 (
            .O(N__48162),
            .I(N__48150));
    Span4Mux_v I__11252 (
            .O(N__48159),
            .I(N__48143));
    Span4Mux_v I__11251 (
            .O(N__48156),
            .I(N__48143));
    LocalMux I__11250 (
            .O(N__48153),
            .I(N__48143));
    LocalMux I__11249 (
            .O(N__48150),
            .I(N__48140));
    Span4Mux_h I__11248 (
            .O(N__48143),
            .I(N__48137));
    Span4Mux_h I__11247 (
            .O(N__48140),
            .I(N__48134));
    Odrv4 I__11246 (
            .O(N__48137),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    Odrv4 I__11245 (
            .O(N__48134),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    CascadeMux I__11244 (
            .O(N__48129),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__11243 (
            .O(N__48126),
            .I(N__48123));
    LocalMux I__11242 (
            .O(N__48123),
            .I(N__48120));
    Odrv12 I__11241 (
            .O(N__48120),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ));
    InMux I__11240 (
            .O(N__48117),
            .I(N__48113));
    CascadeMux I__11239 (
            .O(N__48116),
            .I(N__48110));
    LocalMux I__11238 (
            .O(N__48113),
            .I(N__48106));
    InMux I__11237 (
            .O(N__48110),
            .I(N__48103));
    InMux I__11236 (
            .O(N__48109),
            .I(N__48100));
    Odrv4 I__11235 (
            .O(N__48106),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__11234 (
            .O(N__48103),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    LocalMux I__11233 (
            .O(N__48100),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    CEMux I__11232 (
            .O(N__48093),
            .I(N__48090));
    LocalMux I__11231 (
            .O(N__48090),
            .I(N__48084));
    CEMux I__11230 (
            .O(N__48089),
            .I(N__48081));
    CEMux I__11229 (
            .O(N__48088),
            .I(N__48078));
    CEMux I__11228 (
            .O(N__48087),
            .I(N__48075));
    Span4Mux_h I__11227 (
            .O(N__48084),
            .I(N__48069));
    LocalMux I__11226 (
            .O(N__48081),
            .I(N__48069));
    LocalMux I__11225 (
            .O(N__48078),
            .I(N__48066));
    LocalMux I__11224 (
            .O(N__48075),
            .I(N__48063));
    CEMux I__11223 (
            .O(N__48074),
            .I(N__48060));
    Span4Mux_h I__11222 (
            .O(N__48069),
            .I(N__48057));
    Span4Mux_v I__11221 (
            .O(N__48066),
            .I(N__48054));
    Span4Mux_h I__11220 (
            .O(N__48063),
            .I(N__48051));
    LocalMux I__11219 (
            .O(N__48060),
            .I(N__48048));
    Odrv4 I__11218 (
            .O(N__48057),
            .I(\delay_measurement_inst.delay_hc_timer.N_341_i ));
    Odrv4 I__11217 (
            .O(N__48054),
            .I(\delay_measurement_inst.delay_hc_timer.N_341_i ));
    Odrv4 I__11216 (
            .O(N__48051),
            .I(\delay_measurement_inst.delay_hc_timer.N_341_i ));
    Odrv4 I__11215 (
            .O(N__48048),
            .I(\delay_measurement_inst.delay_hc_timer.N_341_i ));
    InMux I__11214 (
            .O(N__48039),
            .I(N__48033));
    InMux I__11213 (
            .O(N__48038),
            .I(N__48030));
    InMux I__11212 (
            .O(N__48037),
            .I(N__48027));
    InMux I__11211 (
            .O(N__48036),
            .I(N__48024));
    LocalMux I__11210 (
            .O(N__48033),
            .I(N__48019));
    LocalMux I__11209 (
            .O(N__48030),
            .I(N__48019));
    LocalMux I__11208 (
            .O(N__48027),
            .I(N__48016));
    LocalMux I__11207 (
            .O(N__48024),
            .I(N__48013));
    Span4Mux_v I__11206 (
            .O(N__48019),
            .I(N__48010));
    Odrv4 I__11205 (
            .O(N__48016),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv12 I__11204 (
            .O(N__48013),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    Odrv4 I__11203 (
            .O(N__48010),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__11202 (
            .O(N__48003),
            .I(N__48000));
    LocalMux I__11201 (
            .O(N__48000),
            .I(N__47996));
    InMux I__11200 (
            .O(N__47999),
            .I(N__47993));
    Span4Mux_h I__11199 (
            .O(N__47996),
            .I(N__47989));
    LocalMux I__11198 (
            .O(N__47993),
            .I(N__47986));
    InMux I__11197 (
            .O(N__47992),
            .I(N__47983));
    Span4Mux_v I__11196 (
            .O(N__47989),
            .I(N__47978));
    Span4Mux_h I__11195 (
            .O(N__47986),
            .I(N__47978));
    LocalMux I__11194 (
            .O(N__47983),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    Odrv4 I__11193 (
            .O(N__47978),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    CascadeMux I__11192 (
            .O(N__47973),
            .I(N__47970));
    InMux I__11191 (
            .O(N__47970),
            .I(N__47964));
    InMux I__11190 (
            .O(N__47969),
            .I(N__47964));
    LocalMux I__11189 (
            .O(N__47964),
            .I(N__47961));
    Span4Mux_h I__11188 (
            .O(N__47961),
            .I(N__47958));
    Odrv4 I__11187 (
            .O(N__47958),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ));
    CascadeMux I__11186 (
            .O(N__47955),
            .I(N__47951));
    CascadeMux I__11185 (
            .O(N__47954),
            .I(N__47948));
    InMux I__11184 (
            .O(N__47951),
            .I(N__47943));
    InMux I__11183 (
            .O(N__47948),
            .I(N__47943));
    LocalMux I__11182 (
            .O(N__47943),
            .I(N__47940));
    Span4Mux_v I__11181 (
            .O(N__47940),
            .I(N__47937));
    Span4Mux_h I__11180 (
            .O(N__47937),
            .I(N__47934));
    Odrv4 I__11179 (
            .O(N__47934),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ));
    InMux I__11178 (
            .O(N__47931),
            .I(N__47928));
    LocalMux I__11177 (
            .O(N__47928),
            .I(N__47925));
    Odrv12 I__11176 (
            .O(N__47925),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ));
    CascadeMux I__11175 (
            .O(N__47922),
            .I(elapsed_time_ns_1_RNIL73T9_0_9_cascade_));
    CascadeMux I__11174 (
            .O(N__47919),
            .I(N__47916));
    InMux I__11173 (
            .O(N__47916),
            .I(N__47913));
    LocalMux I__11172 (
            .O(N__47913),
            .I(N__47910));
    Odrv12 I__11171 (
            .O(N__47910),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ));
    InMux I__11170 (
            .O(N__47907),
            .I(N__47904));
    LocalMux I__11169 (
            .O(N__47904),
            .I(N__47901));
    Span4Mux_h I__11168 (
            .O(N__47901),
            .I(N__47898));
    Odrv4 I__11167 (
            .O(N__47898),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ));
    InMux I__11166 (
            .O(N__47895),
            .I(N__47889));
    InMux I__11165 (
            .O(N__47894),
            .I(N__47889));
    LocalMux I__11164 (
            .O(N__47889),
            .I(N__47884));
    InMux I__11163 (
            .O(N__47888),
            .I(N__47881));
    InMux I__11162 (
            .O(N__47887),
            .I(N__47878));
    Span4Mux_v I__11161 (
            .O(N__47884),
            .I(N__47875));
    LocalMux I__11160 (
            .O(N__47881),
            .I(N__47872));
    LocalMux I__11159 (
            .O(N__47878),
            .I(N__47869));
    Span4Mux_v I__11158 (
            .O(N__47875),
            .I(N__47866));
    Span4Mux_v I__11157 (
            .O(N__47872),
            .I(N__47861));
    Span4Mux_h I__11156 (
            .O(N__47869),
            .I(N__47861));
    Odrv4 I__11155 (
            .O(N__47866),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    Odrv4 I__11154 (
            .O(N__47861),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__11153 (
            .O(N__47856),
            .I(N__47850));
    InMux I__11152 (
            .O(N__47855),
            .I(N__47847));
    InMux I__11151 (
            .O(N__47854),
            .I(N__47844));
    InMux I__11150 (
            .O(N__47853),
            .I(N__47841));
    LocalMux I__11149 (
            .O(N__47850),
            .I(N__47836));
    LocalMux I__11148 (
            .O(N__47847),
            .I(N__47836));
    LocalMux I__11147 (
            .O(N__47844),
            .I(N__47833));
    LocalMux I__11146 (
            .O(N__47841),
            .I(N__47830));
    Span4Mux_h I__11145 (
            .O(N__47836),
            .I(N__47825));
    Span4Mux_h I__11144 (
            .O(N__47833),
            .I(N__47825));
    Odrv4 I__11143 (
            .O(N__47830),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    Odrv4 I__11142 (
            .O(N__47825),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__11141 (
            .O(N__47820),
            .I(N__47814));
    InMux I__11140 (
            .O(N__47819),
            .I(N__47811));
    InMux I__11139 (
            .O(N__47818),
            .I(N__47808));
    InMux I__11138 (
            .O(N__47817),
            .I(N__47805));
    LocalMux I__11137 (
            .O(N__47814),
            .I(N__47802));
    LocalMux I__11136 (
            .O(N__47811),
            .I(N__47799));
    LocalMux I__11135 (
            .O(N__47808),
            .I(N__47794));
    LocalMux I__11134 (
            .O(N__47805),
            .I(N__47794));
    Span4Mux_h I__11133 (
            .O(N__47802),
            .I(N__47789));
    Span4Mux_h I__11132 (
            .O(N__47799),
            .I(N__47789));
    Odrv4 I__11131 (
            .O(N__47794),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    Odrv4 I__11130 (
            .O(N__47789),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    CascadeMux I__11129 (
            .O(N__47784),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ));
    CascadeMux I__11128 (
            .O(N__47781),
            .I(N__47778));
    InMux I__11127 (
            .O(N__47778),
            .I(N__47775));
    LocalMux I__11126 (
            .O(N__47775),
            .I(N__47772));
    Span4Mux_h I__11125 (
            .O(N__47772),
            .I(N__47769));
    Odrv4 I__11124 (
            .O(N__47769),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    InMux I__11123 (
            .O(N__47766),
            .I(N__47763));
    LocalMux I__11122 (
            .O(N__47763),
            .I(N__47760));
    Sp12to4 I__11121 (
            .O(N__47760),
            .I(N__47757));
    Span12Mux_v I__11120 (
            .O(N__47757),
            .I(N__47754));
    Span12Mux_h I__11119 (
            .O(N__47754),
            .I(N__47751));
    Odrv12 I__11118 (
            .O(N__47751),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    CascadeMux I__11117 (
            .O(N__47748),
            .I(N__47745));
    InMux I__11116 (
            .O(N__47745),
            .I(N__47742));
    LocalMux I__11115 (
            .O(N__47742),
            .I(N__47739));
    Odrv4 I__11114 (
            .O(N__47739),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__11113 (
            .O(N__47736),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    CascadeMux I__11112 (
            .O(N__47733),
            .I(N__47730));
    InMux I__11111 (
            .O(N__47730),
            .I(N__47727));
    LocalMux I__11110 (
            .O(N__47727),
            .I(N__47724));
    Span12Mux_s7_h I__11109 (
            .O(N__47724),
            .I(N__47721));
    Span12Mux_v I__11108 (
            .O(N__47721),
            .I(N__47718));
    Span12Mux_h I__11107 (
            .O(N__47718),
            .I(N__47715));
    Odrv12 I__11106 (
            .O(N__47715),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    CascadeMux I__11105 (
            .O(N__47712),
            .I(N__47709));
    InMux I__11104 (
            .O(N__47709),
            .I(N__47706));
    LocalMux I__11103 (
            .O(N__47706),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__11102 (
            .O(N__47703),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__11101 (
            .O(N__47700),
            .I(N__47697));
    LocalMux I__11100 (
            .O(N__47697),
            .I(N__47694));
    Sp12to4 I__11099 (
            .O(N__47694),
            .I(N__47691));
    Span12Mux_h I__11098 (
            .O(N__47691),
            .I(N__47688));
    Span12Mux_v I__11097 (
            .O(N__47688),
            .I(N__47685));
    Odrv12 I__11096 (
            .O(N__47685),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__11095 (
            .O(N__47682),
            .I(N__47679));
    LocalMux I__11094 (
            .O(N__47679),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__11093 (
            .O(N__47676),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    CascadeMux I__11092 (
            .O(N__47673),
            .I(N__47670));
    InMux I__11091 (
            .O(N__47670),
            .I(N__47667));
    LocalMux I__11090 (
            .O(N__47667),
            .I(N__47664));
    Sp12to4 I__11089 (
            .O(N__47664),
            .I(N__47661));
    Span12Mux_h I__11088 (
            .O(N__47661),
            .I(N__47658));
    Span12Mux_v I__11087 (
            .O(N__47658),
            .I(N__47655));
    Odrv12 I__11086 (
            .O(N__47655),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    CascadeMux I__11085 (
            .O(N__47652),
            .I(N__47649));
    InMux I__11084 (
            .O(N__47649),
            .I(N__47646));
    LocalMux I__11083 (
            .O(N__47646),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__11082 (
            .O(N__47643),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__11081 (
            .O(N__47640),
            .I(N__47637));
    LocalMux I__11080 (
            .O(N__47637),
            .I(N__47634));
    Span12Mux_h I__11079 (
            .O(N__47634),
            .I(N__47631));
    Span12Mux_v I__11078 (
            .O(N__47631),
            .I(N__47628));
    Odrv12 I__11077 (
            .O(N__47628),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    CascadeMux I__11076 (
            .O(N__47625),
            .I(N__47622));
    InMux I__11075 (
            .O(N__47622),
            .I(N__47619));
    LocalMux I__11074 (
            .O(N__47619),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__11073 (
            .O(N__47616),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    CascadeMux I__11072 (
            .O(N__47613),
            .I(N__47603));
    CascadeMux I__11071 (
            .O(N__47612),
            .I(N__47599));
    CascadeMux I__11070 (
            .O(N__47611),
            .I(N__47595));
    CascadeMux I__11069 (
            .O(N__47610),
            .I(N__47591));
    CascadeMux I__11068 (
            .O(N__47609),
            .I(N__47587));
    CascadeMux I__11067 (
            .O(N__47608),
            .I(N__47584));
    InMux I__11066 (
            .O(N__47607),
            .I(N__47581));
    InMux I__11065 (
            .O(N__47606),
            .I(N__47566));
    InMux I__11064 (
            .O(N__47603),
            .I(N__47566));
    InMux I__11063 (
            .O(N__47602),
            .I(N__47566));
    InMux I__11062 (
            .O(N__47599),
            .I(N__47566));
    InMux I__11061 (
            .O(N__47598),
            .I(N__47566));
    InMux I__11060 (
            .O(N__47595),
            .I(N__47566));
    InMux I__11059 (
            .O(N__47594),
            .I(N__47566));
    InMux I__11058 (
            .O(N__47591),
            .I(N__47563));
    InMux I__11057 (
            .O(N__47590),
            .I(N__47556));
    InMux I__11056 (
            .O(N__47587),
            .I(N__47556));
    InMux I__11055 (
            .O(N__47584),
            .I(N__47556));
    LocalMux I__11054 (
            .O(N__47581),
            .I(N__47553));
    LocalMux I__11053 (
            .O(N__47566),
            .I(N__47546));
    LocalMux I__11052 (
            .O(N__47563),
            .I(N__47546));
    LocalMux I__11051 (
            .O(N__47556),
            .I(N__47546));
    Span12Mux_h I__11050 (
            .O(N__47553),
            .I(N__47543));
    Span12Mux_v I__11049 (
            .O(N__47546),
            .I(N__47540));
    Odrv12 I__11048 (
            .O(N__47543),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    Odrv12 I__11047 (
            .O(N__47540),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    CascadeMux I__11046 (
            .O(N__47535),
            .I(N__47532));
    InMux I__11045 (
            .O(N__47532),
            .I(N__47529));
    LocalMux I__11044 (
            .O(N__47529),
            .I(N__47526));
    Sp12to4 I__11043 (
            .O(N__47526),
            .I(N__47523));
    Span12Mux_h I__11042 (
            .O(N__47523),
            .I(N__47520));
    Span12Mux_v I__11041 (
            .O(N__47520),
            .I(N__47517));
    Odrv12 I__11040 (
            .O(N__47517),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    CascadeMux I__11039 (
            .O(N__47514),
            .I(N__47511));
    InMux I__11038 (
            .O(N__47511),
            .I(N__47508));
    LocalMux I__11037 (
            .O(N__47508),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__11036 (
            .O(N__47505),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__11035 (
            .O(N__47502),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__11034 (
            .O(N__47499),
            .I(N__47496));
    LocalMux I__11033 (
            .O(N__47496),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    IoInMux I__11032 (
            .O(N__47493),
            .I(N__47490));
    LocalMux I__11031 (
            .O(N__47490),
            .I(GB_BUFFER_clock_output_0_THRU_CO));
    InMux I__11030 (
            .O(N__47487),
            .I(N__47484));
    LocalMux I__11029 (
            .O(N__47484),
            .I(N__47481));
    Sp12to4 I__11028 (
            .O(N__47481),
            .I(N__47478));
    Span12Mux_v I__11027 (
            .O(N__47478),
            .I(N__47475));
    Span12Mux_h I__11026 (
            .O(N__47475),
            .I(N__47472));
    Odrv12 I__11025 (
            .O(N__47472),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__11024 (
            .O(N__47469),
            .I(N__47466));
    InMux I__11023 (
            .O(N__47466),
            .I(N__47463));
    LocalMux I__11022 (
            .O(N__47463),
            .I(N__47460));
    Span4Mux_h I__11021 (
            .O(N__47460),
            .I(N__47457));
    Span4Mux_h I__11020 (
            .O(N__47457),
            .I(N__47454));
    Odrv4 I__11019 (
            .O(N__47454),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    CascadeMux I__11018 (
            .O(N__47451),
            .I(N__47448));
    InMux I__11017 (
            .O(N__47448),
            .I(N__47445));
    LocalMux I__11016 (
            .O(N__47445),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__11015 (
            .O(N__47442),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__11014 (
            .O(N__47439),
            .I(N__47436));
    LocalMux I__11013 (
            .O(N__47436),
            .I(N__47433));
    Span12Mux_v I__11012 (
            .O(N__47433),
            .I(N__47430));
    Span12Mux_h I__11011 (
            .O(N__47430),
            .I(N__47427));
    Odrv12 I__11010 (
            .O(N__47427),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__11009 (
            .O(N__47424),
            .I(N__47421));
    InMux I__11008 (
            .O(N__47421),
            .I(N__47418));
    LocalMux I__11007 (
            .O(N__47418),
            .I(N__47415));
    Span4Mux_h I__11006 (
            .O(N__47415),
            .I(N__47412));
    Span4Mux_h I__11005 (
            .O(N__47412),
            .I(N__47409));
    Odrv4 I__11004 (
            .O(N__47409),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    CascadeMux I__11003 (
            .O(N__47406),
            .I(N__47403));
    InMux I__11002 (
            .O(N__47403),
            .I(N__47400));
    LocalMux I__11001 (
            .O(N__47400),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__11000 (
            .O(N__47397),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__10999 (
            .O(N__47394),
            .I(N__47391));
    LocalMux I__10998 (
            .O(N__47391),
            .I(N__47388));
    Span12Mux_s8_h I__10997 (
            .O(N__47388),
            .I(N__47385));
    Span12Mux_h I__10996 (
            .O(N__47385),
            .I(N__47382));
    Span12Mux_v I__10995 (
            .O(N__47382),
            .I(N__47379));
    Odrv12 I__10994 (
            .O(N__47379),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__10993 (
            .O(N__47376),
            .I(N__47373));
    InMux I__10992 (
            .O(N__47373),
            .I(N__47370));
    LocalMux I__10991 (
            .O(N__47370),
            .I(N__47367));
    Span4Mux_h I__10990 (
            .O(N__47367),
            .I(N__47364));
    Span4Mux_h I__10989 (
            .O(N__47364),
            .I(N__47361));
    Odrv4 I__10988 (
            .O(N__47361),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    CascadeMux I__10987 (
            .O(N__47358),
            .I(N__47355));
    InMux I__10986 (
            .O(N__47355),
            .I(N__47352));
    LocalMux I__10985 (
            .O(N__47352),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__10984 (
            .O(N__47349),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__10983 (
            .O(N__47346),
            .I(N__47343));
    LocalMux I__10982 (
            .O(N__47343),
            .I(N__47340));
    Span12Mux_s9_h I__10981 (
            .O(N__47340),
            .I(N__47337));
    Span12Mux_v I__10980 (
            .O(N__47337),
            .I(N__47334));
    Span12Mux_h I__10979 (
            .O(N__47334),
            .I(N__47331));
    Odrv12 I__10978 (
            .O(N__47331),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    CascadeMux I__10977 (
            .O(N__47328),
            .I(N__47325));
    InMux I__10976 (
            .O(N__47325),
            .I(N__47322));
    LocalMux I__10975 (
            .O(N__47322),
            .I(N__47319));
    Odrv4 I__10974 (
            .O(N__47319),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__10973 (
            .O(N__47316),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__10972 (
            .O(N__47313),
            .I(N__47310));
    LocalMux I__10971 (
            .O(N__47310),
            .I(N__47307));
    Span12Mux_h I__10970 (
            .O(N__47307),
            .I(N__47304));
    Span12Mux_v I__10969 (
            .O(N__47304),
            .I(N__47301));
    Odrv12 I__10968 (
            .O(N__47301),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    CascadeMux I__10967 (
            .O(N__47298),
            .I(N__47295));
    InMux I__10966 (
            .O(N__47295),
            .I(N__47292));
    LocalMux I__10965 (
            .O(N__47292),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__10964 (
            .O(N__47289),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__10963 (
            .O(N__47286),
            .I(N__47283));
    LocalMux I__10962 (
            .O(N__47283),
            .I(N__47280));
    Span12Mux_h I__10961 (
            .O(N__47280),
            .I(N__47277));
    Span12Mux_v I__10960 (
            .O(N__47277),
            .I(N__47274));
    Odrv12 I__10959 (
            .O(N__47274),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    CascadeMux I__10958 (
            .O(N__47271),
            .I(N__47268));
    InMux I__10957 (
            .O(N__47268),
            .I(N__47265));
    LocalMux I__10956 (
            .O(N__47265),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__10955 (
            .O(N__47262),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    CascadeMux I__10954 (
            .O(N__47259),
            .I(N__47256));
    InMux I__10953 (
            .O(N__47256),
            .I(N__47253));
    LocalMux I__10952 (
            .O(N__47253),
            .I(N__47250));
    Span12Mux_h I__10951 (
            .O(N__47250),
            .I(N__47247));
    Span12Mux_v I__10950 (
            .O(N__47247),
            .I(N__47244));
    Odrv12 I__10949 (
            .O(N__47244),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    CascadeMux I__10948 (
            .O(N__47241),
            .I(N__47238));
    InMux I__10947 (
            .O(N__47238),
            .I(N__47235));
    LocalMux I__10946 (
            .O(N__47235),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__10945 (
            .O(N__47232),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    CascadeMux I__10944 (
            .O(N__47229),
            .I(N__47226));
    InMux I__10943 (
            .O(N__47226),
            .I(N__47223));
    LocalMux I__10942 (
            .O(N__47223),
            .I(N__47220));
    Span12Mux_h I__10941 (
            .O(N__47220),
            .I(N__47217));
    Span12Mux_v I__10940 (
            .O(N__47217),
            .I(N__47214));
    Odrv12 I__10939 (
            .O(N__47214),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    CascadeMux I__10938 (
            .O(N__47211),
            .I(N__47208));
    InMux I__10937 (
            .O(N__47208),
            .I(N__47205));
    LocalMux I__10936 (
            .O(N__47205),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__10935 (
            .O(N__47202),
            .I(bfn_18_23_0_));
    InMux I__10934 (
            .O(N__47199),
            .I(N__47196));
    LocalMux I__10933 (
            .O(N__47196),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt30 ));
    CascadeMux I__10932 (
            .O(N__47193),
            .I(N__47190));
    InMux I__10931 (
            .O(N__47190),
            .I(N__47187));
    LocalMux I__10930 (
            .O(N__47187),
            .I(N__47184));
    Odrv4 I__10929 (
            .O(N__47184),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ));
    InMux I__10928 (
            .O(N__47181),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_0_30 ));
    CascadeMux I__10927 (
            .O(N__47178),
            .I(N__47175));
    InMux I__10926 (
            .O(N__47175),
            .I(N__47169));
    InMux I__10925 (
            .O(N__47174),
            .I(N__47169));
    LocalMux I__10924 (
            .O(N__47169),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_CO ));
    IoInMux I__10923 (
            .O(N__47166),
            .I(N__47137));
    InMux I__10922 (
            .O(N__47165),
            .I(N__47124));
    InMux I__10921 (
            .O(N__47164),
            .I(N__47124));
    InMux I__10920 (
            .O(N__47163),
            .I(N__47124));
    InMux I__10919 (
            .O(N__47162),
            .I(N__47124));
    InMux I__10918 (
            .O(N__47161),
            .I(N__47117));
    InMux I__10917 (
            .O(N__47160),
            .I(N__47117));
    InMux I__10916 (
            .O(N__47159),
            .I(N__47117));
    InMux I__10915 (
            .O(N__47158),
            .I(N__47108));
    InMux I__10914 (
            .O(N__47157),
            .I(N__47108));
    InMux I__10913 (
            .O(N__47156),
            .I(N__47108));
    InMux I__10912 (
            .O(N__47155),
            .I(N__47108));
    InMux I__10911 (
            .O(N__47154),
            .I(N__47098));
    InMux I__10910 (
            .O(N__47153),
            .I(N__47098));
    InMux I__10909 (
            .O(N__47152),
            .I(N__47098));
    InMux I__10908 (
            .O(N__47151),
            .I(N__47098));
    InMux I__10907 (
            .O(N__47150),
            .I(N__47089));
    InMux I__10906 (
            .O(N__47149),
            .I(N__47089));
    InMux I__10905 (
            .O(N__47148),
            .I(N__47089));
    InMux I__10904 (
            .O(N__47147),
            .I(N__47089));
    InMux I__10903 (
            .O(N__47146),
            .I(N__47082));
    InMux I__10902 (
            .O(N__47145),
            .I(N__47082));
    InMux I__10901 (
            .O(N__47144),
            .I(N__47082));
    InMux I__10900 (
            .O(N__47143),
            .I(N__47073));
    InMux I__10899 (
            .O(N__47142),
            .I(N__47073));
    InMux I__10898 (
            .O(N__47141),
            .I(N__47073));
    InMux I__10897 (
            .O(N__47140),
            .I(N__47073));
    LocalMux I__10896 (
            .O(N__47137),
            .I(N__47070));
    InMux I__10895 (
            .O(N__47136),
            .I(N__47061));
    InMux I__10894 (
            .O(N__47135),
            .I(N__47061));
    InMux I__10893 (
            .O(N__47134),
            .I(N__47061));
    InMux I__10892 (
            .O(N__47133),
            .I(N__47061));
    LocalMux I__10891 (
            .O(N__47124),
            .I(N__47056));
    LocalMux I__10890 (
            .O(N__47117),
            .I(N__47056));
    LocalMux I__10889 (
            .O(N__47108),
            .I(N__47053));
    InMux I__10888 (
            .O(N__47107),
            .I(N__47050));
    LocalMux I__10887 (
            .O(N__47098),
            .I(N__47047));
    LocalMux I__10886 (
            .O(N__47089),
            .I(N__47040));
    LocalMux I__10885 (
            .O(N__47082),
            .I(N__47040));
    LocalMux I__10884 (
            .O(N__47073),
            .I(N__47040));
    Span4Mux_s1_v I__10883 (
            .O(N__47070),
            .I(N__47037));
    LocalMux I__10882 (
            .O(N__47061),
            .I(N__47034));
    Span4Mux_v I__10881 (
            .O(N__47056),
            .I(N__47029));
    Span4Mux_v I__10880 (
            .O(N__47053),
            .I(N__47029));
    LocalMux I__10879 (
            .O(N__47050),
            .I(N__47022));
    Span4Mux_h I__10878 (
            .O(N__47047),
            .I(N__47022));
    Span4Mux_v I__10877 (
            .O(N__47040),
            .I(N__47022));
    Span4Mux_h I__10876 (
            .O(N__47037),
            .I(N__47019));
    Span4Mux_h I__10875 (
            .O(N__47034),
            .I(N__47016));
    Span4Mux_v I__10874 (
            .O(N__47029),
            .I(N__47011));
    Span4Mux_v I__10873 (
            .O(N__47022),
            .I(N__47011));
    Span4Mux_h I__10872 (
            .O(N__47019),
            .I(N__47008));
    Span4Mux_v I__10871 (
            .O(N__47016),
            .I(N__47005));
    Span4Mux_h I__10870 (
            .O(N__47011),
            .I(N__47000));
    Span4Mux_v I__10869 (
            .O(N__47008),
            .I(N__47000));
    Odrv4 I__10868 (
            .O(N__47005),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    Odrv4 I__10867 (
            .O(N__47000),
            .I(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ));
    InMux I__10866 (
            .O(N__46995),
            .I(N__46991));
    InMux I__10865 (
            .O(N__46994),
            .I(N__46988));
    LocalMux I__10864 (
            .O(N__46991),
            .I(N__46985));
    LocalMux I__10863 (
            .O(N__46988),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30 ));
    Odrv12 I__10862 (
            .O(N__46985),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30 ));
    InMux I__10861 (
            .O(N__46980),
            .I(N__46977));
    LocalMux I__10860 (
            .O(N__46977),
            .I(N__46972));
    InMux I__10859 (
            .O(N__46976),
            .I(N__46969));
    InMux I__10858 (
            .O(N__46975),
            .I(N__46966));
    Span4Mux_v I__10857 (
            .O(N__46972),
            .I(N__46961));
    LocalMux I__10856 (
            .O(N__46969),
            .I(N__46961));
    LocalMux I__10855 (
            .O(N__46966),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__10854 (
            .O(N__46961),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ));
    InMux I__10853 (
            .O(N__46956),
            .I(N__46953));
    LocalMux I__10852 (
            .O(N__46953),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__10851 (
            .O(N__46950),
            .I(N__46947));
    LocalMux I__10850 (
            .O(N__46947),
            .I(N__46944));
    Span4Mux_v I__10849 (
            .O(N__46944),
            .I(N__46940));
    InMux I__10848 (
            .O(N__46943),
            .I(N__46937));
    Sp12to4 I__10847 (
            .O(N__46940),
            .I(N__46933));
    LocalMux I__10846 (
            .O(N__46937),
            .I(N__46929));
    InMux I__10845 (
            .O(N__46936),
            .I(N__46926));
    Span12Mux_h I__10844 (
            .O(N__46933),
            .I(N__46923));
    InMux I__10843 (
            .O(N__46932),
            .I(N__46920));
    Span4Mux_v I__10842 (
            .O(N__46929),
            .I(N__46915));
    LocalMux I__10841 (
            .O(N__46926),
            .I(N__46915));
    Odrv12 I__10840 (
            .O(N__46923),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__10839 (
            .O(N__46920),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__10838 (
            .O(N__46915),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    CascadeMux I__10837 (
            .O(N__46908),
            .I(N__46905));
    InMux I__10836 (
            .O(N__46905),
            .I(N__46902));
    LocalMux I__10835 (
            .O(N__46902),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    CascadeMux I__10834 (
            .O(N__46899),
            .I(N__46896));
    InMux I__10833 (
            .O(N__46896),
            .I(N__46893));
    LocalMux I__10832 (
            .O(N__46893),
            .I(N__46888));
    CascadeMux I__10831 (
            .O(N__46892),
            .I(N__46885));
    InMux I__10830 (
            .O(N__46891),
            .I(N__46882));
    Span4Mux_v I__10829 (
            .O(N__46888),
            .I(N__46879));
    InMux I__10828 (
            .O(N__46885),
            .I(N__46876));
    LocalMux I__10827 (
            .O(N__46882),
            .I(N__46873));
    Sp12to4 I__10826 (
            .O(N__46879),
            .I(N__46869));
    LocalMux I__10825 (
            .O(N__46876),
            .I(N__46866));
    Span4Mux_h I__10824 (
            .O(N__46873),
            .I(N__46863));
    InMux I__10823 (
            .O(N__46872),
            .I(N__46860));
    Span12Mux_h I__10822 (
            .O(N__46869),
            .I(N__46857));
    Odrv4 I__10821 (
            .O(N__46866),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__10820 (
            .O(N__46863),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    LocalMux I__10819 (
            .O(N__46860),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv12 I__10818 (
            .O(N__46857),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    CascadeMux I__10817 (
            .O(N__46848),
            .I(N__46845));
    InMux I__10816 (
            .O(N__46845),
            .I(N__46842));
    LocalMux I__10815 (
            .O(N__46842),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    CascadeMux I__10814 (
            .O(N__46839),
            .I(N__46835));
    CascadeMux I__10813 (
            .O(N__46838),
            .I(N__46832));
    InMux I__10812 (
            .O(N__46835),
            .I(N__46829));
    InMux I__10811 (
            .O(N__46832),
            .I(N__46826));
    LocalMux I__10810 (
            .O(N__46829),
            .I(N__46822));
    LocalMux I__10809 (
            .O(N__46826),
            .I(N__46819));
    InMux I__10808 (
            .O(N__46825),
            .I(N__46816));
    Span4Mux_v I__10807 (
            .O(N__46822),
            .I(N__46813));
    Span4Mux_v I__10806 (
            .O(N__46819),
            .I(N__46810));
    LocalMux I__10805 (
            .O(N__46816),
            .I(N__46807));
    Sp12to4 I__10804 (
            .O(N__46813),
            .I(N__46801));
    Sp12to4 I__10803 (
            .O(N__46810),
            .I(N__46801));
    Span4Mux_v I__10802 (
            .O(N__46807),
            .I(N__46798));
    InMux I__10801 (
            .O(N__46806),
            .I(N__46795));
    Span12Mux_h I__10800 (
            .O(N__46801),
            .I(N__46792));
    Odrv4 I__10799 (
            .O(N__46798),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    LocalMux I__10798 (
            .O(N__46795),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv12 I__10797 (
            .O(N__46792),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    CascadeMux I__10796 (
            .O(N__46785),
            .I(N__46771));
    CascadeMux I__10795 (
            .O(N__46784),
            .I(N__46758));
    CascadeMux I__10794 (
            .O(N__46783),
            .I(N__46755));
    CascadeMux I__10793 (
            .O(N__46782),
            .I(N__46752));
    CascadeMux I__10792 (
            .O(N__46781),
            .I(N__46745));
    InMux I__10791 (
            .O(N__46780),
            .I(N__46742));
    InMux I__10790 (
            .O(N__46779),
            .I(N__46729));
    InMux I__10789 (
            .O(N__46778),
            .I(N__46729));
    InMux I__10788 (
            .O(N__46777),
            .I(N__46729));
    InMux I__10787 (
            .O(N__46776),
            .I(N__46729));
    InMux I__10786 (
            .O(N__46775),
            .I(N__46729));
    InMux I__10785 (
            .O(N__46774),
            .I(N__46729));
    InMux I__10784 (
            .O(N__46771),
            .I(N__46726));
    InMux I__10783 (
            .O(N__46770),
            .I(N__46721));
    InMux I__10782 (
            .O(N__46769),
            .I(N__46721));
    InMux I__10781 (
            .O(N__46768),
            .I(N__46714));
    InMux I__10780 (
            .O(N__46767),
            .I(N__46714));
    CascadeMux I__10779 (
            .O(N__46766),
            .I(N__46708));
    CascadeMux I__10778 (
            .O(N__46765),
            .I(N__46705));
    CascadeMux I__10777 (
            .O(N__46764),
            .I(N__46702));
    InMux I__10776 (
            .O(N__46763),
            .I(N__46689));
    InMux I__10775 (
            .O(N__46762),
            .I(N__46689));
    InMux I__10774 (
            .O(N__46761),
            .I(N__46689));
    InMux I__10773 (
            .O(N__46758),
            .I(N__46689));
    InMux I__10772 (
            .O(N__46755),
            .I(N__46689));
    InMux I__10771 (
            .O(N__46752),
            .I(N__46689));
    InMux I__10770 (
            .O(N__46751),
            .I(N__46686));
    InMux I__10769 (
            .O(N__46750),
            .I(N__46683));
    InMux I__10768 (
            .O(N__46749),
            .I(N__46676));
    InMux I__10767 (
            .O(N__46748),
            .I(N__46676));
    InMux I__10766 (
            .O(N__46745),
            .I(N__46676));
    LocalMux I__10765 (
            .O(N__46742),
            .I(N__46673));
    LocalMux I__10764 (
            .O(N__46729),
            .I(N__46668));
    LocalMux I__10763 (
            .O(N__46726),
            .I(N__46668));
    LocalMux I__10762 (
            .O(N__46721),
            .I(N__46665));
    InMux I__10761 (
            .O(N__46720),
            .I(N__46660));
    InMux I__10760 (
            .O(N__46719),
            .I(N__46660));
    LocalMux I__10759 (
            .O(N__46714),
            .I(N__46657));
    InMux I__10758 (
            .O(N__46713),
            .I(N__46644));
    InMux I__10757 (
            .O(N__46712),
            .I(N__46644));
    InMux I__10756 (
            .O(N__46711),
            .I(N__46644));
    InMux I__10755 (
            .O(N__46708),
            .I(N__46644));
    InMux I__10754 (
            .O(N__46705),
            .I(N__46644));
    InMux I__10753 (
            .O(N__46702),
            .I(N__46644));
    LocalMux I__10752 (
            .O(N__46689),
            .I(N__46641));
    LocalMux I__10751 (
            .O(N__46686),
            .I(N__46634));
    LocalMux I__10750 (
            .O(N__46683),
            .I(N__46634));
    LocalMux I__10749 (
            .O(N__46676),
            .I(N__46634));
    Span4Mux_v I__10748 (
            .O(N__46673),
            .I(N__46629));
    Span4Mux_v I__10747 (
            .O(N__46668),
            .I(N__46629));
    Span12Mux_h I__10746 (
            .O(N__46665),
            .I(N__46624));
    LocalMux I__10745 (
            .O(N__46660),
            .I(N__46624));
    Span4Mux_h I__10744 (
            .O(N__46657),
            .I(N__46621));
    LocalMux I__10743 (
            .O(N__46644),
            .I(\current_shift_inst.PI_CTRL.N_289 ));
    Odrv4 I__10742 (
            .O(N__46641),
            .I(\current_shift_inst.PI_CTRL.N_289 ));
    Odrv4 I__10741 (
            .O(N__46634),
            .I(\current_shift_inst.PI_CTRL.N_289 ));
    Odrv4 I__10740 (
            .O(N__46629),
            .I(\current_shift_inst.PI_CTRL.N_289 ));
    Odrv12 I__10739 (
            .O(N__46624),
            .I(\current_shift_inst.PI_CTRL.N_289 ));
    Odrv4 I__10738 (
            .O(N__46621),
            .I(\current_shift_inst.PI_CTRL.N_289 ));
    InMux I__10737 (
            .O(N__46608),
            .I(N__46604));
    InMux I__10736 (
            .O(N__46607),
            .I(N__46601));
    LocalMux I__10735 (
            .O(N__46604),
            .I(N__46598));
    LocalMux I__10734 (
            .O(N__46601),
            .I(N__46590));
    Span4Mux_v I__10733 (
            .O(N__46598),
            .I(N__46586));
    InMux I__10732 (
            .O(N__46597),
            .I(N__46576));
    InMux I__10731 (
            .O(N__46596),
            .I(N__46571));
    InMux I__10730 (
            .O(N__46595),
            .I(N__46571));
    InMux I__10729 (
            .O(N__46594),
            .I(N__46566));
    InMux I__10728 (
            .O(N__46593),
            .I(N__46566));
    Span4Mux_v I__10727 (
            .O(N__46590),
            .I(N__46557));
    InMux I__10726 (
            .O(N__46589),
            .I(N__46553));
    Span4Mux_h I__10725 (
            .O(N__46586),
            .I(N__46550));
    InMux I__10724 (
            .O(N__46585),
            .I(N__46547));
    InMux I__10723 (
            .O(N__46584),
            .I(N__46525));
    InMux I__10722 (
            .O(N__46583),
            .I(N__46525));
    InMux I__10721 (
            .O(N__46582),
            .I(N__46525));
    InMux I__10720 (
            .O(N__46581),
            .I(N__46525));
    InMux I__10719 (
            .O(N__46580),
            .I(N__46525));
    InMux I__10718 (
            .O(N__46579),
            .I(N__46525));
    LocalMux I__10717 (
            .O(N__46576),
            .I(N__46522));
    LocalMux I__10716 (
            .O(N__46571),
            .I(N__46517));
    LocalMux I__10715 (
            .O(N__46566),
            .I(N__46517));
    InMux I__10714 (
            .O(N__46565),
            .I(N__46503));
    InMux I__10713 (
            .O(N__46564),
            .I(N__46503));
    InMux I__10712 (
            .O(N__46563),
            .I(N__46503));
    InMux I__10711 (
            .O(N__46562),
            .I(N__46503));
    InMux I__10710 (
            .O(N__46561),
            .I(N__46503));
    InMux I__10709 (
            .O(N__46560),
            .I(N__46503));
    Span4Mux_h I__10708 (
            .O(N__46557),
            .I(N__46500));
    InMux I__10707 (
            .O(N__46556),
            .I(N__46497));
    LocalMux I__10706 (
            .O(N__46553),
            .I(N__46490));
    Span4Mux_h I__10705 (
            .O(N__46550),
            .I(N__46490));
    LocalMux I__10704 (
            .O(N__46547),
            .I(N__46490));
    InMux I__10703 (
            .O(N__46546),
            .I(N__46487));
    InMux I__10702 (
            .O(N__46545),
            .I(N__46482));
    InMux I__10701 (
            .O(N__46544),
            .I(N__46482));
    InMux I__10700 (
            .O(N__46543),
            .I(N__46469));
    InMux I__10699 (
            .O(N__46542),
            .I(N__46469));
    InMux I__10698 (
            .O(N__46541),
            .I(N__46469));
    InMux I__10697 (
            .O(N__46540),
            .I(N__46469));
    InMux I__10696 (
            .O(N__46539),
            .I(N__46469));
    InMux I__10695 (
            .O(N__46538),
            .I(N__46469));
    LocalMux I__10694 (
            .O(N__46525),
            .I(N__46462));
    Span4Mux_v I__10693 (
            .O(N__46522),
            .I(N__46462));
    Span4Mux_v I__10692 (
            .O(N__46517),
            .I(N__46462));
    InMux I__10691 (
            .O(N__46516),
            .I(N__46459));
    LocalMux I__10690 (
            .O(N__46503),
            .I(N__46452));
    Span4Mux_h I__10689 (
            .O(N__46500),
            .I(N__46452));
    LocalMux I__10688 (
            .O(N__46497),
            .I(N__46452));
    Span4Mux_v I__10687 (
            .O(N__46490),
            .I(N__46449));
    LocalMux I__10686 (
            .O(N__46487),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__10685 (
            .O(N__46482),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__10684 (
            .O(N__46469),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__10683 (
            .O(N__46462),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__10682 (
            .O(N__46459),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__10681 (
            .O(N__46452),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__10680 (
            .O(N__46449),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    CascadeMux I__10679 (
            .O(N__46434),
            .I(N__46431));
    InMux I__10678 (
            .O(N__46431),
            .I(N__46428));
    LocalMux I__10677 (
            .O(N__46428),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    CascadeMux I__10676 (
            .O(N__46425),
            .I(N__46413));
    CascadeMux I__10675 (
            .O(N__46424),
            .I(N__46410));
    CascadeMux I__10674 (
            .O(N__46423),
            .I(N__46407));
    CascadeMux I__10673 (
            .O(N__46422),
            .I(N__46404));
    CascadeMux I__10672 (
            .O(N__46421),
            .I(N__46398));
    CascadeMux I__10671 (
            .O(N__46420),
            .I(N__46395));
    CascadeMux I__10670 (
            .O(N__46419),
            .I(N__46380));
    InMux I__10669 (
            .O(N__46418),
            .I(N__46375));
    InMux I__10668 (
            .O(N__46417),
            .I(N__46359));
    InMux I__10667 (
            .O(N__46416),
            .I(N__46359));
    InMux I__10666 (
            .O(N__46413),
            .I(N__46359));
    InMux I__10665 (
            .O(N__46410),
            .I(N__46359));
    InMux I__10664 (
            .O(N__46407),
            .I(N__46359));
    InMux I__10663 (
            .O(N__46404),
            .I(N__46359));
    InMux I__10662 (
            .O(N__46403),
            .I(N__46346));
    InMux I__10661 (
            .O(N__46402),
            .I(N__46346));
    InMux I__10660 (
            .O(N__46401),
            .I(N__46346));
    InMux I__10659 (
            .O(N__46398),
            .I(N__46346));
    InMux I__10658 (
            .O(N__46395),
            .I(N__46346));
    InMux I__10657 (
            .O(N__46394),
            .I(N__46346));
    InMux I__10656 (
            .O(N__46393),
            .I(N__46343));
    InMux I__10655 (
            .O(N__46392),
            .I(N__46330));
    InMux I__10654 (
            .O(N__46391),
            .I(N__46330));
    InMux I__10653 (
            .O(N__46390),
            .I(N__46330));
    InMux I__10652 (
            .O(N__46389),
            .I(N__46330));
    InMux I__10651 (
            .O(N__46388),
            .I(N__46330));
    InMux I__10650 (
            .O(N__46387),
            .I(N__46330));
    CascadeMux I__10649 (
            .O(N__46386),
            .I(N__46326));
    InMux I__10648 (
            .O(N__46385),
            .I(N__46323));
    InMux I__10647 (
            .O(N__46384),
            .I(N__46320));
    InMux I__10646 (
            .O(N__46383),
            .I(N__46315));
    InMux I__10645 (
            .O(N__46380),
            .I(N__46315));
    InMux I__10644 (
            .O(N__46379),
            .I(N__46312));
    InMux I__10643 (
            .O(N__46378),
            .I(N__46309));
    LocalMux I__10642 (
            .O(N__46375),
            .I(N__46306));
    InMux I__10641 (
            .O(N__46374),
            .I(N__46299));
    InMux I__10640 (
            .O(N__46373),
            .I(N__46299));
    InMux I__10639 (
            .O(N__46372),
            .I(N__46299));
    LocalMux I__10638 (
            .O(N__46359),
            .I(N__46294));
    LocalMux I__10637 (
            .O(N__46346),
            .I(N__46294));
    LocalMux I__10636 (
            .O(N__46343),
            .I(N__46289));
    LocalMux I__10635 (
            .O(N__46330),
            .I(N__46289));
    InMux I__10634 (
            .O(N__46329),
            .I(N__46284));
    InMux I__10633 (
            .O(N__46326),
            .I(N__46284));
    LocalMux I__10632 (
            .O(N__46323),
            .I(N__46279));
    LocalMux I__10631 (
            .O(N__46320),
            .I(N__46279));
    LocalMux I__10630 (
            .O(N__46315),
            .I(N__46276));
    LocalMux I__10629 (
            .O(N__46312),
            .I(N__46263));
    LocalMux I__10628 (
            .O(N__46309),
            .I(N__46263));
    Span4Mux_v I__10627 (
            .O(N__46306),
            .I(N__46263));
    LocalMux I__10626 (
            .O(N__46299),
            .I(N__46263));
    Span4Mux_v I__10625 (
            .O(N__46294),
            .I(N__46263));
    Span4Mux_v I__10624 (
            .O(N__46289),
            .I(N__46263));
    LocalMux I__10623 (
            .O(N__46284),
            .I(N__46256));
    Span12Mux_s10_v I__10622 (
            .O(N__46279),
            .I(N__46256));
    Span12Mux_s7_h I__10621 (
            .O(N__46276),
            .I(N__46256));
    Span4Mux_h I__10620 (
            .O(N__46263),
            .I(N__46253));
    Odrv12 I__10619 (
            .O(N__46256),
            .I(\current_shift_inst.PI_CTRL.N_290 ));
    Odrv4 I__10618 (
            .O(N__46253),
            .I(\current_shift_inst.PI_CTRL.N_290 ));
    CascadeMux I__10617 (
            .O(N__46248),
            .I(N__46245));
    InMux I__10616 (
            .O(N__46245),
            .I(N__46242));
    LocalMux I__10615 (
            .O(N__46242),
            .I(N__46239));
    Span4Mux_h I__10614 (
            .O(N__46239),
            .I(N__46236));
    Span4Mux_v I__10613 (
            .O(N__46236),
            .I(N__46231));
    InMux I__10612 (
            .O(N__46235),
            .I(N__46228));
    InMux I__10611 (
            .O(N__46234),
            .I(N__46225));
    Span4Mux_h I__10610 (
            .O(N__46231),
            .I(N__46220));
    LocalMux I__10609 (
            .O(N__46228),
            .I(N__46220));
    LocalMux I__10608 (
            .O(N__46225),
            .I(N__46214));
    Span4Mux_h I__10607 (
            .O(N__46220),
            .I(N__46214));
    InMux I__10606 (
            .O(N__46219),
            .I(N__46211));
    Span4Mux_h I__10605 (
            .O(N__46214),
            .I(N__46208));
    LocalMux I__10604 (
            .O(N__46211),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__10603 (
            .O(N__46208),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__10602 (
            .O(N__46203),
            .I(N__46200));
    LocalMux I__10601 (
            .O(N__46200),
            .I(N__46197));
    Sp12to4 I__10600 (
            .O(N__46197),
            .I(N__46194));
    Span12Mux_h I__10599 (
            .O(N__46194),
            .I(N__46191));
    Span12Mux_v I__10598 (
            .O(N__46191),
            .I(N__46188));
    Odrv12 I__10597 (
            .O(N__46188),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__10596 (
            .O(N__46185),
            .I(N__46182));
    InMux I__10595 (
            .O(N__46182),
            .I(N__46179));
    LocalMux I__10594 (
            .O(N__46179),
            .I(N__46176));
    Span4Mux_h I__10593 (
            .O(N__46176),
            .I(N__46173));
    Span4Mux_h I__10592 (
            .O(N__46173),
            .I(N__46170));
    Odrv4 I__10591 (
            .O(N__46170),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    CascadeMux I__10590 (
            .O(N__46167),
            .I(N__46164));
    InMux I__10589 (
            .O(N__46164),
            .I(N__46161));
    LocalMux I__10588 (
            .O(N__46161),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    CascadeMux I__10587 (
            .O(N__46158),
            .I(N__46155));
    InMux I__10586 (
            .O(N__46155),
            .I(N__46152));
    LocalMux I__10585 (
            .O(N__46152),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ));
    InMux I__10584 (
            .O(N__46149),
            .I(N__46146));
    LocalMux I__10583 (
            .O(N__46146),
            .I(N__46143));
    Span4Mux_v I__10582 (
            .O(N__46143),
            .I(N__46140));
    Odrv4 I__10581 (
            .O(N__46140),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ));
    CascadeMux I__10580 (
            .O(N__46137),
            .I(N__46134));
    InMux I__10579 (
            .O(N__46134),
            .I(N__46131));
    LocalMux I__10578 (
            .O(N__46131),
            .I(N__46128));
    Span4Mux_v I__10577 (
            .O(N__46128),
            .I(N__46125));
    Odrv4 I__10576 (
            .O(N__46125),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt16 ));
    InMux I__10575 (
            .O(N__46122),
            .I(N__46119));
    LocalMux I__10574 (
            .O(N__46119),
            .I(N__46116));
    Odrv12 I__10573 (
            .O(N__46116),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ));
    CascadeMux I__10572 (
            .O(N__46113),
            .I(N__46110));
    InMux I__10571 (
            .O(N__46110),
            .I(N__46107));
    LocalMux I__10570 (
            .O(N__46107),
            .I(N__46104));
    Span4Mux_v I__10569 (
            .O(N__46104),
            .I(N__46101));
    Odrv4 I__10568 (
            .O(N__46101),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt18 ));
    InMux I__10567 (
            .O(N__46098),
            .I(N__46095));
    LocalMux I__10566 (
            .O(N__46095),
            .I(N__46092));
    Span4Mux_h I__10565 (
            .O(N__46092),
            .I(N__46089));
    Span4Mux_v I__10564 (
            .O(N__46089),
            .I(N__46086));
    Odrv4 I__10563 (
            .O(N__46086),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ));
    CascadeMux I__10562 (
            .O(N__46083),
            .I(N__46080));
    InMux I__10561 (
            .O(N__46080),
            .I(N__46077));
    LocalMux I__10560 (
            .O(N__46077),
            .I(N__46074));
    Span4Mux_h I__10559 (
            .O(N__46074),
            .I(N__46071));
    Span4Mux_v I__10558 (
            .O(N__46071),
            .I(N__46068));
    Odrv4 I__10557 (
            .O(N__46068),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt20 ));
    InMux I__10556 (
            .O(N__46065),
            .I(N__46062));
    LocalMux I__10555 (
            .O(N__46062),
            .I(N__46059));
    Odrv4 I__10554 (
            .O(N__46059),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ));
    CascadeMux I__10553 (
            .O(N__46056),
            .I(N__46053));
    InMux I__10552 (
            .O(N__46053),
            .I(N__46050));
    LocalMux I__10551 (
            .O(N__46050),
            .I(N__46047));
    Odrv4 I__10550 (
            .O(N__46047),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt24 ));
    InMux I__10549 (
            .O(N__46044),
            .I(N__46041));
    LocalMux I__10548 (
            .O(N__46041),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ));
    CascadeMux I__10547 (
            .O(N__46038),
            .I(N__46035));
    InMux I__10546 (
            .O(N__46035),
            .I(N__46032));
    LocalMux I__10545 (
            .O(N__46032),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt26 ));
    InMux I__10544 (
            .O(N__46029),
            .I(N__46026));
    LocalMux I__10543 (
            .O(N__46026),
            .I(N__46023));
    Span12Mux_h I__10542 (
            .O(N__46023),
            .I(N__46020));
    Odrv12 I__10541 (
            .O(N__46020),
            .I(\phase_controller_inst2.stoper_hc.un4_running_lt28 ));
    CascadeMux I__10540 (
            .O(N__46017),
            .I(N__46014));
    InMux I__10539 (
            .O(N__46014),
            .I(N__46011));
    LocalMux I__10538 (
            .O(N__46011),
            .I(N__46008));
    Span4Mux_h I__10537 (
            .O(N__46008),
            .I(N__46005));
    Span4Mux_v I__10536 (
            .O(N__46005),
            .I(N__46002));
    Span4Mux_v I__10535 (
            .O(N__46002),
            .I(N__45999));
    Odrv4 I__10534 (
            .O(N__45999),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ));
    InMux I__10533 (
            .O(N__45996),
            .I(N__45992));
    InMux I__10532 (
            .O(N__45995),
            .I(N__45989));
    LocalMux I__10531 (
            .O(N__45992),
            .I(N__45986));
    LocalMux I__10530 (
            .O(N__45989),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    Odrv4 I__10529 (
            .O(N__45986),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__10528 (
            .O(N__45981),
            .I(N__45978));
    InMux I__10527 (
            .O(N__45978),
            .I(N__45975));
    LocalMux I__10526 (
            .O(N__45975),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ));
    InMux I__10525 (
            .O(N__45972),
            .I(N__45969));
    LocalMux I__10524 (
            .O(N__45969),
            .I(N__45965));
    InMux I__10523 (
            .O(N__45968),
            .I(N__45962));
    Span4Mux_v I__10522 (
            .O(N__45965),
            .I(N__45959));
    LocalMux I__10521 (
            .O(N__45962),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    Odrv4 I__10520 (
            .O(N__45959),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__10519 (
            .O(N__45954),
            .I(N__45951));
    LocalMux I__10518 (
            .O(N__45951),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ));
    InMux I__10517 (
            .O(N__45948),
            .I(N__45944));
    InMux I__10516 (
            .O(N__45947),
            .I(N__45941));
    LocalMux I__10515 (
            .O(N__45944),
            .I(N__45938));
    LocalMux I__10514 (
            .O(N__45941),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    Odrv4 I__10513 (
            .O(N__45938),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ));
    InMux I__10512 (
            .O(N__45933),
            .I(N__45930));
    LocalMux I__10511 (
            .O(N__45930),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ));
    InMux I__10510 (
            .O(N__45927),
            .I(N__45924));
    LocalMux I__10509 (
            .O(N__45924),
            .I(N__45920));
    InMux I__10508 (
            .O(N__45923),
            .I(N__45917));
    Span4Mux_v I__10507 (
            .O(N__45920),
            .I(N__45914));
    LocalMux I__10506 (
            .O(N__45917),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    Odrv4 I__10505 (
            .O(N__45914),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__10504 (
            .O(N__45909),
            .I(N__45906));
    InMux I__10503 (
            .O(N__45906),
            .I(N__45903));
    LocalMux I__10502 (
            .O(N__45903),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ));
    InMux I__10501 (
            .O(N__45900),
            .I(N__45897));
    LocalMux I__10500 (
            .O(N__45897),
            .I(N__45894));
    Span4Mux_h I__10499 (
            .O(N__45894),
            .I(N__45891));
    Odrv4 I__10498 (
            .O(N__45891),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ));
    InMux I__10497 (
            .O(N__45888),
            .I(N__45884));
    InMux I__10496 (
            .O(N__45887),
            .I(N__45881));
    LocalMux I__10495 (
            .O(N__45884),
            .I(N__45878));
    LocalMux I__10494 (
            .O(N__45881),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    Odrv4 I__10493 (
            .O(N__45878),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ));
    CascadeMux I__10492 (
            .O(N__45873),
            .I(N__45870));
    InMux I__10491 (
            .O(N__45870),
            .I(N__45867));
    LocalMux I__10490 (
            .O(N__45867),
            .I(N__45864));
    Odrv4 I__10489 (
            .O(N__45864),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ));
    InMux I__10488 (
            .O(N__45861),
            .I(N__45857));
    InMux I__10487 (
            .O(N__45860),
            .I(N__45854));
    LocalMux I__10486 (
            .O(N__45857),
            .I(N__45851));
    LocalMux I__10485 (
            .O(N__45854),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    Odrv4 I__10484 (
            .O(N__45851),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__10483 (
            .O(N__45846),
            .I(N__45843));
    InMux I__10482 (
            .O(N__45843),
            .I(N__45840));
    LocalMux I__10481 (
            .O(N__45840),
            .I(N__45837));
    Span12Mux_v I__10480 (
            .O(N__45837),
            .I(N__45834));
    Odrv12 I__10479 (
            .O(N__45834),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ));
    InMux I__10478 (
            .O(N__45831),
            .I(N__45828));
    LocalMux I__10477 (
            .O(N__45828),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ));
    InMux I__10476 (
            .O(N__45825),
            .I(N__45821));
    InMux I__10475 (
            .O(N__45824),
            .I(N__45818));
    LocalMux I__10474 (
            .O(N__45821),
            .I(N__45815));
    LocalMux I__10473 (
            .O(N__45818),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    Odrv4 I__10472 (
            .O(N__45815),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ));
    InMux I__10471 (
            .O(N__45810),
            .I(N__45807));
    LocalMux I__10470 (
            .O(N__45807),
            .I(N__45804));
    Odrv12 I__10469 (
            .O(N__45804),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ));
    CascadeMux I__10468 (
            .O(N__45801),
            .I(N__45798));
    InMux I__10467 (
            .O(N__45798),
            .I(N__45795));
    LocalMux I__10466 (
            .O(N__45795),
            .I(N__45792));
    Odrv4 I__10465 (
            .O(N__45792),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ));
    InMux I__10464 (
            .O(N__45789),
            .I(N__45786));
    LocalMux I__10463 (
            .O(N__45786),
            .I(N__45783));
    Odrv12 I__10462 (
            .O(N__45783),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ));
    InMux I__10461 (
            .O(N__45780),
            .I(N__45776));
    InMux I__10460 (
            .O(N__45779),
            .I(N__45773));
    LocalMux I__10459 (
            .O(N__45776),
            .I(N__45770));
    LocalMux I__10458 (
            .O(N__45773),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    Odrv4 I__10457 (
            .O(N__45770),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__10456 (
            .O(N__45765),
            .I(N__45762));
    InMux I__10455 (
            .O(N__45762),
            .I(N__45759));
    LocalMux I__10454 (
            .O(N__45759),
            .I(N__45756));
    Odrv4 I__10453 (
            .O(N__45756),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ));
    InMux I__10452 (
            .O(N__45753),
            .I(N__45750));
    LocalMux I__10451 (
            .O(N__45750),
            .I(N__45746));
    InMux I__10450 (
            .O(N__45749),
            .I(N__45743));
    Span4Mux_v I__10449 (
            .O(N__45746),
            .I(N__45740));
    LocalMux I__10448 (
            .O(N__45743),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    Odrv4 I__10447 (
            .O(N__45740),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__10446 (
            .O(N__45735),
            .I(N__45732));
    InMux I__10445 (
            .O(N__45732),
            .I(N__45729));
    LocalMux I__10444 (
            .O(N__45729),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ));
    InMux I__10443 (
            .O(N__45726),
            .I(N__45723));
    LocalMux I__10442 (
            .O(N__45723),
            .I(N__45719));
    InMux I__10441 (
            .O(N__45722),
            .I(N__45716));
    Span4Mux_v I__10440 (
            .O(N__45719),
            .I(N__45713));
    LocalMux I__10439 (
            .O(N__45716),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    Odrv4 I__10438 (
            .O(N__45713),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__10437 (
            .O(N__45708),
            .I(N__45705));
    LocalMux I__10436 (
            .O(N__45705),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ));
    InMux I__10435 (
            .O(N__45702),
            .I(N__45699));
    LocalMux I__10434 (
            .O(N__45699),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ));
    InMux I__10433 (
            .O(N__45696),
            .I(N__45693));
    LocalMux I__10432 (
            .O(N__45693),
            .I(N__45689));
    InMux I__10431 (
            .O(N__45692),
            .I(N__45686));
    Span4Mux_v I__10430 (
            .O(N__45689),
            .I(N__45683));
    LocalMux I__10429 (
            .O(N__45686),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    Odrv4 I__10428 (
            .O(N__45683),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__10427 (
            .O(N__45678),
            .I(N__45675));
    InMux I__10426 (
            .O(N__45675),
            .I(N__45672));
    LocalMux I__10425 (
            .O(N__45672),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ));
    InMux I__10424 (
            .O(N__45669),
            .I(N__45665));
    InMux I__10423 (
            .O(N__45668),
            .I(N__45662));
    LocalMux I__10422 (
            .O(N__45665),
            .I(N__45659));
    LocalMux I__10421 (
            .O(N__45662),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    Odrv4 I__10420 (
            .O(N__45659),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ));
    InMux I__10419 (
            .O(N__45654),
            .I(N__45651));
    LocalMux I__10418 (
            .O(N__45651),
            .I(N__45648));
    Span4Mux_h I__10417 (
            .O(N__45648),
            .I(N__45645));
    Odrv4 I__10416 (
            .O(N__45645),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__10415 (
            .O(N__45642),
            .I(N__45639));
    InMux I__10414 (
            .O(N__45639),
            .I(N__45636));
    LocalMux I__10413 (
            .O(N__45636),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ));
    CascadeMux I__10412 (
            .O(N__45633),
            .I(N__45630));
    InMux I__10411 (
            .O(N__45630),
            .I(N__45627));
    LocalMux I__10410 (
            .O(N__45627),
            .I(N__45624));
    Span4Mux_h I__10409 (
            .O(N__45624),
            .I(N__45621));
    Odrv4 I__10408 (
            .O(N__45621),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ));
    InMux I__10407 (
            .O(N__45618),
            .I(N__45614));
    InMux I__10406 (
            .O(N__45617),
            .I(N__45611));
    LocalMux I__10405 (
            .O(N__45614),
            .I(N__45608));
    LocalMux I__10404 (
            .O(N__45611),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    Odrv4 I__10403 (
            .O(N__45608),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ));
    InMux I__10402 (
            .O(N__45603),
            .I(N__45600));
    LocalMux I__10401 (
            .O(N__45600),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ));
    CascadeMux I__10400 (
            .O(N__45597),
            .I(N__45594));
    InMux I__10399 (
            .O(N__45594),
            .I(N__45591));
    LocalMux I__10398 (
            .O(N__45591),
            .I(N__45588));
    Span4Mux_v I__10397 (
            .O(N__45588),
            .I(N__45585));
    Odrv4 I__10396 (
            .O(N__45585),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ));
    InMux I__10395 (
            .O(N__45582),
            .I(N__45578));
    InMux I__10394 (
            .O(N__45581),
            .I(N__45575));
    LocalMux I__10393 (
            .O(N__45578),
            .I(N__45572));
    LocalMux I__10392 (
            .O(N__45575),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    Odrv4 I__10391 (
            .O(N__45572),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ));
    InMux I__10390 (
            .O(N__45567),
            .I(N__45564));
    LocalMux I__10389 (
            .O(N__45564),
            .I(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ));
    InMux I__10388 (
            .O(N__45561),
            .I(N__45558));
    LocalMux I__10387 (
            .O(N__45558),
            .I(N__45554));
    InMux I__10386 (
            .O(N__45557),
            .I(N__45551));
    Odrv12 I__10385 (
            .O(N__45554),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__10384 (
            .O(N__45551),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    CascadeMux I__10383 (
            .O(N__45546),
            .I(elapsed_time_ns_1_RNI46CN9_0_17_cascade_));
    InMux I__10382 (
            .O(N__45543),
            .I(N__45537));
    InMux I__10381 (
            .O(N__45542),
            .I(N__45532));
    InMux I__10380 (
            .O(N__45541),
            .I(N__45532));
    InMux I__10379 (
            .O(N__45540),
            .I(N__45529));
    LocalMux I__10378 (
            .O(N__45537),
            .I(N__45526));
    LocalMux I__10377 (
            .O(N__45532),
            .I(N__45523));
    LocalMux I__10376 (
            .O(N__45529),
            .I(N__45520));
    Odrv12 I__10375 (
            .O(N__45526),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__10374 (
            .O(N__45523),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    Odrv4 I__10373 (
            .O(N__45520),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    CascadeMux I__10372 (
            .O(N__45513),
            .I(N__45510));
    InMux I__10371 (
            .O(N__45510),
            .I(N__45504));
    InMux I__10370 (
            .O(N__45509),
            .I(N__45504));
    LocalMux I__10369 (
            .O(N__45504),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ));
    InMux I__10368 (
            .O(N__45501),
            .I(N__45497));
    InMux I__10367 (
            .O(N__45500),
            .I(N__45494));
    LocalMux I__10366 (
            .O(N__45497),
            .I(N__45490));
    LocalMux I__10365 (
            .O(N__45494),
            .I(N__45487));
    InMux I__10364 (
            .O(N__45493),
            .I(N__45484));
    Span4Mux_h I__10363 (
            .O(N__45490),
            .I(N__45481));
    Span4Mux_v I__10362 (
            .O(N__45487),
            .I(N__45478));
    LocalMux I__10361 (
            .O(N__45484),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__10360 (
            .O(N__45481),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    Odrv4 I__10359 (
            .O(N__45478),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__10358 (
            .O(N__45471),
            .I(N__45467));
    InMux I__10357 (
            .O(N__45470),
            .I(N__45463));
    LocalMux I__10356 (
            .O(N__45467),
            .I(N__45459));
    InMux I__10355 (
            .O(N__45466),
            .I(N__45456));
    LocalMux I__10354 (
            .O(N__45463),
            .I(N__45453));
    InMux I__10353 (
            .O(N__45462),
            .I(N__45450));
    Span4Mux_v I__10352 (
            .O(N__45459),
            .I(N__45443));
    LocalMux I__10351 (
            .O(N__45456),
            .I(N__45443));
    Span4Mux_h I__10350 (
            .O(N__45453),
            .I(N__45443));
    LocalMux I__10349 (
            .O(N__45450),
            .I(N__45440));
    Odrv4 I__10348 (
            .O(N__45443),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    Odrv4 I__10347 (
            .O(N__45440),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__10346 (
            .O(N__45435),
            .I(N__45429));
    InMux I__10345 (
            .O(N__45434),
            .I(N__45429));
    LocalMux I__10344 (
            .O(N__45429),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ));
    InMux I__10343 (
            .O(N__45426),
            .I(N__45419));
    InMux I__10342 (
            .O(N__45425),
            .I(N__45419));
    InMux I__10341 (
            .O(N__45424),
            .I(N__45416));
    LocalMux I__10340 (
            .O(N__45419),
            .I(N__45412));
    LocalMux I__10339 (
            .O(N__45416),
            .I(N__45409));
    InMux I__10338 (
            .O(N__45415),
            .I(N__45406));
    Span4Mux_v I__10337 (
            .O(N__45412),
            .I(N__45403));
    Span4Mux_v I__10336 (
            .O(N__45409),
            .I(N__45398));
    LocalMux I__10335 (
            .O(N__45406),
            .I(N__45398));
    Odrv4 I__10334 (
            .O(N__45403),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    Odrv4 I__10333 (
            .O(N__45398),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__10332 (
            .O(N__45393),
            .I(N__45390));
    LocalMux I__10331 (
            .O(N__45390),
            .I(N__45387));
    Span4Mux_h I__10330 (
            .O(N__45387),
            .I(N__45384));
    Span4Mux_v I__10329 (
            .O(N__45384),
            .I(N__45380));
    InMux I__10328 (
            .O(N__45383),
            .I(N__45377));
    Odrv4 I__10327 (
            .O(N__45380),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__10326 (
            .O(N__45377),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    InMux I__10325 (
            .O(N__45372),
            .I(N__45369));
    LocalMux I__10324 (
            .O(N__45369),
            .I(N__45365));
    InMux I__10323 (
            .O(N__45368),
            .I(N__45361));
    Span4Mux_h I__10322 (
            .O(N__45365),
            .I(N__45358));
    InMux I__10321 (
            .O(N__45364),
            .I(N__45355));
    LocalMux I__10320 (
            .O(N__45361),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    Odrv4 I__10319 (
            .O(N__45358),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    LocalMux I__10318 (
            .O(N__45355),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__10317 (
            .O(N__45348),
            .I(N__45342));
    InMux I__10316 (
            .O(N__45347),
            .I(N__45339));
    InMux I__10315 (
            .O(N__45346),
            .I(N__45336));
    InMux I__10314 (
            .O(N__45345),
            .I(N__45333));
    LocalMux I__10313 (
            .O(N__45342),
            .I(N__45330));
    LocalMux I__10312 (
            .O(N__45339),
            .I(N__45327));
    LocalMux I__10311 (
            .O(N__45336),
            .I(N__45324));
    LocalMux I__10310 (
            .O(N__45333),
            .I(N__45321));
    Odrv4 I__10309 (
            .O(N__45330),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__10308 (
            .O(N__45327),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__10307 (
            .O(N__45324),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    Odrv4 I__10306 (
            .O(N__45321),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    CascadeMux I__10305 (
            .O(N__45312),
            .I(N__45307));
    InMux I__10304 (
            .O(N__45311),
            .I(N__45304));
    InMux I__10303 (
            .O(N__45310),
            .I(N__45299));
    InMux I__10302 (
            .O(N__45307),
            .I(N__45299));
    LocalMux I__10301 (
            .O(N__45304),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    LocalMux I__10300 (
            .O(N__45299),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ));
    InMux I__10299 (
            .O(N__45294),
            .I(N__45289));
    InMux I__10298 (
            .O(N__45293),
            .I(N__45284));
    InMux I__10297 (
            .O(N__45292),
            .I(N__45284));
    LocalMux I__10296 (
            .O(N__45289),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    LocalMux I__10295 (
            .O(N__45284),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__10294 (
            .O(N__45279),
            .I(N__45276));
    LocalMux I__10293 (
            .O(N__45276),
            .I(N__45271));
    InMux I__10292 (
            .O(N__45275),
            .I(N__45268));
    InMux I__10291 (
            .O(N__45274),
            .I(N__45265));
    Span4Mux_v I__10290 (
            .O(N__45271),
            .I(N__45262));
    LocalMux I__10289 (
            .O(N__45268),
            .I(N__45259));
    LocalMux I__10288 (
            .O(N__45265),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    Odrv4 I__10287 (
            .O(N__45262),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    Odrv4 I__10286 (
            .O(N__45259),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    InMux I__10285 (
            .O(N__45252),
            .I(N__45248));
    InMux I__10284 (
            .O(N__45251),
            .I(N__45243));
    LocalMux I__10283 (
            .O(N__45248),
            .I(N__45240));
    InMux I__10282 (
            .O(N__45247),
            .I(N__45235));
    InMux I__10281 (
            .O(N__45246),
            .I(N__45235));
    LocalMux I__10280 (
            .O(N__45243),
            .I(N__45232));
    Span4Mux_v I__10279 (
            .O(N__45240),
            .I(N__45227));
    LocalMux I__10278 (
            .O(N__45235),
            .I(N__45227));
    Odrv12 I__10277 (
            .O(N__45232),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    Odrv4 I__10276 (
            .O(N__45227),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__10275 (
            .O(N__45222),
            .I(N__45216));
    InMux I__10274 (
            .O(N__45221),
            .I(N__45216));
    LocalMux I__10273 (
            .O(N__45216),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__10272 (
            .O(N__45213),
            .I(N__45210));
    InMux I__10271 (
            .O(N__45210),
            .I(N__45205));
    InMux I__10270 (
            .O(N__45209),
            .I(N__45202));
    InMux I__10269 (
            .O(N__45208),
            .I(N__45199));
    LocalMux I__10268 (
            .O(N__45205),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__10267 (
            .O(N__45202),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    LocalMux I__10266 (
            .O(N__45199),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    CascadeMux I__10265 (
            .O(N__45192),
            .I(N__45187));
    InMux I__10264 (
            .O(N__45191),
            .I(N__45184));
    InMux I__10263 (
            .O(N__45190),
            .I(N__45180));
    InMux I__10262 (
            .O(N__45187),
            .I(N__45177));
    LocalMux I__10261 (
            .O(N__45184),
            .I(N__45174));
    InMux I__10260 (
            .O(N__45183),
            .I(N__45171));
    LocalMux I__10259 (
            .O(N__45180),
            .I(N__45168));
    LocalMux I__10258 (
            .O(N__45177),
            .I(N__45165));
    Span4Mux_h I__10257 (
            .O(N__45174),
            .I(N__45162));
    LocalMux I__10256 (
            .O(N__45171),
            .I(N__45159));
    Span4Mux_v I__10255 (
            .O(N__45168),
            .I(N__45156));
    Span4Mux_h I__10254 (
            .O(N__45165),
            .I(N__45153));
    Span4Mux_v I__10253 (
            .O(N__45162),
            .I(N__45148));
    Span4Mux_h I__10252 (
            .O(N__45159),
            .I(N__45148));
    Odrv4 I__10251 (
            .O(N__45156),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__10250 (
            .O(N__45153),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    Odrv4 I__10249 (
            .O(N__45148),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__10248 (
            .O(N__45141),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__10247 (
            .O(N__45138),
            .I(N__45135));
    InMux I__10246 (
            .O(N__45135),
            .I(N__45130));
    InMux I__10245 (
            .O(N__45134),
            .I(N__45127));
    InMux I__10244 (
            .O(N__45133),
            .I(N__45124));
    LocalMux I__10243 (
            .O(N__45130),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__10242 (
            .O(N__45127),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    LocalMux I__10241 (
            .O(N__45124),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__10240 (
            .O(N__45117),
            .I(bfn_18_13_0_));
    CascadeMux I__10239 (
            .O(N__45114),
            .I(N__45111));
    InMux I__10238 (
            .O(N__45111),
            .I(N__45106));
    InMux I__10237 (
            .O(N__45110),
            .I(N__45103));
    InMux I__10236 (
            .O(N__45109),
            .I(N__45100));
    LocalMux I__10235 (
            .O(N__45106),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__10234 (
            .O(N__45103),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    LocalMux I__10233 (
            .O(N__45100),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__10232 (
            .O(N__45093),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__10231 (
            .O(N__45090),
            .I(N__45086));
    InMux I__10230 (
            .O(N__45089),
            .I(N__45083));
    LocalMux I__10229 (
            .O(N__45086),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    LocalMux I__10228 (
            .O(N__45083),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    CascadeMux I__10227 (
            .O(N__45078),
            .I(N__45075));
    InMux I__10226 (
            .O(N__45075),
            .I(N__45070));
    InMux I__10225 (
            .O(N__45074),
            .I(N__45067));
    InMux I__10224 (
            .O(N__45073),
            .I(N__45064));
    LocalMux I__10223 (
            .O(N__45070),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__10222 (
            .O(N__45067),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    LocalMux I__10221 (
            .O(N__45064),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__10220 (
            .O(N__45057),
            .I(N__45052));
    InMux I__10219 (
            .O(N__45056),
            .I(N__45049));
    InMux I__10218 (
            .O(N__45055),
            .I(N__45046));
    LocalMux I__10217 (
            .O(N__45052),
            .I(N__45042));
    LocalMux I__10216 (
            .O(N__45049),
            .I(N__45037));
    LocalMux I__10215 (
            .O(N__45046),
            .I(N__45037));
    InMux I__10214 (
            .O(N__45045),
            .I(N__45034));
    Span4Mux_h I__10213 (
            .O(N__45042),
            .I(N__45027));
    Span4Mux_v I__10212 (
            .O(N__45037),
            .I(N__45027));
    LocalMux I__10211 (
            .O(N__45034),
            .I(N__45027));
    Span4Mux_h I__10210 (
            .O(N__45027),
            .I(N__45024));
    Odrv4 I__10209 (
            .O(N__45024),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__10208 (
            .O(N__45021),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__10207 (
            .O(N__45018),
            .I(N__45014));
    InMux I__10206 (
            .O(N__45017),
            .I(N__45011));
    LocalMux I__10205 (
            .O(N__45014),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    LocalMux I__10204 (
            .O(N__45011),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    CascadeMux I__10203 (
            .O(N__45006),
            .I(N__45003));
    InMux I__10202 (
            .O(N__45003),
            .I(N__44998));
    InMux I__10201 (
            .O(N__45002),
            .I(N__44995));
    InMux I__10200 (
            .O(N__45001),
            .I(N__44992));
    LocalMux I__10199 (
            .O(N__44998),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__10198 (
            .O(N__44995),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    LocalMux I__10197 (
            .O(N__44992),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__10196 (
            .O(N__44985),
            .I(N__44979));
    InMux I__10195 (
            .O(N__44984),
            .I(N__44976));
    InMux I__10194 (
            .O(N__44983),
            .I(N__44971));
    InMux I__10193 (
            .O(N__44982),
            .I(N__44971));
    LocalMux I__10192 (
            .O(N__44979),
            .I(N__44968));
    LocalMux I__10191 (
            .O(N__44976),
            .I(N__44965));
    LocalMux I__10190 (
            .O(N__44971),
            .I(N__44962));
    Span4Mux_h I__10189 (
            .O(N__44968),
            .I(N__44959));
    Span4Mux_v I__10188 (
            .O(N__44965),
            .I(N__44956));
    Span4Mux_h I__10187 (
            .O(N__44962),
            .I(N__44953));
    Odrv4 I__10186 (
            .O(N__44959),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__10185 (
            .O(N__44956),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    Odrv4 I__10184 (
            .O(N__44953),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__10183 (
            .O(N__44946),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__10182 (
            .O(N__44943),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    InMux I__10181 (
            .O(N__44940),
            .I(N__44937));
    LocalMux I__10180 (
            .O(N__44937),
            .I(N__44933));
    CascadeMux I__10179 (
            .O(N__44936),
            .I(N__44930));
    Span4Mux_v I__10178 (
            .O(N__44933),
            .I(N__44926));
    InMux I__10177 (
            .O(N__44930),
            .I(N__44923));
    InMux I__10176 (
            .O(N__44929),
            .I(N__44920));
    Odrv4 I__10175 (
            .O(N__44926),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__10174 (
            .O(N__44923),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__10173 (
            .O(N__44920),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__10172 (
            .O(N__44913),
            .I(N__44908));
    InMux I__10171 (
            .O(N__44912),
            .I(N__44903));
    InMux I__10170 (
            .O(N__44911),
            .I(N__44903));
    LocalMux I__10169 (
            .O(N__44908),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    LocalMux I__10168 (
            .O(N__44903),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__10167 (
            .O(N__44898),
            .I(N__44895));
    InMux I__10166 (
            .O(N__44895),
            .I(N__44888));
    InMux I__10165 (
            .O(N__44894),
            .I(N__44888));
    InMux I__10164 (
            .O(N__44893),
            .I(N__44885));
    LocalMux I__10163 (
            .O(N__44888),
            .I(N__44882));
    LocalMux I__10162 (
            .O(N__44885),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__10161 (
            .O(N__44882),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__10160 (
            .O(N__44877),
            .I(N__44874));
    InMux I__10159 (
            .O(N__44874),
            .I(N__44869));
    InMux I__10158 (
            .O(N__44873),
            .I(N__44866));
    InMux I__10157 (
            .O(N__44872),
            .I(N__44863));
    LocalMux I__10156 (
            .O(N__44869),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__10155 (
            .O(N__44866),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    LocalMux I__10154 (
            .O(N__44863),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__10153 (
            .O(N__44856),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__10152 (
            .O(N__44853),
            .I(N__44850));
    InMux I__10151 (
            .O(N__44850),
            .I(N__44845));
    InMux I__10150 (
            .O(N__44849),
            .I(N__44842));
    InMux I__10149 (
            .O(N__44848),
            .I(N__44839));
    LocalMux I__10148 (
            .O(N__44845),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__10147 (
            .O(N__44842),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    LocalMux I__10146 (
            .O(N__44839),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__10145 (
            .O(N__44832),
            .I(bfn_18_12_0_));
    CascadeMux I__10144 (
            .O(N__44829),
            .I(N__44826));
    InMux I__10143 (
            .O(N__44826),
            .I(N__44821));
    InMux I__10142 (
            .O(N__44825),
            .I(N__44818));
    InMux I__10141 (
            .O(N__44824),
            .I(N__44815));
    LocalMux I__10140 (
            .O(N__44821),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__10139 (
            .O(N__44818),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    LocalMux I__10138 (
            .O(N__44815),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    CascadeMux I__10137 (
            .O(N__44808),
            .I(N__44802));
    InMux I__10136 (
            .O(N__44807),
            .I(N__44799));
    InMux I__10135 (
            .O(N__44806),
            .I(N__44796));
    InMux I__10134 (
            .O(N__44805),
            .I(N__44793));
    InMux I__10133 (
            .O(N__44802),
            .I(N__44790));
    LocalMux I__10132 (
            .O(N__44799),
            .I(N__44781));
    LocalMux I__10131 (
            .O(N__44796),
            .I(N__44781));
    LocalMux I__10130 (
            .O(N__44793),
            .I(N__44781));
    LocalMux I__10129 (
            .O(N__44790),
            .I(N__44781));
    Span4Mux_v I__10128 (
            .O(N__44781),
            .I(N__44778));
    Odrv4 I__10127 (
            .O(N__44778),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__10126 (
            .O(N__44775),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__10125 (
            .O(N__44772),
            .I(N__44769));
    InMux I__10124 (
            .O(N__44769),
            .I(N__44764));
    InMux I__10123 (
            .O(N__44768),
            .I(N__44761));
    InMux I__10122 (
            .O(N__44767),
            .I(N__44758));
    LocalMux I__10121 (
            .O(N__44764),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__10120 (
            .O(N__44761),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    LocalMux I__10119 (
            .O(N__44758),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__10118 (
            .O(N__44751),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__10117 (
            .O(N__44748),
            .I(N__44745));
    InMux I__10116 (
            .O(N__44745),
            .I(N__44740));
    InMux I__10115 (
            .O(N__44744),
            .I(N__44737));
    InMux I__10114 (
            .O(N__44743),
            .I(N__44734));
    LocalMux I__10113 (
            .O(N__44740),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__10112 (
            .O(N__44737),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    LocalMux I__10111 (
            .O(N__44734),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__10110 (
            .O(N__44727),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__10109 (
            .O(N__44724),
            .I(N__44721));
    InMux I__10108 (
            .O(N__44721),
            .I(N__44716));
    InMux I__10107 (
            .O(N__44720),
            .I(N__44713));
    InMux I__10106 (
            .O(N__44719),
            .I(N__44710));
    LocalMux I__10105 (
            .O(N__44716),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__10104 (
            .O(N__44713),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    LocalMux I__10103 (
            .O(N__44710),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__10102 (
            .O(N__44703),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__10101 (
            .O(N__44700),
            .I(N__44697));
    InMux I__10100 (
            .O(N__44697),
            .I(N__44692));
    InMux I__10099 (
            .O(N__44696),
            .I(N__44689));
    InMux I__10098 (
            .O(N__44695),
            .I(N__44686));
    LocalMux I__10097 (
            .O(N__44692),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__10096 (
            .O(N__44689),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    LocalMux I__10095 (
            .O(N__44686),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__10094 (
            .O(N__44679),
            .I(N__44675));
    InMux I__10093 (
            .O(N__44678),
            .I(N__44672));
    LocalMux I__10092 (
            .O(N__44675),
            .I(N__44665));
    LocalMux I__10091 (
            .O(N__44672),
            .I(N__44665));
    InMux I__10090 (
            .O(N__44671),
            .I(N__44662));
    InMux I__10089 (
            .O(N__44670),
            .I(N__44659));
    Span4Mux_v I__10088 (
            .O(N__44665),
            .I(N__44654));
    LocalMux I__10087 (
            .O(N__44662),
            .I(N__44654));
    LocalMux I__10086 (
            .O(N__44659),
            .I(N__44651));
    Span4Mux_h I__10085 (
            .O(N__44654),
            .I(N__44648));
    Odrv4 I__10084 (
            .O(N__44651),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    Odrv4 I__10083 (
            .O(N__44648),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__10082 (
            .O(N__44643),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__10081 (
            .O(N__44640),
            .I(N__44637));
    InMux I__10080 (
            .O(N__44637),
            .I(N__44632));
    InMux I__10079 (
            .O(N__44636),
            .I(N__44629));
    InMux I__10078 (
            .O(N__44635),
            .I(N__44626));
    LocalMux I__10077 (
            .O(N__44632),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__10076 (
            .O(N__44629),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    LocalMux I__10075 (
            .O(N__44626),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    CascadeMux I__10074 (
            .O(N__44619),
            .I(N__44614));
    InMux I__10073 (
            .O(N__44618),
            .I(N__44610));
    InMux I__10072 (
            .O(N__44617),
            .I(N__44607));
    InMux I__10071 (
            .O(N__44614),
            .I(N__44604));
    InMux I__10070 (
            .O(N__44613),
            .I(N__44601));
    LocalMux I__10069 (
            .O(N__44610),
            .I(N__44596));
    LocalMux I__10068 (
            .O(N__44607),
            .I(N__44596));
    LocalMux I__10067 (
            .O(N__44604),
            .I(N__44593));
    LocalMux I__10066 (
            .O(N__44601),
            .I(N__44590));
    Span4Mux_h I__10065 (
            .O(N__44596),
            .I(N__44587));
    Span4Mux_h I__10064 (
            .O(N__44593),
            .I(N__44584));
    Odrv4 I__10063 (
            .O(N__44590),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__10062 (
            .O(N__44587),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    Odrv4 I__10061 (
            .O(N__44584),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__10060 (
            .O(N__44577),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__10059 (
            .O(N__44574),
            .I(N__44571));
    InMux I__10058 (
            .O(N__44571),
            .I(N__44566));
    InMux I__10057 (
            .O(N__44570),
            .I(N__44563));
    InMux I__10056 (
            .O(N__44569),
            .I(N__44560));
    LocalMux I__10055 (
            .O(N__44566),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__10054 (
            .O(N__44563),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    LocalMux I__10053 (
            .O(N__44560),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__10052 (
            .O(N__44553),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__10051 (
            .O(N__44550),
            .I(N__44547));
    InMux I__10050 (
            .O(N__44547),
            .I(N__44542));
    InMux I__10049 (
            .O(N__44546),
            .I(N__44539));
    InMux I__10048 (
            .O(N__44545),
            .I(N__44536));
    LocalMux I__10047 (
            .O(N__44542),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__10046 (
            .O(N__44539),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    LocalMux I__10045 (
            .O(N__44536),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__10044 (
            .O(N__44529),
            .I(bfn_18_11_0_));
    CascadeMux I__10043 (
            .O(N__44526),
            .I(N__44523));
    InMux I__10042 (
            .O(N__44523),
            .I(N__44518));
    InMux I__10041 (
            .O(N__44522),
            .I(N__44515));
    InMux I__10040 (
            .O(N__44521),
            .I(N__44512));
    LocalMux I__10039 (
            .O(N__44518),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__10038 (
            .O(N__44515),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    LocalMux I__10037 (
            .O(N__44512),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__10036 (
            .O(N__44505),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__10035 (
            .O(N__44502),
            .I(N__44499));
    InMux I__10034 (
            .O(N__44499),
            .I(N__44494));
    InMux I__10033 (
            .O(N__44498),
            .I(N__44491));
    InMux I__10032 (
            .O(N__44497),
            .I(N__44488));
    LocalMux I__10031 (
            .O(N__44494),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__10030 (
            .O(N__44491),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    LocalMux I__10029 (
            .O(N__44488),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__10028 (
            .O(N__44481),
            .I(N__44476));
    CascadeMux I__10027 (
            .O(N__44480),
            .I(N__44472));
    CascadeMux I__10026 (
            .O(N__44479),
            .I(N__44469));
    LocalMux I__10025 (
            .O(N__44476),
            .I(N__44466));
    InMux I__10024 (
            .O(N__44475),
            .I(N__44459));
    InMux I__10023 (
            .O(N__44472),
            .I(N__44459));
    InMux I__10022 (
            .O(N__44469),
            .I(N__44459));
    Span4Mux_v I__10021 (
            .O(N__44466),
            .I(N__44456));
    LocalMux I__10020 (
            .O(N__44459),
            .I(N__44453));
    Odrv4 I__10019 (
            .O(N__44456),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    Odrv4 I__10018 (
            .O(N__44453),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__10017 (
            .O(N__44448),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__10016 (
            .O(N__44445),
            .I(N__44442));
    InMux I__10015 (
            .O(N__44442),
            .I(N__44437));
    InMux I__10014 (
            .O(N__44441),
            .I(N__44434));
    InMux I__10013 (
            .O(N__44440),
            .I(N__44431));
    LocalMux I__10012 (
            .O(N__44437),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__10011 (
            .O(N__44434),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    LocalMux I__10010 (
            .O(N__44431),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__10009 (
            .O(N__44424),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    CascadeMux I__10008 (
            .O(N__44421),
            .I(N__44418));
    InMux I__10007 (
            .O(N__44418),
            .I(N__44413));
    InMux I__10006 (
            .O(N__44417),
            .I(N__44410));
    InMux I__10005 (
            .O(N__44416),
            .I(N__44407));
    LocalMux I__10004 (
            .O(N__44413),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__10003 (
            .O(N__44410),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    LocalMux I__10002 (
            .O(N__44407),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__10001 (
            .O(N__44400),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__10000 (
            .O(N__44397),
            .I(N__44394));
    InMux I__9999 (
            .O(N__44394),
            .I(N__44389));
    InMux I__9998 (
            .O(N__44393),
            .I(N__44386));
    InMux I__9997 (
            .O(N__44392),
            .I(N__44383));
    LocalMux I__9996 (
            .O(N__44389),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__9995 (
            .O(N__44386),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    LocalMux I__9994 (
            .O(N__44383),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__9993 (
            .O(N__44376),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__9992 (
            .O(N__44373),
            .I(N__44370));
    InMux I__9991 (
            .O(N__44370),
            .I(N__44365));
    InMux I__9990 (
            .O(N__44369),
            .I(N__44362));
    InMux I__9989 (
            .O(N__44368),
            .I(N__44359));
    LocalMux I__9988 (
            .O(N__44365),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__9987 (
            .O(N__44362),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    LocalMux I__9986 (
            .O(N__44359),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__9985 (
            .O(N__44352),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__9984 (
            .O(N__44349),
            .I(N__44346));
    LocalMux I__9983 (
            .O(N__44346),
            .I(N__44342));
    InMux I__9982 (
            .O(N__44345),
            .I(N__44339));
    Odrv4 I__9981 (
            .O(N__44342),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    LocalMux I__9980 (
            .O(N__44339),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    CascadeMux I__9979 (
            .O(N__44334),
            .I(elapsed_time_ns_1_RNI02CN9_0_13_cascade_));
    InMux I__9978 (
            .O(N__44331),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__9977 (
            .O(N__44328),
            .I(N__44325));
    InMux I__9976 (
            .O(N__44325),
            .I(N__44320));
    InMux I__9975 (
            .O(N__44324),
            .I(N__44317));
    InMux I__9974 (
            .O(N__44323),
            .I(N__44314));
    LocalMux I__9973 (
            .O(N__44320),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__9972 (
            .O(N__44317),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    LocalMux I__9971 (
            .O(N__44314),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__9970 (
            .O(N__44307),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__9969 (
            .O(N__44304),
            .I(N__44301));
    InMux I__9968 (
            .O(N__44301),
            .I(N__44296));
    InMux I__9967 (
            .O(N__44300),
            .I(N__44293));
    InMux I__9966 (
            .O(N__44299),
            .I(N__44290));
    LocalMux I__9965 (
            .O(N__44296),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__9964 (
            .O(N__44293),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    LocalMux I__9963 (
            .O(N__44290),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__9962 (
            .O(N__44283),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__9961 (
            .O(N__44280),
            .I(N__44277));
    InMux I__9960 (
            .O(N__44277),
            .I(N__44272));
    InMux I__9959 (
            .O(N__44276),
            .I(N__44269));
    InMux I__9958 (
            .O(N__44275),
            .I(N__44266));
    LocalMux I__9957 (
            .O(N__44272),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__9956 (
            .O(N__44269),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    LocalMux I__9955 (
            .O(N__44266),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__9954 (
            .O(N__44259),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9953 (
            .O(N__44256),
            .I(N__44253));
    InMux I__9952 (
            .O(N__44253),
            .I(N__44248));
    InMux I__9951 (
            .O(N__44252),
            .I(N__44245));
    InMux I__9950 (
            .O(N__44251),
            .I(N__44242));
    LocalMux I__9949 (
            .O(N__44248),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__9948 (
            .O(N__44245),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    LocalMux I__9947 (
            .O(N__44242),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__9946 (
            .O(N__44235),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__9945 (
            .O(N__44232),
            .I(N__44229));
    InMux I__9944 (
            .O(N__44229),
            .I(N__44224));
    InMux I__9943 (
            .O(N__44228),
            .I(N__44221));
    InMux I__9942 (
            .O(N__44227),
            .I(N__44218));
    LocalMux I__9941 (
            .O(N__44224),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__9940 (
            .O(N__44221),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    LocalMux I__9939 (
            .O(N__44218),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__9938 (
            .O(N__44211),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__9937 (
            .O(N__44208),
            .I(N__44205));
    InMux I__9936 (
            .O(N__44205),
            .I(N__44200));
    CascadeMux I__9935 (
            .O(N__44204),
            .I(N__44197));
    InMux I__9934 (
            .O(N__44203),
            .I(N__44194));
    LocalMux I__9933 (
            .O(N__44200),
            .I(N__44191));
    InMux I__9932 (
            .O(N__44197),
            .I(N__44188));
    LocalMux I__9931 (
            .O(N__44194),
            .I(N__44185));
    Span4Mux_v I__9930 (
            .O(N__44191),
            .I(N__44180));
    LocalMux I__9929 (
            .O(N__44188),
            .I(N__44180));
    Span12Mux_s4_v I__9928 (
            .O(N__44185),
            .I(N__44177));
    Span4Mux_h I__9927 (
            .O(N__44180),
            .I(N__44174));
    Odrv12 I__9926 (
            .O(N__44177),
            .I(\phase_controller_inst2.tr_time_passed ));
    Odrv4 I__9925 (
            .O(N__44174),
            .I(\phase_controller_inst2.tr_time_passed ));
    InMux I__9924 (
            .O(N__44169),
            .I(N__44165));
    InMux I__9923 (
            .O(N__44168),
            .I(N__44162));
    LocalMux I__9922 (
            .O(N__44165),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    LocalMux I__9921 (
            .O(N__44162),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ));
    CascadeMux I__9920 (
            .O(N__44157),
            .I(N__44154));
    InMux I__9919 (
            .O(N__44154),
            .I(N__44151));
    LocalMux I__9918 (
            .O(N__44151),
            .I(N__44148));
    Odrv12 I__9917 (
            .O(N__44148),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ));
    InMux I__9916 (
            .O(N__44145),
            .I(N__44141));
    CascadeMux I__9915 (
            .O(N__44144),
            .I(N__44138));
    LocalMux I__9914 (
            .O(N__44141),
            .I(N__44134));
    InMux I__9913 (
            .O(N__44138),
            .I(N__44131));
    CascadeMux I__9912 (
            .O(N__44137),
            .I(N__44128));
    Span4Mux_h I__9911 (
            .O(N__44134),
            .I(N__44121));
    LocalMux I__9910 (
            .O(N__44131),
            .I(N__44121));
    InMux I__9909 (
            .O(N__44128),
            .I(N__44118));
    InMux I__9908 (
            .O(N__44127),
            .I(N__44115));
    InMux I__9907 (
            .O(N__44126),
            .I(N__44112));
    Span4Mux_h I__9906 (
            .O(N__44121),
            .I(N__44107));
    LocalMux I__9905 (
            .O(N__44118),
            .I(N__44107));
    LocalMux I__9904 (
            .O(N__44115),
            .I(N__44104));
    LocalMux I__9903 (
            .O(N__44112),
            .I(N__44101));
    Span4Mux_h I__9902 (
            .O(N__44107),
            .I(N__44098));
    Span12Mux_h I__9901 (
            .O(N__44104),
            .I(N__44095));
    Span12Mux_v I__9900 (
            .O(N__44101),
            .I(N__44092));
    Span4Mux_v I__9899 (
            .O(N__44098),
            .I(N__44089));
    Odrv12 I__9898 (
            .O(N__44095),
            .I(\phase_controller_inst2.start_latched ));
    Odrv12 I__9897 (
            .O(N__44092),
            .I(\phase_controller_inst2.start_latched ));
    Odrv4 I__9896 (
            .O(N__44089),
            .I(\phase_controller_inst2.start_latched ));
    InMux I__9895 (
            .O(N__44082),
            .I(N__44078));
    InMux I__9894 (
            .O(N__44081),
            .I(N__44075));
    LocalMux I__9893 (
            .O(N__44078),
            .I(N__44069));
    LocalMux I__9892 (
            .O(N__44075),
            .I(N__44069));
    InMux I__9891 (
            .O(N__44074),
            .I(N__44066));
    Span4Mux_h I__9890 (
            .O(N__44069),
            .I(N__44063));
    LocalMux I__9889 (
            .O(N__44066),
            .I(\phase_controller_inst2.running ));
    Odrv4 I__9888 (
            .O(N__44063),
            .I(\phase_controller_inst2.running ));
    InMux I__9887 (
            .O(N__44058),
            .I(N__44052));
    InMux I__9886 (
            .O(N__44057),
            .I(N__44052));
    LocalMux I__9885 (
            .O(N__44052),
            .I(N__44049));
    Odrv12 I__9884 (
            .O(N__44049),
            .I(\phase_controller_inst2.N_39 ));
    CEMux I__9883 (
            .O(N__44046),
            .I(N__44043));
    LocalMux I__9882 (
            .O(N__44043),
            .I(N__44040));
    Odrv12 I__9881 (
            .O(N__44040),
            .I(\phase_controller_inst2.stoper_tr.N_39_0 ));
    InMux I__9880 (
            .O(N__44037),
            .I(N__44031));
    InMux I__9879 (
            .O(N__44036),
            .I(N__44031));
    LocalMux I__9878 (
            .O(N__44031),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ));
    InMux I__9877 (
            .O(N__44028),
            .I(N__44025));
    LocalMux I__9876 (
            .O(N__44025),
            .I(N__44022));
    Span4Mux_h I__9875 (
            .O(N__44022),
            .I(N__44019));
    Odrv4 I__9874 (
            .O(N__44019),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ));
    InMux I__9873 (
            .O(N__44016),
            .I(N__44013));
    LocalMux I__9872 (
            .O(N__44013),
            .I(N__44010));
    Span4Mux_v I__9871 (
            .O(N__44010),
            .I(N__44007));
    Odrv4 I__9870 (
            .O(N__44007),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ));
    InMux I__9869 (
            .O(N__44004),
            .I(N__44001));
    LocalMux I__9868 (
            .O(N__44001),
            .I(N__43998));
    Span4Mux_h I__9867 (
            .O(N__43998),
            .I(N__43995));
    Odrv4 I__9866 (
            .O(N__43995),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    CascadeMux I__9865 (
            .O(N__43992),
            .I(N__43989));
    InMux I__9864 (
            .O(N__43989),
            .I(N__43986));
    LocalMux I__9863 (
            .O(N__43986),
            .I(N__43983));
    Span4Mux_h I__9862 (
            .O(N__43983),
            .I(N__43980));
    Span4Mux_v I__9861 (
            .O(N__43980),
            .I(N__43974));
    InMux I__9860 (
            .O(N__43979),
            .I(N__43971));
    InMux I__9859 (
            .O(N__43978),
            .I(N__43968));
    CascadeMux I__9858 (
            .O(N__43977),
            .I(N__43965));
    Span4Mux_h I__9857 (
            .O(N__43974),
            .I(N__43962));
    LocalMux I__9856 (
            .O(N__43971),
            .I(N__43957));
    LocalMux I__9855 (
            .O(N__43968),
            .I(N__43957));
    InMux I__9854 (
            .O(N__43965),
            .I(N__43954));
    Span4Mux_h I__9853 (
            .O(N__43962),
            .I(N__43951));
    Span4Mux_h I__9852 (
            .O(N__43957),
            .I(N__43948));
    LocalMux I__9851 (
            .O(N__43954),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__9850 (
            .O(N__43951),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__9849 (
            .O(N__43948),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__9848 (
            .O(N__43941),
            .I(N__43938));
    LocalMux I__9847 (
            .O(N__43938),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__9846 (
            .O(N__43935),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__9845 (
            .O(N__43932),
            .I(N__43929));
    InMux I__9844 (
            .O(N__43929),
            .I(N__43926));
    LocalMux I__9843 (
            .O(N__43926),
            .I(N__43923));
    Span4Mux_h I__9842 (
            .O(N__43923),
            .I(N__43919));
    CascadeMux I__9841 (
            .O(N__43922),
            .I(N__43916));
    Span4Mux_v I__9840 (
            .O(N__43919),
            .I(N__43912));
    InMux I__9839 (
            .O(N__43916),
            .I(N__43909));
    InMux I__9838 (
            .O(N__43915),
            .I(N__43906));
    Span4Mux_h I__9837 (
            .O(N__43912),
            .I(N__43902));
    LocalMux I__9836 (
            .O(N__43909),
            .I(N__43897));
    LocalMux I__9835 (
            .O(N__43906),
            .I(N__43897));
    InMux I__9834 (
            .O(N__43905),
            .I(N__43894));
    Span4Mux_h I__9833 (
            .O(N__43902),
            .I(N__43891));
    Span4Mux_h I__9832 (
            .O(N__43897),
            .I(N__43888));
    LocalMux I__9831 (
            .O(N__43894),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__9830 (
            .O(N__43891),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__9829 (
            .O(N__43888),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__9828 (
            .O(N__43881),
            .I(N__43878));
    LocalMux I__9827 (
            .O(N__43878),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__9826 (
            .O(N__43875),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__9825 (
            .O(N__43872),
            .I(N__43869));
    InMux I__9824 (
            .O(N__43869),
            .I(N__43866));
    LocalMux I__9823 (
            .O(N__43866),
            .I(N__43862));
    CascadeMux I__9822 (
            .O(N__43865),
            .I(N__43859));
    Span4Mux_v I__9821 (
            .O(N__43862),
            .I(N__43856));
    InMux I__9820 (
            .O(N__43859),
            .I(N__43852));
    Span4Mux_h I__9819 (
            .O(N__43856),
            .I(N__43849));
    InMux I__9818 (
            .O(N__43855),
            .I(N__43846));
    LocalMux I__9817 (
            .O(N__43852),
            .I(N__43843));
    Span4Mux_h I__9816 (
            .O(N__43849),
            .I(N__43835));
    LocalMux I__9815 (
            .O(N__43846),
            .I(N__43835));
    Span4Mux_h I__9814 (
            .O(N__43843),
            .I(N__43835));
    InMux I__9813 (
            .O(N__43842),
            .I(N__43832));
    Span4Mux_h I__9812 (
            .O(N__43835),
            .I(N__43829));
    LocalMux I__9811 (
            .O(N__43832),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__9810 (
            .O(N__43829),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    CascadeMux I__9809 (
            .O(N__43824),
            .I(N__43821));
    InMux I__9808 (
            .O(N__43821),
            .I(N__43818));
    LocalMux I__9807 (
            .O(N__43818),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__9806 (
            .O(N__43815),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__9805 (
            .O(N__43812),
            .I(N__43809));
    InMux I__9804 (
            .O(N__43809),
            .I(N__43806));
    LocalMux I__9803 (
            .O(N__43806),
            .I(N__43803));
    Span4Mux_v I__9802 (
            .O(N__43803),
            .I(N__43798));
    CascadeMux I__9801 (
            .O(N__43802),
            .I(N__43795));
    InMux I__9800 (
            .O(N__43801),
            .I(N__43792));
    Span4Mux_v I__9799 (
            .O(N__43798),
            .I(N__43789));
    InMux I__9798 (
            .O(N__43795),
            .I(N__43786));
    LocalMux I__9797 (
            .O(N__43792),
            .I(N__43782));
    Span4Mux_h I__9796 (
            .O(N__43789),
            .I(N__43779));
    LocalMux I__9795 (
            .O(N__43786),
            .I(N__43776));
    InMux I__9794 (
            .O(N__43785),
            .I(N__43773));
    Span4Mux_v I__9793 (
            .O(N__43782),
            .I(N__43770));
    Span4Mux_h I__9792 (
            .O(N__43779),
            .I(N__43765));
    Span4Mux_v I__9791 (
            .O(N__43776),
            .I(N__43765));
    LocalMux I__9790 (
            .O(N__43773),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__9789 (
            .O(N__43770),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__9788 (
            .O(N__43765),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    CascadeMux I__9787 (
            .O(N__43758),
            .I(N__43755));
    InMux I__9786 (
            .O(N__43755),
            .I(N__43752));
    LocalMux I__9785 (
            .O(N__43752),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__9784 (
            .O(N__43749),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__9783 (
            .O(N__43746),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__9782 (
            .O(N__43743),
            .I(N__43740));
    LocalMux I__9781 (
            .O(N__43740),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ));
    InMux I__9780 (
            .O(N__43737),
            .I(N__43734));
    LocalMux I__9779 (
            .O(N__43734),
            .I(N__43731));
    Span4Mux_h I__9778 (
            .O(N__43731),
            .I(N__43728));
    Sp12to4 I__9777 (
            .O(N__43728),
            .I(N__43725));
    Span12Mux_v I__9776 (
            .O(N__43725),
            .I(N__43722));
    Span12Mux_h I__9775 (
            .O(N__43722),
            .I(N__43719));
    Odrv12 I__9774 (
            .O(N__43719),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    CascadeMux I__9773 (
            .O(N__43716),
            .I(N__43713));
    InMux I__9772 (
            .O(N__43713),
            .I(N__43710));
    LocalMux I__9771 (
            .O(N__43710),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ));
    InMux I__9770 (
            .O(N__43707),
            .I(N__43704));
    LocalMux I__9769 (
            .O(N__43704),
            .I(\phase_controller_inst1.stateZ0Z_5 ));
    IoInMux I__9768 (
            .O(N__43701),
            .I(N__43697));
    InMux I__9767 (
            .O(N__43700),
            .I(N__43694));
    LocalMux I__9766 (
            .O(N__43697),
            .I(test_c));
    LocalMux I__9765 (
            .O(N__43694),
            .I(test_c));
    InMux I__9764 (
            .O(N__43689),
            .I(N__43683));
    InMux I__9763 (
            .O(N__43688),
            .I(N__43683));
    LocalMux I__9762 (
            .O(N__43683),
            .I(N__43680));
    Span4Mux_s3_v I__9761 (
            .O(N__43680),
            .I(N__43677));
    Span4Mux_h I__9760 (
            .O(N__43677),
            .I(N__43673));
    CEMux I__9759 (
            .O(N__43676),
            .I(N__43670));
    Span4Mux_h I__9758 (
            .O(N__43673),
            .I(N__43664));
    LocalMux I__9757 (
            .O(N__43670),
            .I(N__43664));
    CEMux I__9756 (
            .O(N__43669),
            .I(N__43660));
    Span4Mux_h I__9755 (
            .O(N__43664),
            .I(N__43656));
    CEMux I__9754 (
            .O(N__43663),
            .I(N__43653));
    LocalMux I__9753 (
            .O(N__43660),
            .I(N__43650));
    CEMux I__9752 (
            .O(N__43659),
            .I(N__43647));
    Span4Mux_h I__9751 (
            .O(N__43656),
            .I(N__43642));
    LocalMux I__9750 (
            .O(N__43653),
            .I(N__43642));
    Span4Mux_s1_v I__9749 (
            .O(N__43650),
            .I(N__43638));
    LocalMux I__9748 (
            .O(N__43647),
            .I(N__43635));
    Span4Mux_v I__9747 (
            .O(N__43642),
            .I(N__43632));
    CEMux I__9746 (
            .O(N__43641),
            .I(N__43629));
    Span4Mux_v I__9745 (
            .O(N__43638),
            .I(N__43620));
    Span4Mux_h I__9744 (
            .O(N__43635),
            .I(N__43620));
    Span4Mux_v I__9743 (
            .O(N__43632),
            .I(N__43617));
    LocalMux I__9742 (
            .O(N__43629),
            .I(N__43614));
    CEMux I__9741 (
            .O(N__43628),
            .I(N__43611));
    CEMux I__9740 (
            .O(N__43627),
            .I(N__43608));
    InMux I__9739 (
            .O(N__43626),
            .I(N__43603));
    CEMux I__9738 (
            .O(N__43625),
            .I(N__43600));
    Sp12to4 I__9737 (
            .O(N__43620),
            .I(N__43596));
    Sp12to4 I__9736 (
            .O(N__43617),
            .I(N__43591));
    Sp12to4 I__9735 (
            .O(N__43614),
            .I(N__43591));
    LocalMux I__9734 (
            .O(N__43611),
            .I(N__43588));
    LocalMux I__9733 (
            .O(N__43608),
            .I(N__43585));
    CEMux I__9732 (
            .O(N__43607),
            .I(N__43582));
    InMux I__9731 (
            .O(N__43606),
            .I(N__43579));
    LocalMux I__9730 (
            .O(N__43603),
            .I(N__43574));
    LocalMux I__9729 (
            .O(N__43600),
            .I(N__43574));
    CEMux I__9728 (
            .O(N__43599),
            .I(N__43571));
    Span12Mux_s11_v I__9727 (
            .O(N__43596),
            .I(N__43566));
    Span12Mux_h I__9726 (
            .O(N__43591),
            .I(N__43566));
    Span4Mux_h I__9725 (
            .O(N__43588),
            .I(N__43559));
    Span4Mux_h I__9724 (
            .O(N__43585),
            .I(N__43559));
    LocalMux I__9723 (
            .O(N__43582),
            .I(N__43559));
    LocalMux I__9722 (
            .O(N__43579),
            .I(N__43556));
    Span4Mux_h I__9721 (
            .O(N__43574),
            .I(N__43553));
    LocalMux I__9720 (
            .O(N__43571),
            .I(N__43550));
    Span12Mux_v I__9719 (
            .O(N__43566),
            .I(N__43547));
    Span4Mux_h I__9718 (
            .O(N__43559),
            .I(N__43542));
    Span4Mux_h I__9717 (
            .O(N__43556),
            .I(N__43542));
    Sp12to4 I__9716 (
            .O(N__43553),
            .I(N__43539));
    Span4Mux_h I__9715 (
            .O(N__43550),
            .I(N__43536));
    Odrv12 I__9714 (
            .O(N__43547),
            .I(start_stop_c));
    Odrv4 I__9713 (
            .O(N__43542),
            .I(start_stop_c));
    Odrv12 I__9712 (
            .O(N__43539),
            .I(start_stop_c));
    Odrv4 I__9711 (
            .O(N__43536),
            .I(start_stop_c));
    CascadeMux I__9710 (
            .O(N__43527),
            .I(N__43524));
    InMux I__9709 (
            .O(N__43524),
            .I(N__43521));
    LocalMux I__9708 (
            .O(N__43521),
            .I(N__43518));
    Span4Mux_h I__9707 (
            .O(N__43518),
            .I(N__43515));
    Span4Mux_v I__9706 (
            .O(N__43515),
            .I(N__43509));
    InMux I__9705 (
            .O(N__43514),
            .I(N__43506));
    InMux I__9704 (
            .O(N__43513),
            .I(N__43503));
    InMux I__9703 (
            .O(N__43512),
            .I(N__43500));
    Sp12to4 I__9702 (
            .O(N__43509),
            .I(N__43495));
    LocalMux I__9701 (
            .O(N__43506),
            .I(N__43495));
    LocalMux I__9700 (
            .O(N__43503),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__9699 (
            .O(N__43500),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__9698 (
            .O(N__43495),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__9697 (
            .O(N__43488),
            .I(N__43485));
    InMux I__9696 (
            .O(N__43485),
            .I(N__43482));
    LocalMux I__9695 (
            .O(N__43482),
            .I(N__43479));
    Odrv4 I__9694 (
            .O(N__43479),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    InMux I__9693 (
            .O(N__43476),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    CascadeMux I__9692 (
            .O(N__43473),
            .I(N__43470));
    InMux I__9691 (
            .O(N__43470),
            .I(N__43467));
    LocalMux I__9690 (
            .O(N__43467),
            .I(N__43463));
    InMux I__9689 (
            .O(N__43466),
            .I(N__43458));
    Sp12to4 I__9688 (
            .O(N__43463),
            .I(N__43455));
    InMux I__9687 (
            .O(N__43462),
            .I(N__43452));
    InMux I__9686 (
            .O(N__43461),
            .I(N__43449));
    LocalMux I__9685 (
            .O(N__43458),
            .I(N__43446));
    Span12Mux_v I__9684 (
            .O(N__43455),
            .I(N__43443));
    LocalMux I__9683 (
            .O(N__43452),
            .I(N__43440));
    LocalMux I__9682 (
            .O(N__43449),
            .I(N__43437));
    Span4Mux_h I__9681 (
            .O(N__43446),
            .I(N__43434));
    Odrv12 I__9680 (
            .O(N__43443),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__9679 (
            .O(N__43440),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__9678 (
            .O(N__43437),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__9677 (
            .O(N__43434),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    InMux I__9676 (
            .O(N__43425),
            .I(N__43422));
    LocalMux I__9675 (
            .O(N__43422),
            .I(N__43419));
    Odrv4 I__9674 (
            .O(N__43419),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__9673 (
            .O(N__43416),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    InMux I__9672 (
            .O(N__43413),
            .I(N__43410));
    LocalMux I__9671 (
            .O(N__43410),
            .I(N__43407));
    Span4Mux_v I__9670 (
            .O(N__43407),
            .I(N__43404));
    Sp12to4 I__9669 (
            .O(N__43404),
            .I(N__43399));
    InMux I__9668 (
            .O(N__43403),
            .I(N__43396));
    InMux I__9667 (
            .O(N__43402),
            .I(N__43392));
    Span12Mux_h I__9666 (
            .O(N__43399),
            .I(N__43389));
    LocalMux I__9665 (
            .O(N__43396),
            .I(N__43386));
    InMux I__9664 (
            .O(N__43395),
            .I(N__43383));
    LocalMux I__9663 (
            .O(N__43392),
            .I(N__43380));
    Odrv12 I__9662 (
            .O(N__43389),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv4 I__9661 (
            .O(N__43386),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__9660 (
            .O(N__43383),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    Odrv12 I__9659 (
            .O(N__43380),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__9658 (
            .O(N__43371),
            .I(N__43368));
    LocalMux I__9657 (
            .O(N__43368),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__9656 (
            .O(N__43365),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    CascadeMux I__9655 (
            .O(N__43362),
            .I(N__43359));
    InMux I__9654 (
            .O(N__43359),
            .I(N__43355));
    CascadeMux I__9653 (
            .O(N__43358),
            .I(N__43352));
    LocalMux I__9652 (
            .O(N__43355),
            .I(N__43349));
    InMux I__9651 (
            .O(N__43352),
            .I(N__43345));
    Span4Mux_v I__9650 (
            .O(N__43349),
            .I(N__43342));
    CascadeMux I__9649 (
            .O(N__43348),
            .I(N__43339));
    LocalMux I__9648 (
            .O(N__43345),
            .I(N__43336));
    Sp12to4 I__9647 (
            .O(N__43342),
            .I(N__43332));
    InMux I__9646 (
            .O(N__43339),
            .I(N__43329));
    Span4Mux_v I__9645 (
            .O(N__43336),
            .I(N__43326));
    InMux I__9644 (
            .O(N__43335),
            .I(N__43323));
    Span12Mux_h I__9643 (
            .O(N__43332),
            .I(N__43320));
    LocalMux I__9642 (
            .O(N__43329),
            .I(N__43317));
    Span4Mux_h I__9641 (
            .O(N__43326),
            .I(N__43314));
    LocalMux I__9640 (
            .O(N__43323),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv12 I__9639 (
            .O(N__43320),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__9638 (
            .O(N__43317),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__9637 (
            .O(N__43314),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__9636 (
            .O(N__43305),
            .I(N__43302));
    LocalMux I__9635 (
            .O(N__43302),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__9634 (
            .O(N__43299),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__9633 (
            .O(N__43296),
            .I(N__43293));
    InMux I__9632 (
            .O(N__43293),
            .I(N__43290));
    LocalMux I__9631 (
            .O(N__43290),
            .I(N__43287));
    Span4Mux_h I__9630 (
            .O(N__43287),
            .I(N__43283));
    InMux I__9629 (
            .O(N__43286),
            .I(N__43279));
    Span4Mux_v I__9628 (
            .O(N__43283),
            .I(N__43276));
    InMux I__9627 (
            .O(N__43282),
            .I(N__43273));
    LocalMux I__9626 (
            .O(N__43279),
            .I(N__43269));
    Span4Mux_h I__9625 (
            .O(N__43276),
            .I(N__43264));
    LocalMux I__9624 (
            .O(N__43273),
            .I(N__43264));
    InMux I__9623 (
            .O(N__43272),
            .I(N__43261));
    Span4Mux_v I__9622 (
            .O(N__43269),
            .I(N__43256));
    Span4Mux_h I__9621 (
            .O(N__43264),
            .I(N__43256));
    LocalMux I__9620 (
            .O(N__43261),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    Odrv4 I__9619 (
            .O(N__43256),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__9618 (
            .O(N__43251),
            .I(N__43248));
    LocalMux I__9617 (
            .O(N__43248),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__9616 (
            .O(N__43245),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__9615 (
            .O(N__43242),
            .I(N__43239));
    InMux I__9614 (
            .O(N__43239),
            .I(N__43236));
    LocalMux I__9613 (
            .O(N__43236),
            .I(N__43233));
    Span4Mux_v I__9612 (
            .O(N__43233),
            .I(N__43228));
    CascadeMux I__9611 (
            .O(N__43232),
            .I(N__43225));
    InMux I__9610 (
            .O(N__43231),
            .I(N__43222));
    Span4Mux_h I__9609 (
            .O(N__43228),
            .I(N__43219));
    InMux I__9608 (
            .O(N__43225),
            .I(N__43215));
    LocalMux I__9607 (
            .O(N__43222),
            .I(N__43212));
    Span4Mux_h I__9606 (
            .O(N__43219),
            .I(N__43209));
    InMux I__9605 (
            .O(N__43218),
            .I(N__43206));
    LocalMux I__9604 (
            .O(N__43215),
            .I(N__43203));
    Span4Mux_v I__9603 (
            .O(N__43212),
            .I(N__43200));
    Span4Mux_h I__9602 (
            .O(N__43209),
            .I(N__43197));
    LocalMux I__9601 (
            .O(N__43206),
            .I(N__43190));
    Span4Mux_v I__9600 (
            .O(N__43203),
            .I(N__43190));
    Span4Mux_h I__9599 (
            .O(N__43200),
            .I(N__43190));
    Odrv4 I__9598 (
            .O(N__43197),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    Odrv4 I__9597 (
            .O(N__43190),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    CascadeMux I__9596 (
            .O(N__43185),
            .I(N__43182));
    InMux I__9595 (
            .O(N__43182),
            .I(N__43179));
    LocalMux I__9594 (
            .O(N__43179),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__9593 (
            .O(N__43176),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__9592 (
            .O(N__43173),
            .I(N__43170));
    InMux I__9591 (
            .O(N__43170),
            .I(N__43167));
    LocalMux I__9590 (
            .O(N__43167),
            .I(N__43162));
    InMux I__9589 (
            .O(N__43166),
            .I(N__43159));
    InMux I__9588 (
            .O(N__43165),
            .I(N__43156));
    Sp12to4 I__9587 (
            .O(N__43162),
            .I(N__43152));
    LocalMux I__9586 (
            .O(N__43159),
            .I(N__43147));
    LocalMux I__9585 (
            .O(N__43156),
            .I(N__43147));
    InMux I__9584 (
            .O(N__43155),
            .I(N__43144));
    Span12Mux_v I__9583 (
            .O(N__43152),
            .I(N__43141));
    Span4Mux_h I__9582 (
            .O(N__43147),
            .I(N__43138));
    LocalMux I__9581 (
            .O(N__43144),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv12 I__9580 (
            .O(N__43141),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    Odrv4 I__9579 (
            .O(N__43138),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    CascadeMux I__9578 (
            .O(N__43131),
            .I(N__43128));
    InMux I__9577 (
            .O(N__43128),
            .I(N__43125));
    LocalMux I__9576 (
            .O(N__43125),
            .I(N__43122));
    Odrv4 I__9575 (
            .O(N__43122),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__9574 (
            .O(N__43119),
            .I(bfn_17_23_0_));
    CascadeMux I__9573 (
            .O(N__43116),
            .I(N__43113));
    InMux I__9572 (
            .O(N__43113),
            .I(N__43110));
    LocalMux I__9571 (
            .O(N__43110),
            .I(N__43107));
    Span4Mux_v I__9570 (
            .O(N__43107),
            .I(N__43103));
    InMux I__9569 (
            .O(N__43106),
            .I(N__43100));
    Span4Mux_h I__9568 (
            .O(N__43103),
            .I(N__43097));
    LocalMux I__9567 (
            .O(N__43100),
            .I(N__43093));
    Span4Mux_h I__9566 (
            .O(N__43097),
            .I(N__43089));
    InMux I__9565 (
            .O(N__43096),
            .I(N__43086));
    Span4Mux_v I__9564 (
            .O(N__43093),
            .I(N__43083));
    InMux I__9563 (
            .O(N__43092),
            .I(N__43080));
    Span4Mux_h I__9562 (
            .O(N__43089),
            .I(N__43077));
    LocalMux I__9561 (
            .O(N__43086),
            .I(N__43074));
    Span4Mux_h I__9560 (
            .O(N__43083),
            .I(N__43071));
    LocalMux I__9559 (
            .O(N__43080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__9558 (
            .O(N__43077),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__9557 (
            .O(N__43074),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    Odrv4 I__9556 (
            .O(N__43071),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__9555 (
            .O(N__43062),
            .I(N__43059));
    LocalMux I__9554 (
            .O(N__43059),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__9553 (
            .O(N__43056),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__9552 (
            .O(N__43053),
            .I(N__43050));
    InMux I__9551 (
            .O(N__43050),
            .I(N__43047));
    LocalMux I__9550 (
            .O(N__43047),
            .I(N__43044));
    Span4Mux_h I__9549 (
            .O(N__43044),
            .I(N__43041));
    Span4Mux_h I__9548 (
            .O(N__43041),
            .I(N__43038));
    Odrv4 I__9547 (
            .O(N__43038),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__9546 (
            .O(N__43035),
            .I(N__43032));
    LocalMux I__9545 (
            .O(N__43032),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__9544 (
            .O(N__43029),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__9543 (
            .O(N__43026),
            .I(N__43023));
    InMux I__9542 (
            .O(N__43023),
            .I(N__43020));
    LocalMux I__9541 (
            .O(N__43020),
            .I(N__43017));
    Span4Mux_h I__9540 (
            .O(N__43017),
            .I(N__43014));
    Span4Mux_h I__9539 (
            .O(N__43014),
            .I(N__43011));
    Odrv4 I__9538 (
            .O(N__43011),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__9537 (
            .O(N__43008),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    CascadeMux I__9536 (
            .O(N__43005),
            .I(N__43002));
    InMux I__9535 (
            .O(N__43002),
            .I(N__42999));
    LocalMux I__9534 (
            .O(N__42999),
            .I(N__42996));
    Span4Mux_v I__9533 (
            .O(N__42996),
            .I(N__42993));
    Sp12to4 I__9532 (
            .O(N__42993),
            .I(N__42990));
    Odrv12 I__9531 (
            .O(N__42990),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__9530 (
            .O(N__42987),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    InMux I__9529 (
            .O(N__42984),
            .I(N__42981));
    LocalMux I__9528 (
            .O(N__42981),
            .I(N__42978));
    Span4Mux_h I__9527 (
            .O(N__42978),
            .I(N__42974));
    InMux I__9526 (
            .O(N__42977),
            .I(N__42971));
    Span4Mux_v I__9525 (
            .O(N__42974),
            .I(N__42968));
    LocalMux I__9524 (
            .O(N__42971),
            .I(N__42965));
    Span4Mux_h I__9523 (
            .O(N__42968),
            .I(N__42960));
    Span4Mux_h I__9522 (
            .O(N__42965),
            .I(N__42960));
    Span4Mux_h I__9521 (
            .O(N__42960),
            .I(N__42955));
    InMux I__9520 (
            .O(N__42959),
            .I(N__42952));
    InMux I__9519 (
            .O(N__42958),
            .I(N__42949));
    Odrv4 I__9518 (
            .O(N__42955),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__9517 (
            .O(N__42952),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__9516 (
            .O(N__42949),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    CascadeMux I__9515 (
            .O(N__42942),
            .I(N__42939));
    InMux I__9514 (
            .O(N__42939),
            .I(N__42936));
    LocalMux I__9513 (
            .O(N__42936),
            .I(N__42933));
    Span4Mux_v I__9512 (
            .O(N__42933),
            .I(N__42930));
    Span4Mux_h I__9511 (
            .O(N__42930),
            .I(N__42927));
    Odrv4 I__9510 (
            .O(N__42927),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__9509 (
            .O(N__42924),
            .I(N__42921));
    LocalMux I__9508 (
            .O(N__42921),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__9507 (
            .O(N__42918),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__9506 (
            .O(N__42915),
            .I(N__42912));
    InMux I__9505 (
            .O(N__42912),
            .I(N__42909));
    LocalMux I__9504 (
            .O(N__42909),
            .I(N__42906));
    Span4Mux_h I__9503 (
            .O(N__42906),
            .I(N__42902));
    InMux I__9502 (
            .O(N__42905),
            .I(N__42899));
    Span4Mux_v I__9501 (
            .O(N__42902),
            .I(N__42894));
    LocalMux I__9500 (
            .O(N__42899),
            .I(N__42894));
    Span4Mux_h I__9499 (
            .O(N__42894),
            .I(N__42889));
    InMux I__9498 (
            .O(N__42893),
            .I(N__42886));
    InMux I__9497 (
            .O(N__42892),
            .I(N__42883));
    Span4Mux_h I__9496 (
            .O(N__42889),
            .I(N__42880));
    LocalMux I__9495 (
            .O(N__42886),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    LocalMux I__9494 (
            .O(N__42883),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__9493 (
            .O(N__42880),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    CascadeMux I__9492 (
            .O(N__42873),
            .I(N__42870));
    InMux I__9491 (
            .O(N__42870),
            .I(N__42867));
    LocalMux I__9490 (
            .O(N__42867),
            .I(N__42864));
    Span4Mux_h I__9489 (
            .O(N__42864),
            .I(N__42861));
    Span4Mux_h I__9488 (
            .O(N__42861),
            .I(N__42858));
    Odrv4 I__9487 (
            .O(N__42858),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__9486 (
            .O(N__42855),
            .I(N__42852));
    LocalMux I__9485 (
            .O(N__42852),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__9484 (
            .O(N__42849),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__9483 (
            .O(N__42846),
            .I(N__42843));
    InMux I__9482 (
            .O(N__42843),
            .I(N__42840));
    LocalMux I__9481 (
            .O(N__42840),
            .I(N__42837));
    Span4Mux_v I__9480 (
            .O(N__42837),
            .I(N__42832));
    InMux I__9479 (
            .O(N__42836),
            .I(N__42829));
    InMux I__9478 (
            .O(N__42835),
            .I(N__42826));
    Sp12to4 I__9477 (
            .O(N__42832),
            .I(N__42822));
    LocalMux I__9476 (
            .O(N__42829),
            .I(N__42819));
    LocalMux I__9475 (
            .O(N__42826),
            .I(N__42816));
    InMux I__9474 (
            .O(N__42825),
            .I(N__42813));
    Span12Mux_h I__9473 (
            .O(N__42822),
            .I(N__42810));
    Span12Mux_h I__9472 (
            .O(N__42819),
            .I(N__42807));
    Odrv4 I__9471 (
            .O(N__42816),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__9470 (
            .O(N__42813),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv12 I__9469 (
            .O(N__42810),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    Odrv12 I__9468 (
            .O(N__42807),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    CascadeMux I__9467 (
            .O(N__42798),
            .I(N__42795));
    InMux I__9466 (
            .O(N__42795),
            .I(N__42792));
    LocalMux I__9465 (
            .O(N__42792),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__9464 (
            .O(N__42789),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    CascadeMux I__9463 (
            .O(N__42786),
            .I(N__42783));
    InMux I__9462 (
            .O(N__42783),
            .I(N__42780));
    LocalMux I__9461 (
            .O(N__42780),
            .I(N__42777));
    Span4Mux_h I__9460 (
            .O(N__42777),
            .I(N__42773));
    InMux I__9459 (
            .O(N__42776),
            .I(N__42769));
    Span4Mux_v I__9458 (
            .O(N__42773),
            .I(N__42766));
    InMux I__9457 (
            .O(N__42772),
            .I(N__42763));
    LocalMux I__9456 (
            .O(N__42769),
            .I(N__42759));
    Span4Mux_h I__9455 (
            .O(N__42766),
            .I(N__42754));
    LocalMux I__9454 (
            .O(N__42763),
            .I(N__42754));
    InMux I__9453 (
            .O(N__42762),
            .I(N__42751));
    Span4Mux_v I__9452 (
            .O(N__42759),
            .I(N__42746));
    Span4Mux_h I__9451 (
            .O(N__42754),
            .I(N__42746));
    LocalMux I__9450 (
            .O(N__42751),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__9449 (
            .O(N__42746),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__9448 (
            .O(N__42741),
            .I(N__42738));
    LocalMux I__9447 (
            .O(N__42738),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__9446 (
            .O(N__42735),
            .I(bfn_17_22_0_));
    CascadeMux I__9445 (
            .O(N__42732),
            .I(N__42729));
    InMux I__9444 (
            .O(N__42729),
            .I(N__42726));
    LocalMux I__9443 (
            .O(N__42726),
            .I(N__42723));
    Span4Mux_h I__9442 (
            .O(N__42723),
            .I(N__42720));
    Span4Mux_v I__9441 (
            .O(N__42720),
            .I(N__42714));
    InMux I__9440 (
            .O(N__42719),
            .I(N__42711));
    InMux I__9439 (
            .O(N__42718),
            .I(N__42708));
    InMux I__9438 (
            .O(N__42717),
            .I(N__42705));
    Span4Mux_h I__9437 (
            .O(N__42714),
            .I(N__42700));
    LocalMux I__9436 (
            .O(N__42711),
            .I(N__42700));
    LocalMux I__9435 (
            .O(N__42708),
            .I(N__42697));
    LocalMux I__9434 (
            .O(N__42705),
            .I(N__42694));
    Span4Mux_h I__9433 (
            .O(N__42700),
            .I(N__42691));
    Odrv4 I__9432 (
            .O(N__42697),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__9431 (
            .O(N__42694),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    Odrv4 I__9430 (
            .O(N__42691),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    CascadeMux I__9429 (
            .O(N__42684),
            .I(N__42681));
    InMux I__9428 (
            .O(N__42681),
            .I(N__42678));
    LocalMux I__9427 (
            .O(N__42678),
            .I(N__42675));
    Odrv4 I__9426 (
            .O(N__42675),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__9425 (
            .O(N__42672),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__9424 (
            .O(N__42669),
            .I(N__42666));
    InMux I__9423 (
            .O(N__42666),
            .I(N__42663));
    LocalMux I__9422 (
            .O(N__42663),
            .I(N__42660));
    Span4Mux_v I__9421 (
            .O(N__42660),
            .I(N__42656));
    InMux I__9420 (
            .O(N__42659),
            .I(N__42651));
    Span4Mux_v I__9419 (
            .O(N__42656),
            .I(N__42648));
    InMux I__9418 (
            .O(N__42655),
            .I(N__42645));
    InMux I__9417 (
            .O(N__42654),
            .I(N__42642));
    LocalMux I__9416 (
            .O(N__42651),
            .I(N__42639));
    Span4Mux_h I__9415 (
            .O(N__42648),
            .I(N__42636));
    LocalMux I__9414 (
            .O(N__42645),
            .I(N__42633));
    LocalMux I__9413 (
            .O(N__42642),
            .I(N__42630));
    Span4Mux_h I__9412 (
            .O(N__42639),
            .I(N__42623));
    Span4Mux_h I__9411 (
            .O(N__42636),
            .I(N__42623));
    Span4Mux_h I__9410 (
            .O(N__42633),
            .I(N__42623));
    Odrv4 I__9409 (
            .O(N__42630),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__9408 (
            .O(N__42623),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    CascadeMux I__9407 (
            .O(N__42618),
            .I(N__42615));
    InMux I__9406 (
            .O(N__42615),
            .I(N__42612));
    LocalMux I__9405 (
            .O(N__42612),
            .I(N__42609));
    Span4Mux_h I__9404 (
            .O(N__42609),
            .I(N__42606));
    Span4Mux_h I__9403 (
            .O(N__42606),
            .I(N__42603));
    Odrv4 I__9402 (
            .O(N__42603),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    CascadeMux I__9401 (
            .O(N__42600),
            .I(N__42597));
    InMux I__9400 (
            .O(N__42597),
            .I(N__42594));
    LocalMux I__9399 (
            .O(N__42594),
            .I(N__42591));
    Span4Mux_v I__9398 (
            .O(N__42591),
            .I(N__42588));
    Odrv4 I__9397 (
            .O(N__42588),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__9396 (
            .O(N__42585),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__9395 (
            .O(N__42582),
            .I(N__42579));
    LocalMux I__9394 (
            .O(N__42579),
            .I(N__42576));
    Span12Mux_v I__9393 (
            .O(N__42576),
            .I(N__42573));
    Odrv12 I__9392 (
            .O(N__42573),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__9391 (
            .O(N__42570),
            .I(N__42565));
    CascadeMux I__9390 (
            .O(N__42569),
            .I(N__42562));
    InMux I__9389 (
            .O(N__42568),
            .I(N__42558));
    LocalMux I__9388 (
            .O(N__42565),
            .I(N__42555));
    InMux I__9387 (
            .O(N__42562),
            .I(N__42552));
    InMux I__9386 (
            .O(N__42561),
            .I(N__42549));
    LocalMux I__9385 (
            .O(N__42558),
            .I(N__42546));
    Span4Mux_h I__9384 (
            .O(N__42555),
            .I(N__42543));
    LocalMux I__9383 (
            .O(N__42552),
            .I(N__42538));
    LocalMux I__9382 (
            .O(N__42549),
            .I(N__42538));
    Span4Mux_h I__9381 (
            .O(N__42546),
            .I(N__42535));
    Span4Mux_h I__9380 (
            .O(N__42543),
            .I(N__42532));
    Span12Mux_h I__9379 (
            .O(N__42538),
            .I(N__42529));
    Span4Mux_v I__9378 (
            .O(N__42535),
            .I(N__42524));
    Span4Mux_h I__9377 (
            .O(N__42532),
            .I(N__42524));
    Odrv12 I__9376 (
            .O(N__42529),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__9375 (
            .O(N__42524),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__9374 (
            .O(N__42519),
            .I(N__42516));
    LocalMux I__9373 (
            .O(N__42516),
            .I(N__42513));
    Span12Mux_s9_h I__9372 (
            .O(N__42513),
            .I(N__42510));
    Odrv12 I__9371 (
            .O(N__42510),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__9370 (
            .O(N__42507),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__9369 (
            .O(N__42504),
            .I(N__42501));
    InMux I__9368 (
            .O(N__42501),
            .I(N__42498));
    LocalMux I__9367 (
            .O(N__42498),
            .I(N__42495));
    Span4Mux_v I__9366 (
            .O(N__42495),
            .I(N__42492));
    Span4Mux_h I__9365 (
            .O(N__42492),
            .I(N__42489));
    Odrv4 I__9364 (
            .O(N__42489),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__9363 (
            .O(N__42486),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__9362 (
            .O(N__42483),
            .I(N__42480));
    InMux I__9361 (
            .O(N__42480),
            .I(N__42477));
    LocalMux I__9360 (
            .O(N__42477),
            .I(N__42474));
    Span4Mux_h I__9359 (
            .O(N__42474),
            .I(N__42471));
    Span4Mux_h I__9358 (
            .O(N__42471),
            .I(N__42468));
    Odrv4 I__9357 (
            .O(N__42468),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__9356 (
            .O(N__42465),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__9355 (
            .O(N__42462),
            .I(N__42459));
    InMux I__9354 (
            .O(N__42459),
            .I(N__42453));
    InMux I__9353 (
            .O(N__42458),
            .I(N__42450));
    InMux I__9352 (
            .O(N__42457),
            .I(N__42447));
    InMux I__9351 (
            .O(N__42456),
            .I(N__42444));
    LocalMux I__9350 (
            .O(N__42453),
            .I(N__42441));
    LocalMux I__9349 (
            .O(N__42450),
            .I(N__42438));
    LocalMux I__9348 (
            .O(N__42447),
            .I(N__42433));
    LocalMux I__9347 (
            .O(N__42444),
            .I(N__42433));
    Span12Mux_h I__9346 (
            .O(N__42441),
            .I(N__42430));
    Span4Mux_v I__9345 (
            .O(N__42438),
            .I(N__42425));
    Span4Mux_v I__9344 (
            .O(N__42433),
            .I(N__42425));
    Odrv12 I__9343 (
            .O(N__42430),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__9342 (
            .O(N__42425),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__9341 (
            .O(N__42420),
            .I(N__42417));
    InMux I__9340 (
            .O(N__42417),
            .I(N__42414));
    LocalMux I__9339 (
            .O(N__42414),
            .I(N__42411));
    Span4Mux_h I__9338 (
            .O(N__42411),
            .I(N__42408));
    Span4Mux_h I__9337 (
            .O(N__42408),
            .I(N__42405));
    Odrv4 I__9336 (
            .O(N__42405),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    CascadeMux I__9335 (
            .O(N__42402),
            .I(N__42399));
    InMux I__9334 (
            .O(N__42399),
            .I(N__42396));
    LocalMux I__9333 (
            .O(N__42396),
            .I(N__42393));
    Span4Mux_h I__9332 (
            .O(N__42393),
            .I(N__42390));
    Odrv4 I__9331 (
            .O(N__42390),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    InMux I__9330 (
            .O(N__42387),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    CascadeMux I__9329 (
            .O(N__42384),
            .I(N__42381));
    InMux I__9328 (
            .O(N__42381),
            .I(N__42378));
    LocalMux I__9327 (
            .O(N__42378),
            .I(N__42375));
    Sp12to4 I__9326 (
            .O(N__42375),
            .I(N__42370));
    InMux I__9325 (
            .O(N__42374),
            .I(N__42366));
    InMux I__9324 (
            .O(N__42373),
            .I(N__42363));
    Span12Mux_h I__9323 (
            .O(N__42370),
            .I(N__42360));
    InMux I__9322 (
            .O(N__42369),
            .I(N__42357));
    LocalMux I__9321 (
            .O(N__42366),
            .I(N__42354));
    LocalMux I__9320 (
            .O(N__42363),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv12 I__9319 (
            .O(N__42360),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__9318 (
            .O(N__42357),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__9317 (
            .O(N__42354),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    CascadeMux I__9316 (
            .O(N__42345),
            .I(N__42342));
    InMux I__9315 (
            .O(N__42342),
            .I(N__42339));
    LocalMux I__9314 (
            .O(N__42339),
            .I(N__42336));
    Span4Mux_h I__9313 (
            .O(N__42336),
            .I(N__42333));
    Span4Mux_h I__9312 (
            .O(N__42333),
            .I(N__42330));
    Odrv4 I__9311 (
            .O(N__42330),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__9310 (
            .O(N__42327),
            .I(N__42324));
    LocalMux I__9309 (
            .O(N__42324),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__9308 (
            .O(N__42321),
            .I(bfn_17_21_0_));
    CascadeMux I__9307 (
            .O(N__42318),
            .I(N__42315));
    InMux I__9306 (
            .O(N__42315),
            .I(N__42312));
    LocalMux I__9305 (
            .O(N__42312),
            .I(N__42309));
    Span4Mux_h I__9304 (
            .O(N__42309),
            .I(N__42305));
    InMux I__9303 (
            .O(N__42308),
            .I(N__42302));
    Span4Mux_v I__9302 (
            .O(N__42305),
            .I(N__42296));
    LocalMux I__9301 (
            .O(N__42302),
            .I(N__42296));
    CascadeMux I__9300 (
            .O(N__42301),
            .I(N__42293));
    Span4Mux_h I__9299 (
            .O(N__42296),
            .I(N__42289));
    InMux I__9298 (
            .O(N__42293),
            .I(N__42286));
    InMux I__9297 (
            .O(N__42292),
            .I(N__42283));
    Span4Mux_h I__9296 (
            .O(N__42289),
            .I(N__42280));
    LocalMux I__9295 (
            .O(N__42286),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    LocalMux I__9294 (
            .O(N__42283),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__9293 (
            .O(N__42280),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__9292 (
            .O(N__42273),
            .I(N__42270));
    InMux I__9291 (
            .O(N__42270),
            .I(N__42267));
    LocalMux I__9290 (
            .O(N__42267),
            .I(N__42264));
    Span4Mux_h I__9289 (
            .O(N__42264),
            .I(N__42261));
    Span4Mux_h I__9288 (
            .O(N__42261),
            .I(N__42258));
    Span4Mux_s0_h I__9287 (
            .O(N__42258),
            .I(N__42255));
    Odrv4 I__9286 (
            .O(N__42255),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__9285 (
            .O(N__42252),
            .I(N__42249));
    LocalMux I__9284 (
            .O(N__42249),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    InMux I__9283 (
            .O(N__42246),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__9282 (
            .O(N__42243),
            .I(N__42240));
    InMux I__9281 (
            .O(N__42240),
            .I(N__42237));
    LocalMux I__9280 (
            .O(N__42237),
            .I(N__42233));
    InMux I__9279 (
            .O(N__42236),
            .I(N__42230));
    Span4Mux_v I__9278 (
            .O(N__42233),
            .I(N__42227));
    LocalMux I__9277 (
            .O(N__42230),
            .I(N__42223));
    Sp12to4 I__9276 (
            .O(N__42227),
            .I(N__42219));
    InMux I__9275 (
            .O(N__42226),
            .I(N__42216));
    Span12Mux_v I__9274 (
            .O(N__42223),
            .I(N__42213));
    InMux I__9273 (
            .O(N__42222),
            .I(N__42210));
    Span12Mux_h I__9272 (
            .O(N__42219),
            .I(N__42207));
    LocalMux I__9271 (
            .O(N__42216),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv12 I__9270 (
            .O(N__42213),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__9269 (
            .O(N__42210),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv12 I__9268 (
            .O(N__42207),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__9267 (
            .O(N__42198),
            .I(N__42195));
    LocalMux I__9266 (
            .O(N__42195),
            .I(N__42192));
    Span4Mux_v I__9265 (
            .O(N__42192),
            .I(N__42188));
    InMux I__9264 (
            .O(N__42191),
            .I(N__42184));
    Span4Mux_v I__9263 (
            .O(N__42188),
            .I(N__42181));
    InMux I__9262 (
            .O(N__42187),
            .I(N__42178));
    LocalMux I__9261 (
            .O(N__42184),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    Odrv4 I__9260 (
            .O(N__42181),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    LocalMux I__9259 (
            .O(N__42178),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__9258 (
            .O(N__42171),
            .I(N__42165));
    InMux I__9257 (
            .O(N__42170),
            .I(N__42165));
    LocalMux I__9256 (
            .O(N__42165),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ));
    CascadeMux I__9255 (
            .O(N__42162),
            .I(N__42159));
    InMux I__9254 (
            .O(N__42159),
            .I(N__42156));
    LocalMux I__9253 (
            .O(N__42156),
            .I(N__42153));
    Span4Mux_h I__9252 (
            .O(N__42153),
            .I(N__42149));
    InMux I__9251 (
            .O(N__42152),
            .I(N__42146));
    Sp12to4 I__9250 (
            .O(N__42149),
            .I(N__42143));
    LocalMux I__9249 (
            .O(N__42146),
            .I(N__42140));
    Span12Mux_v I__9248 (
            .O(N__42143),
            .I(N__42137));
    Odrv4 I__9247 (
            .O(N__42140),
            .I(\phase_controller_inst2.stoper_hc.N_47 ));
    Odrv12 I__9246 (
            .O(N__42137),
            .I(\phase_controller_inst2.stoper_hc.N_47 ));
    InMux I__9245 (
            .O(N__42132),
            .I(N__42129));
    LocalMux I__9244 (
            .O(N__42129),
            .I(N__42125));
    InMux I__9243 (
            .O(N__42128),
            .I(N__42122));
    Span4Mux_v I__9242 (
            .O(N__42125),
            .I(N__42119));
    LocalMux I__9241 (
            .O(N__42122),
            .I(N__42116));
    Sp12to4 I__9240 (
            .O(N__42119),
            .I(N__42112));
    Span12Mux_v I__9239 (
            .O(N__42116),
            .I(N__42109));
    InMux I__9238 (
            .O(N__42115),
            .I(N__42106));
    Span12Mux_h I__9237 (
            .O(N__42112),
            .I(N__42103));
    Span12Mux_v I__9236 (
            .O(N__42109),
            .I(N__42098));
    LocalMux I__9235 (
            .O(N__42106),
            .I(N__42098));
    Span12Mux_v I__9234 (
            .O(N__42103),
            .I(N__42093));
    Span12Mux_h I__9233 (
            .O(N__42098),
            .I(N__42093));
    Odrv12 I__9232 (
            .O(N__42093),
            .I(il_max_comp2_c));
    InMux I__9231 (
            .O(N__42090),
            .I(N__42084));
    InMux I__9230 (
            .O(N__42089),
            .I(N__42084));
    LocalMux I__9229 (
            .O(N__42084),
            .I(N__42080));
    InMux I__9228 (
            .O(N__42083),
            .I(N__42077));
    Span4Mux_v I__9227 (
            .O(N__42080),
            .I(N__42074));
    LocalMux I__9226 (
            .O(N__42077),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    Odrv4 I__9225 (
            .O(N__42074),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__9224 (
            .O(N__42069),
            .I(N__42065));
    CascadeMux I__9223 (
            .O(N__42068),
            .I(N__42061));
    LocalMux I__9222 (
            .O(N__42065),
            .I(N__42058));
    InMux I__9221 (
            .O(N__42064),
            .I(N__42053));
    InMux I__9220 (
            .O(N__42061),
            .I(N__42053));
    Span4Mux_v I__9219 (
            .O(N__42058),
            .I(N__42050));
    LocalMux I__9218 (
            .O(N__42053),
            .I(N__42046));
    Span4Mux_v I__9217 (
            .O(N__42050),
            .I(N__42042));
    InMux I__9216 (
            .O(N__42049),
            .I(N__42039));
    Span4Mux_v I__9215 (
            .O(N__42046),
            .I(N__42036));
    InMux I__9214 (
            .O(N__42045),
            .I(N__42033));
    Span4Mux_v I__9213 (
            .O(N__42042),
            .I(N__42030));
    LocalMux I__9212 (
            .O(N__42039),
            .I(N__42025));
    Span4Mux_h I__9211 (
            .O(N__42036),
            .I(N__42025));
    LocalMux I__9210 (
            .O(N__42033),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__9209 (
            .O(N__42030),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__9208 (
            .O(N__42025),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__9207 (
            .O(N__42018),
            .I(N__42014));
    InMux I__9206 (
            .O(N__42017),
            .I(N__42011));
    LocalMux I__9205 (
            .O(N__42014),
            .I(N__42006));
    LocalMux I__9204 (
            .O(N__42011),
            .I(N__42006));
    Span4Mux_v I__9203 (
            .O(N__42006),
            .I(N__42000));
    InMux I__9202 (
            .O(N__42005),
            .I(N__41993));
    InMux I__9201 (
            .O(N__42004),
            .I(N__41993));
    InMux I__9200 (
            .O(N__42003),
            .I(N__41993));
    Odrv4 I__9199 (
            .O(N__42000),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__9198 (
            .O(N__41993),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__9197 (
            .O(N__41988),
            .I(N__41985));
    LocalMux I__9196 (
            .O(N__41985),
            .I(N__41981));
    InMux I__9195 (
            .O(N__41984),
            .I(N__41978));
    Span4Mux_h I__9194 (
            .O(N__41981),
            .I(N__41975));
    LocalMux I__9193 (
            .O(N__41978),
            .I(N__41972));
    Span4Mux_v I__9192 (
            .O(N__41975),
            .I(N__41969));
    Span4Mux_h I__9191 (
            .O(N__41972),
            .I(N__41964));
    Span4Mux_v I__9190 (
            .O(N__41969),
            .I(N__41964));
    Odrv4 I__9189 (
            .O(N__41964),
            .I(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971Z0Z_30 ));
    InMux I__9188 (
            .O(N__41961),
            .I(N__41958));
    LocalMux I__9187 (
            .O(N__41958),
            .I(N__41955));
    Span4Mux_v I__9186 (
            .O(N__41955),
            .I(N__41952));
    Span4Mux_h I__9185 (
            .O(N__41952),
            .I(N__41949));
    Odrv4 I__9184 (
            .O(N__41949),
            .I(\phase_controller_inst2.stoper_hc.mZ0Z16 ));
    CascadeMux I__9183 (
            .O(N__41946),
            .I(N__41943));
    InMux I__9182 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__9181 (
            .O(N__41940),
            .I(N__41937));
    Span4Mux_h I__9180 (
            .O(N__41937),
            .I(N__41934));
    Sp12to4 I__9179 (
            .O(N__41934),
            .I(N__41931));
    Span12Mux_v I__9178 (
            .O(N__41931),
            .I(N__41928));
    Odrv12 I__9177 (
            .O(N__41928),
            .I(\phase_controller_inst2.stoper_hc.m28_ns_1 ));
    InMux I__9176 (
            .O(N__41925),
            .I(N__41919));
    InMux I__9175 (
            .O(N__41924),
            .I(N__41919));
    LocalMux I__9174 (
            .O(N__41919),
            .I(N__41915));
    InMux I__9173 (
            .O(N__41918),
            .I(N__41912));
    Span4Mux_h I__9172 (
            .O(N__41915),
            .I(N__41909));
    LocalMux I__9171 (
            .O(N__41912),
            .I(N__41905));
    Span4Mux_v I__9170 (
            .O(N__41909),
            .I(N__41902));
    InMux I__9169 (
            .O(N__41908),
            .I(N__41899));
    Span12Mux_h I__9168 (
            .O(N__41905),
            .I(N__41896));
    Span4Mux_v I__9167 (
            .O(N__41902),
            .I(N__41893));
    LocalMux I__9166 (
            .O(N__41899),
            .I(N__41888));
    Span12Mux_v I__9165 (
            .O(N__41896),
            .I(N__41885));
    Span4Mux_v I__9164 (
            .O(N__41893),
            .I(N__41882));
    InMux I__9163 (
            .O(N__41892),
            .I(N__41879));
    InMux I__9162 (
            .O(N__41891),
            .I(N__41876));
    Span4Mux_h I__9161 (
            .O(N__41888),
            .I(N__41873));
    Odrv12 I__9160 (
            .O(N__41885),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    Odrv4 I__9159 (
            .O(N__41882),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    LocalMux I__9158 (
            .O(N__41879),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    LocalMux I__9157 (
            .O(N__41876),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    Odrv4 I__9156 (
            .O(N__41873),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    InMux I__9155 (
            .O(N__41862),
            .I(N__41859));
    LocalMux I__9154 (
            .O(N__41859),
            .I(N__41853));
    CascadeMux I__9153 (
            .O(N__41858),
            .I(N__41850));
    CascadeMux I__9152 (
            .O(N__41857),
            .I(N__41847));
    CascadeMux I__9151 (
            .O(N__41856),
            .I(N__41844));
    Span4Mux_h I__9150 (
            .O(N__41853),
            .I(N__41840));
    InMux I__9149 (
            .O(N__41850),
            .I(N__41837));
    InMux I__9148 (
            .O(N__41847),
            .I(N__41832));
    InMux I__9147 (
            .O(N__41844),
            .I(N__41832));
    InMux I__9146 (
            .O(N__41843),
            .I(N__41829));
    Sp12to4 I__9145 (
            .O(N__41840),
            .I(N__41820));
    LocalMux I__9144 (
            .O(N__41837),
            .I(N__41820));
    LocalMux I__9143 (
            .O(N__41832),
            .I(N__41820));
    LocalMux I__9142 (
            .O(N__41829),
            .I(N__41820));
    Span12Mux_s6_v I__9141 (
            .O(N__41820),
            .I(N__41816));
    InMux I__9140 (
            .O(N__41819),
            .I(N__41813));
    Span12Mux_v I__9139 (
            .O(N__41816),
            .I(N__41810));
    LocalMux I__9138 (
            .O(N__41813),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__9137 (
            .O(N__41810),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    CascadeMux I__9136 (
            .O(N__41805),
            .I(N__41802));
    InMux I__9135 (
            .O(N__41802),
            .I(N__41799));
    LocalMux I__9134 (
            .O(N__41799),
            .I(N__41796));
    Span4Mux_v I__9133 (
            .O(N__41796),
            .I(N__41791));
    InMux I__9132 (
            .O(N__41795),
            .I(N__41787));
    CascadeMux I__9131 (
            .O(N__41794),
            .I(N__41784));
    Span4Mux_v I__9130 (
            .O(N__41791),
            .I(N__41781));
    InMux I__9129 (
            .O(N__41790),
            .I(N__41778));
    LocalMux I__9128 (
            .O(N__41787),
            .I(N__41774));
    InMux I__9127 (
            .O(N__41784),
            .I(N__41771));
    Span4Mux_h I__9126 (
            .O(N__41781),
            .I(N__41768));
    LocalMux I__9125 (
            .O(N__41778),
            .I(N__41765));
    InMux I__9124 (
            .O(N__41777),
            .I(N__41762));
    Span12Mux_h I__9123 (
            .O(N__41774),
            .I(N__41759));
    LocalMux I__9122 (
            .O(N__41771),
            .I(N__41756));
    Span4Mux_h I__9121 (
            .O(N__41768),
            .I(N__41751));
    Span4Mux_v I__9120 (
            .O(N__41765),
            .I(N__41751));
    LocalMux I__9119 (
            .O(N__41762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv12 I__9118 (
            .O(N__41759),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__9117 (
            .O(N__41756),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    Odrv4 I__9116 (
            .O(N__41751),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    CascadeMux I__9115 (
            .O(N__41742),
            .I(N__41739));
    InMux I__9114 (
            .O(N__41739),
            .I(N__41735));
    CascadeMux I__9113 (
            .O(N__41738),
            .I(N__41732));
    LocalMux I__9112 (
            .O(N__41735),
            .I(N__41729));
    InMux I__9111 (
            .O(N__41732),
            .I(N__41726));
    Span4Mux_v I__9110 (
            .O(N__41729),
            .I(N__41723));
    LocalMux I__9109 (
            .O(N__41726),
            .I(N__41720));
    Span4Mux_h I__9108 (
            .O(N__41723),
            .I(N__41717));
    Span4Mux_h I__9107 (
            .O(N__41720),
            .I(N__41714));
    Span4Mux_h I__9106 (
            .O(N__41717),
            .I(N__41711));
    Span4Mux_h I__9105 (
            .O(N__41714),
            .I(N__41708));
    Odrv4 I__9104 (
            .O(N__41711),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    Odrv4 I__9103 (
            .O(N__41708),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__9102 (
            .O(N__41703),
            .I(N__41700));
    InMux I__9101 (
            .O(N__41700),
            .I(N__41697));
    LocalMux I__9100 (
            .O(N__41697),
            .I(N__41694));
    Span4Mux_v I__9099 (
            .O(N__41694),
            .I(N__41689));
    InMux I__9098 (
            .O(N__41693),
            .I(N__41686));
    InMux I__9097 (
            .O(N__41692),
            .I(N__41683));
    Sp12to4 I__9096 (
            .O(N__41689),
            .I(N__41680));
    LocalMux I__9095 (
            .O(N__41686),
            .I(N__41677));
    LocalMux I__9094 (
            .O(N__41683),
            .I(N__41672));
    Span12Mux_h I__9093 (
            .O(N__41680),
            .I(N__41672));
    Span4Mux_h I__9092 (
            .O(N__41677),
            .I(N__41669));
    Odrv12 I__9091 (
            .O(N__41672),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    Odrv4 I__9090 (
            .O(N__41669),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    CascadeMux I__9089 (
            .O(N__41664),
            .I(N__41661));
    InMux I__9088 (
            .O(N__41661),
            .I(N__41658));
    LocalMux I__9087 (
            .O(N__41658),
            .I(N__41655));
    Span4Mux_h I__9086 (
            .O(N__41655),
            .I(N__41652));
    Span4Mux_h I__9085 (
            .O(N__41652),
            .I(N__41649));
    Odrv4 I__9084 (
            .O(N__41649),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__9083 (
            .O(N__41646),
            .I(N__41643));
    LocalMux I__9082 (
            .O(N__41643),
            .I(N__41640));
    Span4Mux_v I__9081 (
            .O(N__41640),
            .I(N__41637));
    Odrv4 I__9080 (
            .O(N__41637),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ));
    InMux I__9079 (
            .O(N__41634),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__9078 (
            .O(N__41631),
            .I(N__41628));
    InMux I__9077 (
            .O(N__41628),
            .I(N__41624));
    InMux I__9076 (
            .O(N__41627),
            .I(N__41621));
    LocalMux I__9075 (
            .O(N__41624),
            .I(N__41618));
    LocalMux I__9074 (
            .O(N__41621),
            .I(N__41615));
    Span4Mux_h I__9073 (
            .O(N__41618),
            .I(N__41610));
    Span4Mux_h I__9072 (
            .O(N__41615),
            .I(N__41607));
    InMux I__9071 (
            .O(N__41614),
            .I(N__41604));
    InMux I__9070 (
            .O(N__41613),
            .I(N__41601));
    Span4Mux_v I__9069 (
            .O(N__41610),
            .I(N__41596));
    Span4Mux_h I__9068 (
            .O(N__41607),
            .I(N__41596));
    LocalMux I__9067 (
            .O(N__41604),
            .I(N__41591));
    LocalMux I__9066 (
            .O(N__41601),
            .I(N__41591));
    Odrv4 I__9065 (
            .O(N__41596),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    Odrv12 I__9064 (
            .O(N__41591),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__9063 (
            .O(N__41586),
            .I(N__41583));
    InMux I__9062 (
            .O(N__41583),
            .I(N__41580));
    LocalMux I__9061 (
            .O(N__41580),
            .I(N__41577));
    Span4Mux_h I__9060 (
            .O(N__41577),
            .I(N__41574));
    Span4Mux_h I__9059 (
            .O(N__41574),
            .I(N__41571));
    Odrv4 I__9058 (
            .O(N__41571),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__9057 (
            .O(N__41568),
            .I(N__41565));
    LocalMux I__9056 (
            .O(N__41565),
            .I(N__41562));
    Span12Mux_s11_h I__9055 (
            .O(N__41562),
            .I(N__41559));
    Odrv12 I__9054 (
            .O(N__41559),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ));
    InMux I__9053 (
            .O(N__41556),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__9052 (
            .O(N__41553),
            .I(N__41549));
    InMux I__9051 (
            .O(N__41552),
            .I(N__41544));
    InMux I__9050 (
            .O(N__41549),
            .I(N__41544));
    LocalMux I__9049 (
            .O(N__41544),
            .I(N__41541));
    Span4Mux_v I__9048 (
            .O(N__41541),
            .I(N__41537));
    InMux I__9047 (
            .O(N__41540),
            .I(N__41534));
    Span4Mux_h I__9046 (
            .O(N__41537),
            .I(N__41531));
    LocalMux I__9045 (
            .O(N__41534),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__9044 (
            .O(N__41531),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ));
    InMux I__9043 (
            .O(N__41526),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__9042 (
            .O(N__41523),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__9041 (
            .O(N__41520),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ));
    CascadeMux I__9040 (
            .O(N__41517),
            .I(N__41512));
    InMux I__9039 (
            .O(N__41516),
            .I(N__41509));
    InMux I__9038 (
            .O(N__41515),
            .I(N__41504));
    InMux I__9037 (
            .O(N__41512),
            .I(N__41504));
    LocalMux I__9036 (
            .O(N__41509),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    LocalMux I__9035 (
            .O(N__41504),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__9034 (
            .O(N__41499),
            .I(N__41494));
    InMux I__9033 (
            .O(N__41498),
            .I(N__41489));
    InMux I__9032 (
            .O(N__41497),
            .I(N__41489));
    LocalMux I__9031 (
            .O(N__41494),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    LocalMux I__9030 (
            .O(N__41489),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ));
    InMux I__9029 (
            .O(N__41484),
            .I(N__41480));
    InMux I__9028 (
            .O(N__41483),
            .I(N__41477));
    LocalMux I__9027 (
            .O(N__41480),
            .I(N__41473));
    LocalMux I__9026 (
            .O(N__41477),
            .I(N__41470));
    InMux I__9025 (
            .O(N__41476),
            .I(N__41467));
    Span4Mux_v I__9024 (
            .O(N__41473),
            .I(N__41464));
    Span4Mux_h I__9023 (
            .O(N__41470),
            .I(N__41461));
    LocalMux I__9022 (
            .O(N__41467),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv4 I__9021 (
            .O(N__41464),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv4 I__9020 (
            .O(N__41461),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__9019 (
            .O(N__41454),
            .I(N__41448));
    InMux I__9018 (
            .O(N__41453),
            .I(N__41448));
    LocalMux I__9017 (
            .O(N__41448),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ));
    CascadeMux I__9016 (
            .O(N__41445),
            .I(N__41441));
    InMux I__9015 (
            .O(N__41444),
            .I(N__41437));
    InMux I__9014 (
            .O(N__41441),
            .I(N__41432));
    InMux I__9013 (
            .O(N__41440),
            .I(N__41432));
    LocalMux I__9012 (
            .O(N__41437),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__9011 (
            .O(N__41432),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__9010 (
            .O(N__41427),
            .I(N__41424));
    InMux I__9009 (
            .O(N__41424),
            .I(N__41418));
    InMux I__9008 (
            .O(N__41423),
            .I(N__41418));
    LocalMux I__9007 (
            .O(N__41418),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ));
    InMux I__9006 (
            .O(N__41415),
            .I(N__41410));
    InMux I__9005 (
            .O(N__41414),
            .I(N__41405));
    InMux I__9004 (
            .O(N__41413),
            .I(N__41405));
    LocalMux I__9003 (
            .O(N__41410),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__9002 (
            .O(N__41405),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ));
    CascadeMux I__9001 (
            .O(N__41400),
            .I(N__41397));
    InMux I__9000 (
            .O(N__41397),
            .I(N__41391));
    InMux I__8999 (
            .O(N__41396),
            .I(N__41391));
    LocalMux I__8998 (
            .O(N__41391),
            .I(N__41387));
    InMux I__8997 (
            .O(N__41390),
            .I(N__41384));
    Span4Mux_h I__8996 (
            .O(N__41387),
            .I(N__41381));
    LocalMux I__8995 (
            .O(N__41384),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__8994 (
            .O(N__41381),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__8993 (
            .O(N__41376),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__8992 (
            .O(N__41373),
            .I(N__41366));
    InMux I__8991 (
            .O(N__41372),
            .I(N__41366));
    InMux I__8990 (
            .O(N__41371),
            .I(N__41363));
    LocalMux I__8989 (
            .O(N__41366),
            .I(N__41360));
    LocalMux I__8988 (
            .O(N__41363),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__8987 (
            .O(N__41360),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__8986 (
            .O(N__41355),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__8985 (
            .O(N__41352),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__8984 (
            .O(N__41349),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__8983 (
            .O(N__41346),
            .I(N__41339));
    InMux I__8982 (
            .O(N__41345),
            .I(N__41339));
    InMux I__8981 (
            .O(N__41344),
            .I(N__41336));
    LocalMux I__8980 (
            .O(N__41339),
            .I(N__41333));
    LocalMux I__8979 (
            .O(N__41336),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__8978 (
            .O(N__41333),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__8977 (
            .O(N__41328),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__8976 (
            .O(N__41325),
            .I(N__41320));
    InMux I__8975 (
            .O(N__41324),
            .I(N__41315));
    InMux I__8974 (
            .O(N__41323),
            .I(N__41315));
    LocalMux I__8973 (
            .O(N__41320),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__8972 (
            .O(N__41315),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__8971 (
            .O(N__41310),
            .I(bfn_17_17_0_));
    InMux I__8970 (
            .O(N__41307),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__8969 (
            .O(N__41304),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__8968 (
            .O(N__41301),
            .I(N__41295));
    InMux I__8967 (
            .O(N__41300),
            .I(N__41295));
    LocalMux I__8966 (
            .O(N__41295),
            .I(N__41292));
    Span4Mux_v I__8965 (
            .O(N__41292),
            .I(N__41288));
    InMux I__8964 (
            .O(N__41291),
            .I(N__41285));
    Span4Mux_h I__8963 (
            .O(N__41288),
            .I(N__41282));
    LocalMux I__8962 (
            .O(N__41285),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__8961 (
            .O(N__41282),
            .I(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ));
    InMux I__8960 (
            .O(N__41277),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__8959 (
            .O(N__41274),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__8958 (
            .O(N__41271),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__8957 (
            .O(N__41268),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__8956 (
            .O(N__41265),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__8955 (
            .O(N__41262),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__8954 (
            .O(N__41259),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__8953 (
            .O(N__41256),
            .I(bfn_17_16_0_));
    InMux I__8952 (
            .O(N__41253),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__8951 (
            .O(N__41250),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__8950 (
            .O(N__41247),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__8949 (
            .O(N__41244),
            .I(N__41240));
    CascadeMux I__8948 (
            .O(N__41243),
            .I(N__41237));
    InMux I__8947 (
            .O(N__41240),
            .I(N__41232));
    InMux I__8946 (
            .O(N__41237),
            .I(N__41232));
    LocalMux I__8945 (
            .O(N__41232),
            .I(\phase_controller_inst2.stoper_hc.N_265_i ));
    InMux I__8944 (
            .O(N__41229),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__8943 (
            .O(N__41226),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__8942 (
            .O(N__41223),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__8941 (
            .O(N__41220),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__8940 (
            .O(N__41217),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__8939 (
            .O(N__41214),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__8938 (
            .O(N__41211),
            .I(bfn_17_15_0_));
    InMux I__8937 (
            .O(N__41208),
            .I(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__8936 (
            .O(N__41205),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    InMux I__8935 (
            .O(N__41202),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    InMux I__8934 (
            .O(N__41199),
            .I(bfn_17_13_0_));
    InMux I__8933 (
            .O(N__41196),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    InMux I__8932 (
            .O(N__41193),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    InMux I__8931 (
            .O(N__41190),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__8930 (
            .O(N__41187),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__8929 (
            .O(N__41184),
            .I(N__41168));
    InMux I__8928 (
            .O(N__41183),
            .I(N__41168));
    InMux I__8927 (
            .O(N__41182),
            .I(N__41168));
    InMux I__8926 (
            .O(N__41181),
            .I(N__41168));
    InMux I__8925 (
            .O(N__41180),
            .I(N__41143));
    InMux I__8924 (
            .O(N__41179),
            .I(N__41143));
    InMux I__8923 (
            .O(N__41178),
            .I(N__41143));
    InMux I__8922 (
            .O(N__41177),
            .I(N__41143));
    LocalMux I__8921 (
            .O(N__41168),
            .I(N__41134));
    InMux I__8920 (
            .O(N__41167),
            .I(N__41125));
    InMux I__8919 (
            .O(N__41166),
            .I(N__41125));
    InMux I__8918 (
            .O(N__41165),
            .I(N__41125));
    InMux I__8917 (
            .O(N__41164),
            .I(N__41125));
    InMux I__8916 (
            .O(N__41163),
            .I(N__41116));
    InMux I__8915 (
            .O(N__41162),
            .I(N__41116));
    InMux I__8914 (
            .O(N__41161),
            .I(N__41116));
    InMux I__8913 (
            .O(N__41160),
            .I(N__41116));
    InMux I__8912 (
            .O(N__41159),
            .I(N__41107));
    InMux I__8911 (
            .O(N__41158),
            .I(N__41107));
    InMux I__8910 (
            .O(N__41157),
            .I(N__41107));
    InMux I__8909 (
            .O(N__41156),
            .I(N__41107));
    InMux I__8908 (
            .O(N__41155),
            .I(N__41098));
    InMux I__8907 (
            .O(N__41154),
            .I(N__41098));
    InMux I__8906 (
            .O(N__41153),
            .I(N__41098));
    InMux I__8905 (
            .O(N__41152),
            .I(N__41098));
    LocalMux I__8904 (
            .O(N__41143),
            .I(N__41095));
    InMux I__8903 (
            .O(N__41142),
            .I(N__41090));
    InMux I__8902 (
            .O(N__41141),
            .I(N__41090));
    InMux I__8901 (
            .O(N__41140),
            .I(N__41081));
    InMux I__8900 (
            .O(N__41139),
            .I(N__41081));
    InMux I__8899 (
            .O(N__41138),
            .I(N__41081));
    InMux I__8898 (
            .O(N__41137),
            .I(N__41081));
    Span4Mux_v I__8897 (
            .O(N__41134),
            .I(N__41078));
    LocalMux I__8896 (
            .O(N__41125),
            .I(N__41069));
    LocalMux I__8895 (
            .O(N__41116),
            .I(N__41069));
    LocalMux I__8894 (
            .O(N__41107),
            .I(N__41069));
    LocalMux I__8893 (
            .O(N__41098),
            .I(N__41069));
    Span4Mux_h I__8892 (
            .O(N__41095),
            .I(N__41066));
    LocalMux I__8891 (
            .O(N__41090),
            .I(N__41057));
    LocalMux I__8890 (
            .O(N__41081),
            .I(N__41057));
    Span4Mux_h I__8889 (
            .O(N__41078),
            .I(N__41057));
    Span4Mux_v I__8888 (
            .O(N__41069),
            .I(N__41057));
    Odrv4 I__8887 (
            .O(N__41066),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__8886 (
            .O(N__41057),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    InMux I__8885 (
            .O(N__41052),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    CEMux I__8884 (
            .O(N__41049),
            .I(N__41045));
    CEMux I__8883 (
            .O(N__41048),
            .I(N__41042));
    LocalMux I__8882 (
            .O(N__41045),
            .I(N__41037));
    LocalMux I__8881 (
            .O(N__41042),
            .I(N__41034));
    CEMux I__8880 (
            .O(N__41041),
            .I(N__41031));
    CEMux I__8879 (
            .O(N__41040),
            .I(N__41028));
    Span4Mux_v I__8878 (
            .O(N__41037),
            .I(N__41025));
    Span4Mux_h I__8877 (
            .O(N__41034),
            .I(N__41022));
    LocalMux I__8876 (
            .O(N__41031),
            .I(N__41019));
    LocalMux I__8875 (
            .O(N__41028),
            .I(N__41016));
    Span4Mux_v I__8874 (
            .O(N__41025),
            .I(N__41013));
    Span4Mux_v I__8873 (
            .O(N__41022),
            .I(N__41010));
    Span4Mux_h I__8872 (
            .O(N__41019),
            .I(N__41007));
    Span4Mux_h I__8871 (
            .O(N__41016),
            .I(N__41004));
    Odrv4 I__8870 (
            .O(N__41013),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    Odrv4 I__8869 (
            .O(N__41010),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    Odrv4 I__8868 (
            .O(N__41007),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    Odrv4 I__8867 (
            .O(N__41004),
            .I(\delay_measurement_inst.delay_hc_timer.N_342_i ));
    InMux I__8866 (
            .O(N__40995),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__8865 (
            .O(N__40992),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    InMux I__8864 (
            .O(N__40989),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    InMux I__8863 (
            .O(N__40986),
            .I(bfn_17_12_0_));
    InMux I__8862 (
            .O(N__40983),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__8861 (
            .O(N__40980),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__8860 (
            .O(N__40977),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    InMux I__8859 (
            .O(N__40974),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    InMux I__8858 (
            .O(N__40971),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__8857 (
            .O(N__40968),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    InMux I__8856 (
            .O(N__40965),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__8855 (
            .O(N__40962),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    InMux I__8854 (
            .O(N__40959),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__8853 (
            .O(N__40956),
            .I(bfn_17_11_0_));
    InMux I__8852 (
            .O(N__40953),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    InMux I__8851 (
            .O(N__40950),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__8850 (
            .O(N__40947),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    InMux I__8849 (
            .O(N__40944),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    InMux I__8848 (
            .O(N__40941),
            .I(N__40935));
    InMux I__8847 (
            .O(N__40940),
            .I(N__40935));
    LocalMux I__8846 (
            .O(N__40935),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ));
    InMux I__8845 (
            .O(N__40932),
            .I(N__40929));
    LocalMux I__8844 (
            .O(N__40929),
            .I(N__40925));
    InMux I__8843 (
            .O(N__40928),
            .I(N__40921));
    Span4Mux_v I__8842 (
            .O(N__40925),
            .I(N__40918));
    InMux I__8841 (
            .O(N__40924),
            .I(N__40915));
    LocalMux I__8840 (
            .O(N__40921),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    Odrv4 I__8839 (
            .O(N__40918),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    LocalMux I__8838 (
            .O(N__40915),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    CascadeMux I__8837 (
            .O(N__40908),
            .I(N__40905));
    InMux I__8836 (
            .O(N__40905),
            .I(N__40902));
    LocalMux I__8835 (
            .O(N__40902),
            .I(N__40899));
    Odrv4 I__8834 (
            .O(N__40899),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt22 ));
    InMux I__8833 (
            .O(N__40896),
            .I(N__40890));
    InMux I__8832 (
            .O(N__40895),
            .I(N__40890));
    LocalMux I__8831 (
            .O(N__40890),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ));
    InMux I__8830 (
            .O(N__40887),
            .I(N__40881));
    InMux I__8829 (
            .O(N__40886),
            .I(N__40881));
    LocalMux I__8828 (
            .O(N__40881),
            .I(N__40877));
    InMux I__8827 (
            .O(N__40880),
            .I(N__40874));
    Span4Mux_h I__8826 (
            .O(N__40877),
            .I(N__40871));
    LocalMux I__8825 (
            .O(N__40874),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    Odrv4 I__8824 (
            .O(N__40871),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ));
    InMux I__8823 (
            .O(N__40866),
            .I(N__40860));
    InMux I__8822 (
            .O(N__40865),
            .I(N__40860));
    LocalMux I__8821 (
            .O(N__40860),
            .I(N__40856));
    InMux I__8820 (
            .O(N__40859),
            .I(N__40853));
    Span4Mux_h I__8819 (
            .O(N__40856),
            .I(N__40850));
    LocalMux I__8818 (
            .O(N__40853),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    Odrv4 I__8817 (
            .O(N__40850),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ));
    InMux I__8816 (
            .O(N__40845),
            .I(N__40842));
    LocalMux I__8815 (
            .O(N__40842),
            .I(N__40839));
    Odrv4 I__8814 (
            .O(N__40839),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ));
    InMux I__8813 (
            .O(N__40836),
            .I(bfn_17_10_0_));
    InMux I__8812 (
            .O(N__40833),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    InMux I__8811 (
            .O(N__40830),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__8810 (
            .O(N__40827),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    InMux I__8809 (
            .O(N__40824),
            .I(N__40821));
    LocalMux I__8808 (
            .O(N__40821),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt16 ));
    InMux I__8807 (
            .O(N__40818),
            .I(N__40812));
    InMux I__8806 (
            .O(N__40817),
            .I(N__40812));
    LocalMux I__8805 (
            .O(N__40812),
            .I(N__40808));
    InMux I__8804 (
            .O(N__40811),
            .I(N__40805));
    Span4Mux_v I__8803 (
            .O(N__40808),
            .I(N__40802));
    LocalMux I__8802 (
            .O(N__40805),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    Odrv4 I__8801 (
            .O(N__40802),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ));
    CascadeMux I__8800 (
            .O(N__40797),
            .I(N__40792));
    CascadeMux I__8799 (
            .O(N__40796),
            .I(N__40789));
    InMux I__8798 (
            .O(N__40795),
            .I(N__40786));
    InMux I__8797 (
            .O(N__40792),
            .I(N__40783));
    InMux I__8796 (
            .O(N__40789),
            .I(N__40780));
    LocalMux I__8795 (
            .O(N__40786),
            .I(N__40773));
    LocalMux I__8794 (
            .O(N__40783),
            .I(N__40773));
    LocalMux I__8793 (
            .O(N__40780),
            .I(N__40773));
    Odrv4 I__8792 (
            .O(N__40773),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ));
    CascadeMux I__8791 (
            .O(N__40770),
            .I(N__40767));
    InMux I__8790 (
            .O(N__40767),
            .I(N__40764));
    LocalMux I__8789 (
            .O(N__40764),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ));
    InMux I__8788 (
            .O(N__40761),
            .I(N__40755));
    InMux I__8787 (
            .O(N__40760),
            .I(N__40755));
    LocalMux I__8786 (
            .O(N__40755),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ));
    InMux I__8785 (
            .O(N__40752),
            .I(N__40749));
    LocalMux I__8784 (
            .O(N__40749),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ));
    InMux I__8783 (
            .O(N__40746),
            .I(N__40743));
    LocalMux I__8782 (
            .O(N__40743),
            .I(N__40740));
    Span4Mux_v I__8781 (
            .O(N__40740),
            .I(N__40737));
    Span4Mux_v I__8780 (
            .O(N__40737),
            .I(N__40733));
    InMux I__8779 (
            .O(N__40736),
            .I(N__40730));
    Odrv4 I__8778 (
            .O(N__40733),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    LocalMux I__8777 (
            .O(N__40730),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    CascadeMux I__8776 (
            .O(N__40725),
            .I(N__40722));
    InMux I__8775 (
            .O(N__40722),
            .I(N__40719));
    LocalMux I__8774 (
            .O(N__40719),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ));
    InMux I__8773 (
            .O(N__40716),
            .I(N__40713));
    LocalMux I__8772 (
            .O(N__40713),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ));
    InMux I__8771 (
            .O(N__40710),
            .I(N__40707));
    LocalMux I__8770 (
            .O(N__40707),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ));
    CascadeMux I__8769 (
            .O(N__40704),
            .I(N__40701));
    InMux I__8768 (
            .O(N__40701),
            .I(N__40698));
    LocalMux I__8767 (
            .O(N__40698),
            .I(N__40695));
    Odrv4 I__8766 (
            .O(N__40695),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt26 ));
    CascadeMux I__8765 (
            .O(N__40692),
            .I(N__40687));
    InMux I__8764 (
            .O(N__40691),
            .I(N__40684));
    InMux I__8763 (
            .O(N__40690),
            .I(N__40679));
    InMux I__8762 (
            .O(N__40687),
            .I(N__40679));
    LocalMux I__8761 (
            .O(N__40684),
            .I(N__40674));
    LocalMux I__8760 (
            .O(N__40679),
            .I(N__40674));
    Odrv4 I__8759 (
            .O(N__40674),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ));
    CascadeMux I__8758 (
            .O(N__40671),
            .I(N__40666));
    InMux I__8757 (
            .O(N__40670),
            .I(N__40663));
    InMux I__8756 (
            .O(N__40669),
            .I(N__40658));
    InMux I__8755 (
            .O(N__40666),
            .I(N__40658));
    LocalMux I__8754 (
            .O(N__40663),
            .I(N__40653));
    LocalMux I__8753 (
            .O(N__40658),
            .I(N__40653));
    Odrv4 I__8752 (
            .O(N__40653),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ));
    InMux I__8751 (
            .O(N__40650),
            .I(N__40647));
    LocalMux I__8750 (
            .O(N__40647),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ));
    CascadeMux I__8749 (
            .O(N__40644),
            .I(N__40639));
    CascadeMux I__8748 (
            .O(N__40643),
            .I(N__40636));
    InMux I__8747 (
            .O(N__40642),
            .I(N__40632));
    InMux I__8746 (
            .O(N__40639),
            .I(N__40628));
    InMux I__8745 (
            .O(N__40636),
            .I(N__40625));
    InMux I__8744 (
            .O(N__40635),
            .I(N__40622));
    LocalMux I__8743 (
            .O(N__40632),
            .I(N__40619));
    InMux I__8742 (
            .O(N__40631),
            .I(N__40616));
    LocalMux I__8741 (
            .O(N__40628),
            .I(N__40610));
    LocalMux I__8740 (
            .O(N__40625),
            .I(N__40610));
    LocalMux I__8739 (
            .O(N__40622),
            .I(N__40603));
    Span4Mux_s2_v I__8738 (
            .O(N__40619),
            .I(N__40603));
    LocalMux I__8737 (
            .O(N__40616),
            .I(N__40603));
    InMux I__8736 (
            .O(N__40615),
            .I(N__40600));
    Span4Mux_h I__8735 (
            .O(N__40610),
            .I(N__40597));
    Span4Mux_h I__8734 (
            .O(N__40603),
            .I(N__40594));
    LocalMux I__8733 (
            .O(N__40600),
            .I(\phase_controller_inst1.stoper_hc.hc_time_passed ));
    Odrv4 I__8732 (
            .O(N__40597),
            .I(\phase_controller_inst1.stoper_hc.hc_time_passed ));
    Odrv4 I__8731 (
            .O(N__40594),
            .I(\phase_controller_inst1.stoper_hc.hc_time_passed ));
    InMux I__8730 (
            .O(N__40587),
            .I(N__40583));
    InMux I__8729 (
            .O(N__40586),
            .I(N__40580));
    LocalMux I__8728 (
            .O(N__40583),
            .I(\phase_controller_inst1.stoper_hc.N_45 ));
    LocalMux I__8727 (
            .O(N__40580),
            .I(\phase_controller_inst1.stoper_hc.N_45 ));
    InMux I__8726 (
            .O(N__40575),
            .I(N__40571));
    InMux I__8725 (
            .O(N__40574),
            .I(N__40567));
    LocalMux I__8724 (
            .O(N__40571),
            .I(N__40564));
    InMux I__8723 (
            .O(N__40570),
            .I(N__40561));
    LocalMux I__8722 (
            .O(N__40567),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    Odrv4 I__8721 (
            .O(N__40564),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    LocalMux I__8720 (
            .O(N__40561),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ));
    CascadeMux I__8719 (
            .O(N__40554),
            .I(N__40547));
    InMux I__8718 (
            .O(N__40553),
            .I(N__40544));
    InMux I__8717 (
            .O(N__40552),
            .I(N__40539));
    InMux I__8716 (
            .O(N__40551),
            .I(N__40539));
    InMux I__8715 (
            .O(N__40550),
            .I(N__40536));
    InMux I__8714 (
            .O(N__40547),
            .I(N__40533));
    LocalMux I__8713 (
            .O(N__40544),
            .I(N__40530));
    LocalMux I__8712 (
            .O(N__40539),
            .I(N__40527));
    LocalMux I__8711 (
            .O(N__40536),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__8710 (
            .O(N__40533),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8709 (
            .O(N__40530),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    Odrv4 I__8708 (
            .O(N__40527),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__8707 (
            .O(N__40518),
            .I(N__40513));
    InMux I__8706 (
            .O(N__40517),
            .I(N__40508));
    InMux I__8705 (
            .O(N__40516),
            .I(N__40505));
    LocalMux I__8704 (
            .O(N__40513),
            .I(N__40502));
    InMux I__8703 (
            .O(N__40512),
            .I(N__40497));
    InMux I__8702 (
            .O(N__40511),
            .I(N__40497));
    LocalMux I__8701 (
            .O(N__40508),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__8700 (
            .O(N__40505),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__8699 (
            .O(N__40502),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__8698 (
            .O(N__40497),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    CascadeMux I__8697 (
            .O(N__40488),
            .I(N__40483));
    CascadeMux I__8696 (
            .O(N__40487),
            .I(N__40480));
    InMux I__8695 (
            .O(N__40486),
            .I(N__40477));
    InMux I__8694 (
            .O(N__40483),
            .I(N__40474));
    InMux I__8693 (
            .O(N__40480),
            .I(N__40471));
    LocalMux I__8692 (
            .O(N__40477),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__8691 (
            .O(N__40474),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__8690 (
            .O(N__40471),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    InMux I__8689 (
            .O(N__40464),
            .I(N__40460));
    InMux I__8688 (
            .O(N__40463),
            .I(N__40457));
    LocalMux I__8687 (
            .O(N__40460),
            .I(N__40454));
    LocalMux I__8686 (
            .O(N__40457),
            .I(N__40451));
    Odrv4 I__8685 (
            .O(N__40454),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    Odrv12 I__8684 (
            .O(N__40451),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ));
    InMux I__8683 (
            .O(N__40446),
            .I(N__40443));
    LocalMux I__8682 (
            .O(N__40443),
            .I(\phase_controller_inst1.stoper_hc.N_46 ));
    CascadeMux I__8681 (
            .O(N__40440),
            .I(\phase_controller_inst1.stoper_hc.N_46_cascade_ ));
    CEMux I__8680 (
            .O(N__40437),
            .I(N__40434));
    LocalMux I__8679 (
            .O(N__40434),
            .I(N__40431));
    Odrv4 I__8678 (
            .O(N__40431),
            .I(\phase_controller_inst1.stoper_hc.N_46_0 ));
    CascadeMux I__8677 (
            .O(N__40428),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ));
    CascadeMux I__8676 (
            .O(N__40425),
            .I(\current_shift_inst.PI_CTRL.N_287_cascade_ ));
    InMux I__8675 (
            .O(N__40422),
            .I(N__40419));
    LocalMux I__8674 (
            .O(N__40419),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ));
    InMux I__8673 (
            .O(N__40416),
            .I(N__40413));
    LocalMux I__8672 (
            .O(N__40413),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ));
    CascadeMux I__8671 (
            .O(N__40410),
            .I(N__40407));
    InMux I__8670 (
            .O(N__40407),
            .I(N__40402));
    InMux I__8669 (
            .O(N__40406),
            .I(N__40399));
    InMux I__8668 (
            .O(N__40405),
            .I(N__40396));
    LocalMux I__8667 (
            .O(N__40402),
            .I(N__40391));
    LocalMux I__8666 (
            .O(N__40399),
            .I(N__40391));
    LocalMux I__8665 (
            .O(N__40396),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv4 I__8664 (
            .O(N__40391),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__8663 (
            .O(N__40386),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__8662 (
            .O(N__40383),
            .I(N__40376));
    InMux I__8661 (
            .O(N__40382),
            .I(N__40376));
    InMux I__8660 (
            .O(N__40381),
            .I(N__40373));
    LocalMux I__8659 (
            .O(N__40376),
            .I(N__40370));
    LocalMux I__8658 (
            .O(N__40373),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv4 I__8657 (
            .O(N__40370),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__8656 (
            .O(N__40365),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__8655 (
            .O(N__40362),
            .I(N__40358));
    InMux I__8654 (
            .O(N__40361),
            .I(N__40355));
    LocalMux I__8653 (
            .O(N__40358),
            .I(N__40352));
    LocalMux I__8652 (
            .O(N__40355),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv4 I__8651 (
            .O(N__40352),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    InMux I__8650 (
            .O(N__40347),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__8649 (
            .O(N__40344),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    CascadeMux I__8648 (
            .O(N__40341),
            .I(N__40338));
    InMux I__8647 (
            .O(N__40338),
            .I(N__40334));
    InMux I__8646 (
            .O(N__40337),
            .I(N__40331));
    LocalMux I__8645 (
            .O(N__40334),
            .I(N__40328));
    LocalMux I__8644 (
            .O(N__40331),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__8643 (
            .O(N__40328),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CEMux I__8642 (
            .O(N__40323),
            .I(N__40319));
    CEMux I__8641 (
            .O(N__40322),
            .I(N__40316));
    LocalMux I__8640 (
            .O(N__40319),
            .I(N__40311));
    LocalMux I__8639 (
            .O(N__40316),
            .I(N__40308));
    CEMux I__8638 (
            .O(N__40315),
            .I(N__40305));
    CEMux I__8637 (
            .O(N__40314),
            .I(N__40302));
    Span4Mux_v I__8636 (
            .O(N__40311),
            .I(N__40299));
    Span4Mux_h I__8635 (
            .O(N__40308),
            .I(N__40296));
    LocalMux I__8634 (
            .O(N__40305),
            .I(N__40291));
    LocalMux I__8633 (
            .O(N__40302),
            .I(N__40291));
    Odrv4 I__8632 (
            .O(N__40299),
            .I(\current_shift_inst.timer_s1.N_340_i ));
    Odrv4 I__8631 (
            .O(N__40296),
            .I(\current_shift_inst.timer_s1.N_340_i ));
    Odrv4 I__8630 (
            .O(N__40291),
            .I(\current_shift_inst.timer_s1.N_340_i ));
    CascadeMux I__8629 (
            .O(N__40284),
            .I(N__40281));
    InMux I__8628 (
            .O(N__40281),
            .I(N__40275));
    InMux I__8627 (
            .O(N__40280),
            .I(N__40275));
    LocalMux I__8626 (
            .O(N__40275),
            .I(N__40272));
    Span4Mux_v I__8625 (
            .O(N__40272),
            .I(N__40269));
    Odrv4 I__8624 (
            .O(N__40269),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ));
    CascadeMux I__8623 (
            .O(N__40266),
            .I(N__40262));
    InMux I__8622 (
            .O(N__40265),
            .I(N__40257));
    InMux I__8621 (
            .O(N__40262),
            .I(N__40257));
    LocalMux I__8620 (
            .O(N__40257),
            .I(N__40254));
    Odrv12 I__8619 (
            .O(N__40254),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ));
    CascadeMux I__8618 (
            .O(N__40251),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_));
    InMux I__8617 (
            .O(N__40248),
            .I(N__40245));
    LocalMux I__8616 (
            .O(N__40245),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ));
    InMux I__8615 (
            .O(N__40242),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__8614 (
            .O(N__40239),
            .I(N__40232));
    InMux I__8613 (
            .O(N__40238),
            .I(N__40232));
    InMux I__8612 (
            .O(N__40237),
            .I(N__40229));
    LocalMux I__8611 (
            .O(N__40232),
            .I(N__40226));
    LocalMux I__8610 (
            .O(N__40229),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv4 I__8609 (
            .O(N__40226),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__8608 (
            .O(N__40221),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__8607 (
            .O(N__40218),
            .I(N__40211));
    InMux I__8606 (
            .O(N__40217),
            .I(N__40211));
    InMux I__8605 (
            .O(N__40216),
            .I(N__40208));
    LocalMux I__8604 (
            .O(N__40211),
            .I(N__40205));
    LocalMux I__8603 (
            .O(N__40208),
            .I(N__40200));
    Span4Mux_h I__8602 (
            .O(N__40205),
            .I(N__40200));
    Odrv4 I__8601 (
            .O(N__40200),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__8600 (
            .O(N__40197),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    CascadeMux I__8599 (
            .O(N__40194),
            .I(N__40190));
    InMux I__8598 (
            .O(N__40193),
            .I(N__40186));
    InMux I__8597 (
            .O(N__40190),
            .I(N__40183));
    InMux I__8596 (
            .O(N__40189),
            .I(N__40180));
    LocalMux I__8595 (
            .O(N__40186),
            .I(N__40175));
    LocalMux I__8594 (
            .O(N__40183),
            .I(N__40175));
    LocalMux I__8593 (
            .O(N__40180),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv4 I__8592 (
            .O(N__40175),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__8591 (
            .O(N__40170),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    CascadeMux I__8590 (
            .O(N__40167),
            .I(N__40163));
    InMux I__8589 (
            .O(N__40166),
            .I(N__40159));
    InMux I__8588 (
            .O(N__40163),
            .I(N__40156));
    InMux I__8587 (
            .O(N__40162),
            .I(N__40153));
    LocalMux I__8586 (
            .O(N__40159),
            .I(N__40148));
    LocalMux I__8585 (
            .O(N__40156),
            .I(N__40148));
    LocalMux I__8584 (
            .O(N__40153),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv4 I__8583 (
            .O(N__40148),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__8582 (
            .O(N__40143),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    CascadeMux I__8581 (
            .O(N__40140),
            .I(N__40136));
    CascadeMux I__8580 (
            .O(N__40139),
            .I(N__40133));
    InMux I__8579 (
            .O(N__40136),
            .I(N__40127));
    InMux I__8578 (
            .O(N__40133),
            .I(N__40127));
    InMux I__8577 (
            .O(N__40132),
            .I(N__40124));
    LocalMux I__8576 (
            .O(N__40127),
            .I(N__40121));
    LocalMux I__8575 (
            .O(N__40124),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__8574 (
            .O(N__40121),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__8573 (
            .O(N__40116),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    CascadeMux I__8572 (
            .O(N__40113),
            .I(N__40109));
    CascadeMux I__8571 (
            .O(N__40112),
            .I(N__40106));
    InMux I__8570 (
            .O(N__40109),
            .I(N__40100));
    InMux I__8569 (
            .O(N__40106),
            .I(N__40100));
    InMux I__8568 (
            .O(N__40105),
            .I(N__40097));
    LocalMux I__8567 (
            .O(N__40100),
            .I(N__40094));
    LocalMux I__8566 (
            .O(N__40097),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__8565 (
            .O(N__40094),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__8564 (
            .O(N__40089),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    CascadeMux I__8563 (
            .O(N__40086),
            .I(N__40083));
    InMux I__8562 (
            .O(N__40083),
            .I(N__40078));
    InMux I__8561 (
            .O(N__40082),
            .I(N__40075));
    InMux I__8560 (
            .O(N__40081),
            .I(N__40072));
    LocalMux I__8559 (
            .O(N__40078),
            .I(N__40067));
    LocalMux I__8558 (
            .O(N__40075),
            .I(N__40067));
    LocalMux I__8557 (
            .O(N__40072),
            .I(N__40062));
    Span4Mux_v I__8556 (
            .O(N__40067),
            .I(N__40062));
    Odrv4 I__8555 (
            .O(N__40062),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__8554 (
            .O(N__40059),
            .I(bfn_16_17_0_));
    CascadeMux I__8553 (
            .O(N__40056),
            .I(N__40053));
    InMux I__8552 (
            .O(N__40053),
            .I(N__40049));
    InMux I__8551 (
            .O(N__40052),
            .I(N__40046));
    LocalMux I__8550 (
            .O(N__40049),
            .I(N__40040));
    LocalMux I__8549 (
            .O(N__40046),
            .I(N__40040));
    InMux I__8548 (
            .O(N__40045),
            .I(N__40037));
    Span4Mux_v I__8547 (
            .O(N__40040),
            .I(N__40034));
    LocalMux I__8546 (
            .O(N__40037),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv4 I__8545 (
            .O(N__40034),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__8544 (
            .O(N__40029),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    CascadeMux I__8543 (
            .O(N__40026),
            .I(N__40022));
    CascadeMux I__8542 (
            .O(N__40025),
            .I(N__40019));
    InMux I__8541 (
            .O(N__40022),
            .I(N__40016));
    InMux I__8540 (
            .O(N__40019),
            .I(N__40012));
    LocalMux I__8539 (
            .O(N__40016),
            .I(N__40009));
    InMux I__8538 (
            .O(N__40015),
            .I(N__40006));
    LocalMux I__8537 (
            .O(N__40012),
            .I(N__40003));
    Span4Mux_v I__8536 (
            .O(N__40009),
            .I(N__40000));
    LocalMux I__8535 (
            .O(N__40006),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv12 I__8534 (
            .O(N__40003),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv4 I__8533 (
            .O(N__40000),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__8532 (
            .O(N__39993),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__8531 (
            .O(N__39990),
            .I(N__39983));
    InMux I__8530 (
            .O(N__39989),
            .I(N__39983));
    InMux I__8529 (
            .O(N__39988),
            .I(N__39980));
    LocalMux I__8528 (
            .O(N__39983),
            .I(N__39977));
    LocalMux I__8527 (
            .O(N__39980),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__8526 (
            .O(N__39977),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__8525 (
            .O(N__39972),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__8524 (
            .O(N__39969),
            .I(N__39962));
    InMux I__8523 (
            .O(N__39968),
            .I(N__39962));
    InMux I__8522 (
            .O(N__39967),
            .I(N__39959));
    LocalMux I__8521 (
            .O(N__39962),
            .I(N__39956));
    LocalMux I__8520 (
            .O(N__39959),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv12 I__8519 (
            .O(N__39956),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__8518 (
            .O(N__39951),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    CascadeMux I__8517 (
            .O(N__39948),
            .I(N__39944));
    InMux I__8516 (
            .O(N__39947),
            .I(N__39940));
    InMux I__8515 (
            .O(N__39944),
            .I(N__39937));
    InMux I__8514 (
            .O(N__39943),
            .I(N__39934));
    LocalMux I__8513 (
            .O(N__39940),
            .I(N__39929));
    LocalMux I__8512 (
            .O(N__39937),
            .I(N__39929));
    LocalMux I__8511 (
            .O(N__39934),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__8510 (
            .O(N__39929),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__8509 (
            .O(N__39924),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    CascadeMux I__8508 (
            .O(N__39921),
            .I(N__39917));
    CascadeMux I__8507 (
            .O(N__39920),
            .I(N__39914));
    InMux I__8506 (
            .O(N__39917),
            .I(N__39908));
    InMux I__8505 (
            .O(N__39914),
            .I(N__39908));
    InMux I__8504 (
            .O(N__39913),
            .I(N__39905));
    LocalMux I__8503 (
            .O(N__39908),
            .I(N__39902));
    LocalMux I__8502 (
            .O(N__39905),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv4 I__8501 (
            .O(N__39902),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__8500 (
            .O(N__39897),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    CascadeMux I__8499 (
            .O(N__39894),
            .I(N__39890));
    CascadeMux I__8498 (
            .O(N__39893),
            .I(N__39887));
    InMux I__8497 (
            .O(N__39890),
            .I(N__39881));
    InMux I__8496 (
            .O(N__39887),
            .I(N__39881));
    InMux I__8495 (
            .O(N__39886),
            .I(N__39878));
    LocalMux I__8494 (
            .O(N__39881),
            .I(N__39875));
    LocalMux I__8493 (
            .O(N__39878),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__8492 (
            .O(N__39875),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__8491 (
            .O(N__39870),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__8490 (
            .O(N__39867),
            .I(N__39860));
    InMux I__8489 (
            .O(N__39866),
            .I(N__39860));
    InMux I__8488 (
            .O(N__39865),
            .I(N__39857));
    LocalMux I__8487 (
            .O(N__39860),
            .I(N__39854));
    LocalMux I__8486 (
            .O(N__39857),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv4 I__8485 (
            .O(N__39854),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__8484 (
            .O(N__39849),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    CascadeMux I__8483 (
            .O(N__39846),
            .I(N__39843));
    InMux I__8482 (
            .O(N__39843),
            .I(N__39838));
    InMux I__8481 (
            .O(N__39842),
            .I(N__39835));
    InMux I__8480 (
            .O(N__39841),
            .I(N__39832));
    LocalMux I__8479 (
            .O(N__39838),
            .I(N__39827));
    LocalMux I__8478 (
            .O(N__39835),
            .I(N__39827));
    LocalMux I__8477 (
            .O(N__39832),
            .I(N__39822));
    Span4Mux_v I__8476 (
            .O(N__39827),
            .I(N__39822));
    Odrv4 I__8475 (
            .O(N__39822),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__8474 (
            .O(N__39819),
            .I(bfn_16_16_0_));
    CascadeMux I__8473 (
            .O(N__39816),
            .I(N__39812));
    CascadeMux I__8472 (
            .O(N__39815),
            .I(N__39809));
    InMux I__8471 (
            .O(N__39812),
            .I(N__39806));
    InMux I__8470 (
            .O(N__39809),
            .I(N__39803));
    LocalMux I__8469 (
            .O(N__39806),
            .I(N__39799));
    LocalMux I__8468 (
            .O(N__39803),
            .I(N__39796));
    InMux I__8467 (
            .O(N__39802),
            .I(N__39793));
    Span4Mux_h I__8466 (
            .O(N__39799),
            .I(N__39788));
    Span4Mux_v I__8465 (
            .O(N__39796),
            .I(N__39788));
    LocalMux I__8464 (
            .O(N__39793),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv4 I__8463 (
            .O(N__39788),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__8462 (
            .O(N__39783),
            .I(N__39779));
    CascadeMux I__8461 (
            .O(N__39782),
            .I(N__39776));
    LocalMux I__8460 (
            .O(N__39779),
            .I(N__39773));
    InMux I__8459 (
            .O(N__39776),
            .I(N__39769));
    Span4Mux_h I__8458 (
            .O(N__39773),
            .I(N__39766));
    InMux I__8457 (
            .O(N__39772),
            .I(N__39763));
    LocalMux I__8456 (
            .O(N__39769),
            .I(N__39760));
    Odrv4 I__8455 (
            .O(N__39766),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__8454 (
            .O(N__39763),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv12 I__8453 (
            .O(N__39760),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__8452 (
            .O(N__39753),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__8451 (
            .O(N__39750),
            .I(N__39743));
    InMux I__8450 (
            .O(N__39749),
            .I(N__39743));
    InMux I__8449 (
            .O(N__39748),
            .I(N__39740));
    LocalMux I__8448 (
            .O(N__39743),
            .I(N__39737));
    LocalMux I__8447 (
            .O(N__39740),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv12 I__8446 (
            .O(N__39737),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__8445 (
            .O(N__39732),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__8444 (
            .O(N__39729),
            .I(N__39722));
    InMux I__8443 (
            .O(N__39728),
            .I(N__39722));
    InMux I__8442 (
            .O(N__39727),
            .I(N__39719));
    LocalMux I__8441 (
            .O(N__39722),
            .I(N__39716));
    LocalMux I__8440 (
            .O(N__39719),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv12 I__8439 (
            .O(N__39716),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__8438 (
            .O(N__39711),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    CascadeMux I__8437 (
            .O(N__39708),
            .I(N__39704));
    CascadeMux I__8436 (
            .O(N__39707),
            .I(N__39701));
    InMux I__8435 (
            .O(N__39704),
            .I(N__39695));
    InMux I__8434 (
            .O(N__39701),
            .I(N__39695));
    InMux I__8433 (
            .O(N__39700),
            .I(N__39692));
    LocalMux I__8432 (
            .O(N__39695),
            .I(N__39689));
    LocalMux I__8431 (
            .O(N__39692),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__8430 (
            .O(N__39689),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__8429 (
            .O(N__39684),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    CascadeMux I__8428 (
            .O(N__39681),
            .I(N__39677));
    CascadeMux I__8427 (
            .O(N__39680),
            .I(N__39674));
    InMux I__8426 (
            .O(N__39677),
            .I(N__39668));
    InMux I__8425 (
            .O(N__39674),
            .I(N__39668));
    InMux I__8424 (
            .O(N__39673),
            .I(N__39665));
    LocalMux I__8423 (
            .O(N__39668),
            .I(N__39662));
    LocalMux I__8422 (
            .O(N__39665),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv4 I__8421 (
            .O(N__39662),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__8420 (
            .O(N__39657),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__8419 (
            .O(N__39654),
            .I(N__39647));
    InMux I__8418 (
            .O(N__39653),
            .I(N__39647));
    InMux I__8417 (
            .O(N__39652),
            .I(N__39644));
    LocalMux I__8416 (
            .O(N__39647),
            .I(N__39641));
    LocalMux I__8415 (
            .O(N__39644),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__8414 (
            .O(N__39641),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__8413 (
            .O(N__39636),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__8412 (
            .O(N__39633),
            .I(N__39626));
    InMux I__8411 (
            .O(N__39632),
            .I(N__39626));
    InMux I__8410 (
            .O(N__39631),
            .I(N__39623));
    LocalMux I__8409 (
            .O(N__39626),
            .I(N__39620));
    LocalMux I__8408 (
            .O(N__39623),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__8407 (
            .O(N__39620),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__8406 (
            .O(N__39615),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    CascadeMux I__8405 (
            .O(N__39612),
            .I(N__39608));
    CascadeMux I__8404 (
            .O(N__39611),
            .I(N__39605));
    InMux I__8403 (
            .O(N__39608),
            .I(N__39601));
    InMux I__8402 (
            .O(N__39605),
            .I(N__39598));
    InMux I__8401 (
            .O(N__39604),
            .I(N__39595));
    LocalMux I__8400 (
            .O(N__39601),
            .I(N__39590));
    LocalMux I__8399 (
            .O(N__39598),
            .I(N__39590));
    LocalMux I__8398 (
            .O(N__39595),
            .I(N__39585));
    Span4Mux_v I__8397 (
            .O(N__39590),
            .I(N__39585));
    Odrv4 I__8396 (
            .O(N__39585),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__8395 (
            .O(N__39582),
            .I(bfn_16_15_0_));
    InMux I__8394 (
            .O(N__39579),
            .I(N__39574));
    InMux I__8393 (
            .O(N__39578),
            .I(N__39571));
    InMux I__8392 (
            .O(N__39577),
            .I(N__39568));
    LocalMux I__8391 (
            .O(N__39574),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    LocalMux I__8390 (
            .O(N__39571),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    LocalMux I__8389 (
            .O(N__39568),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    InMux I__8388 (
            .O(N__39561),
            .I(N__39556));
    InMux I__8387 (
            .O(N__39560),
            .I(N__39553));
    InMux I__8386 (
            .O(N__39559),
            .I(N__39550));
    LocalMux I__8385 (
            .O(N__39556),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__8384 (
            .O(N__39553),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    LocalMux I__8383 (
            .O(N__39550),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    InMux I__8382 (
            .O(N__39543),
            .I(N__39540));
    LocalMux I__8381 (
            .O(N__39540),
            .I(N__39536));
    InMux I__8380 (
            .O(N__39539),
            .I(N__39532));
    Span4Mux_h I__8379 (
            .O(N__39536),
            .I(N__39529));
    InMux I__8378 (
            .O(N__39535),
            .I(N__39526));
    LocalMux I__8377 (
            .O(N__39532),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    Odrv4 I__8376 (
            .O(N__39529),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__8375 (
            .O(N__39526),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__8374 (
            .O(N__39519),
            .I(N__39514));
    InMux I__8373 (
            .O(N__39518),
            .I(N__39511));
    InMux I__8372 (
            .O(N__39517),
            .I(N__39508));
    LocalMux I__8371 (
            .O(N__39514),
            .I(N__39505));
    LocalMux I__8370 (
            .O(N__39511),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    LocalMux I__8369 (
            .O(N__39508),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    Odrv4 I__8368 (
            .O(N__39505),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    InMux I__8367 (
            .O(N__39498),
            .I(N__39492));
    InMux I__8366 (
            .O(N__39497),
            .I(N__39492));
    LocalMux I__8365 (
            .O(N__39492),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ));
    CascadeMux I__8364 (
            .O(N__39489),
            .I(N__39486));
    InMux I__8363 (
            .O(N__39486),
            .I(N__39480));
    InMux I__8362 (
            .O(N__39485),
            .I(N__39480));
    LocalMux I__8361 (
            .O(N__39480),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ));
    InMux I__8360 (
            .O(N__39477),
            .I(N__39473));
    InMux I__8359 (
            .O(N__39476),
            .I(N__39469));
    LocalMux I__8358 (
            .O(N__39473),
            .I(N__39466));
    InMux I__8357 (
            .O(N__39472),
            .I(N__39463));
    LocalMux I__8356 (
            .O(N__39469),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    Odrv4 I__8355 (
            .O(N__39466),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    LocalMux I__8354 (
            .O(N__39463),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    InMux I__8353 (
            .O(N__39456),
            .I(N__39452));
    CascadeMux I__8352 (
            .O(N__39455),
            .I(N__39449));
    LocalMux I__8351 (
            .O(N__39452),
            .I(N__39446));
    InMux I__8350 (
            .O(N__39449),
            .I(N__39442));
    Span4Mux_h I__8349 (
            .O(N__39446),
            .I(N__39439));
    InMux I__8348 (
            .O(N__39445),
            .I(N__39436));
    LocalMux I__8347 (
            .O(N__39442),
            .I(N__39433));
    Odrv4 I__8346 (
            .O(N__39439),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__8345 (
            .O(N__39436),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__8344 (
            .O(N__39433),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__8343 (
            .O(N__39426),
            .I(bfn_16_14_0_));
    InMux I__8342 (
            .O(N__39423),
            .I(N__39417));
    InMux I__8341 (
            .O(N__39422),
            .I(N__39417));
    LocalMux I__8340 (
            .O(N__39417),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ));
    InMux I__8339 (
            .O(N__39414),
            .I(N__39407));
    InMux I__8338 (
            .O(N__39413),
            .I(N__39407));
    InMux I__8337 (
            .O(N__39412),
            .I(N__39404));
    LocalMux I__8336 (
            .O(N__39407),
            .I(N__39401));
    LocalMux I__8335 (
            .O(N__39404),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    Odrv4 I__8334 (
            .O(N__39401),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ));
    InMux I__8333 (
            .O(N__39396),
            .I(N__39390));
    InMux I__8332 (
            .O(N__39395),
            .I(N__39390));
    LocalMux I__8331 (
            .O(N__39390),
            .I(N__39386));
    InMux I__8330 (
            .O(N__39389),
            .I(N__39383));
    Span4Mux_v I__8329 (
            .O(N__39386),
            .I(N__39380));
    LocalMux I__8328 (
            .O(N__39383),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    Odrv4 I__8327 (
            .O(N__39380),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ));
    InMux I__8326 (
            .O(N__39375),
            .I(N__39372));
    LocalMux I__8325 (
            .O(N__39372),
            .I(N__39369));
    Odrv4 I__8324 (
            .O(N__39369),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ));
    InMux I__8323 (
            .O(N__39366),
            .I(N__39363));
    LocalMux I__8322 (
            .O(N__39363),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ));
    InMux I__8321 (
            .O(N__39360),
            .I(N__39357));
    LocalMux I__8320 (
            .O(N__39357),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    InMux I__8319 (
            .O(N__39354),
            .I(N__39347));
    InMux I__8318 (
            .O(N__39353),
            .I(N__39347));
    InMux I__8317 (
            .O(N__39352),
            .I(N__39344));
    LocalMux I__8316 (
            .O(N__39347),
            .I(N__39341));
    LocalMux I__8315 (
            .O(N__39344),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    Odrv4 I__8314 (
            .O(N__39341),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ));
    CascadeMux I__8313 (
            .O(N__39336),
            .I(N__39332));
    InMux I__8312 (
            .O(N__39335),
            .I(N__39326));
    InMux I__8311 (
            .O(N__39332),
            .I(N__39326));
    InMux I__8310 (
            .O(N__39331),
            .I(N__39323));
    LocalMux I__8309 (
            .O(N__39326),
            .I(N__39320));
    LocalMux I__8308 (
            .O(N__39323),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    Odrv4 I__8307 (
            .O(N__39320),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ));
    InMux I__8306 (
            .O(N__39315),
            .I(N__39312));
    LocalMux I__8305 (
            .O(N__39312),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ));
    CascadeMux I__8304 (
            .O(N__39309),
            .I(elapsed_time_ns_1_RNI13CN9_0_14_cascade_));
    InMux I__8303 (
            .O(N__39306),
            .I(N__39303));
    LocalMux I__8302 (
            .O(N__39303),
            .I(N__39300));
    Odrv4 I__8301 (
            .O(N__39300),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ));
    InMux I__8300 (
            .O(N__39297),
            .I(N__39291));
    InMux I__8299 (
            .O(N__39296),
            .I(N__39291));
    LocalMux I__8298 (
            .O(N__39291),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ));
    CascadeMux I__8297 (
            .O(N__39288),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_ ));
    InMux I__8296 (
            .O(N__39285),
            .I(N__39282));
    LocalMux I__8295 (
            .O(N__39282),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    CascadeMux I__8294 (
            .O(N__39279),
            .I(N__39276));
    InMux I__8293 (
            .O(N__39276),
            .I(N__39273));
    LocalMux I__8292 (
            .O(N__39273),
            .I(N__39270));
    Odrv4 I__8291 (
            .O(N__39270),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt20 ));
    InMux I__8290 (
            .O(N__39267),
            .I(N__39264));
    LocalMux I__8289 (
            .O(N__39264),
            .I(N__39261));
    Odrv4 I__8288 (
            .O(N__39261),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt24 ));
    CascadeMux I__8287 (
            .O(N__39258),
            .I(N__39255));
    InMux I__8286 (
            .O(N__39255),
            .I(N__39252));
    LocalMux I__8285 (
            .O(N__39252),
            .I(N__39249));
    Span4Mux_v I__8284 (
            .O(N__39249),
            .I(N__39246));
    Odrv4 I__8283 (
            .O(N__39246),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ));
    InMux I__8282 (
            .O(N__39243),
            .I(N__39240));
    LocalMux I__8281 (
            .O(N__39240),
            .I(N__39237));
    Span4Mux_h I__8280 (
            .O(N__39237),
            .I(N__39234));
    Odrv4 I__8279 (
            .O(N__39234),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ));
    CascadeMux I__8278 (
            .O(N__39231),
            .I(N__39228));
    InMux I__8277 (
            .O(N__39228),
            .I(N__39225));
    LocalMux I__8276 (
            .O(N__39225),
            .I(N__39222));
    Span4Mux_h I__8275 (
            .O(N__39222),
            .I(N__39219));
    Odrv4 I__8274 (
            .O(N__39219),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt28 ));
    InMux I__8273 (
            .O(N__39216),
            .I(N__39213));
    LocalMux I__8272 (
            .O(N__39213),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ));
    CascadeMux I__8271 (
            .O(N__39210),
            .I(N__39207));
    InMux I__8270 (
            .O(N__39207),
            .I(N__39204));
    LocalMux I__8269 (
            .O(N__39204),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt30 ));
    InMux I__8268 (
            .O(N__39201),
            .I(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ));
    CascadeMux I__8267 (
            .O(N__39198),
            .I(N__39195));
    InMux I__8266 (
            .O(N__39195),
            .I(N__39192));
    LocalMux I__8265 (
            .O(N__39192),
            .I(\phase_controller_inst1.stoper_hc.un4_running_lt18 ));
    InMux I__8264 (
            .O(N__39189),
            .I(N__39185));
    InMux I__8263 (
            .O(N__39188),
            .I(N__39182));
    LocalMux I__8262 (
            .O(N__39185),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    LocalMux I__8261 (
            .O(N__39182),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ));
    InMux I__8260 (
            .O(N__39177),
            .I(N__39174));
    LocalMux I__8259 (
            .O(N__39174),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ));
    InMux I__8258 (
            .O(N__39171),
            .I(N__39167));
    InMux I__8257 (
            .O(N__39170),
            .I(N__39164));
    LocalMux I__8256 (
            .O(N__39167),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    LocalMux I__8255 (
            .O(N__39164),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ));
    CascadeMux I__8254 (
            .O(N__39159),
            .I(N__39156));
    InMux I__8253 (
            .O(N__39156),
            .I(N__39153));
    LocalMux I__8252 (
            .O(N__39153),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ));
    InMux I__8251 (
            .O(N__39150),
            .I(N__39146));
    InMux I__8250 (
            .O(N__39149),
            .I(N__39143));
    LocalMux I__8249 (
            .O(N__39146),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    LocalMux I__8248 (
            .O(N__39143),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ));
    CascadeMux I__8247 (
            .O(N__39138),
            .I(N__39135));
    InMux I__8246 (
            .O(N__39135),
            .I(N__39132));
    LocalMux I__8245 (
            .O(N__39132),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ));
    InMux I__8244 (
            .O(N__39129),
            .I(N__39125));
    InMux I__8243 (
            .O(N__39128),
            .I(N__39122));
    LocalMux I__8242 (
            .O(N__39125),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    LocalMux I__8241 (
            .O(N__39122),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ));
    InMux I__8240 (
            .O(N__39117),
            .I(N__39114));
    LocalMux I__8239 (
            .O(N__39114),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ));
    InMux I__8238 (
            .O(N__39111),
            .I(N__39108));
    LocalMux I__8237 (
            .O(N__39108),
            .I(N__39105));
    Odrv4 I__8236 (
            .O(N__39105),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ));
    InMux I__8235 (
            .O(N__39102),
            .I(N__39098));
    InMux I__8234 (
            .O(N__39101),
            .I(N__39095));
    LocalMux I__8233 (
            .O(N__39098),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    LocalMux I__8232 (
            .O(N__39095),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ));
    CascadeMux I__8231 (
            .O(N__39090),
            .I(N__39087));
    InMux I__8230 (
            .O(N__39087),
            .I(N__39084));
    LocalMux I__8229 (
            .O(N__39084),
            .I(N__39081));
    Odrv4 I__8228 (
            .O(N__39081),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ));
    InMux I__8227 (
            .O(N__39078),
            .I(N__39074));
    InMux I__8226 (
            .O(N__39077),
            .I(N__39071));
    LocalMux I__8225 (
            .O(N__39074),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    LocalMux I__8224 (
            .O(N__39071),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ));
    CascadeMux I__8223 (
            .O(N__39066),
            .I(N__39063));
    InMux I__8222 (
            .O(N__39063),
            .I(N__39060));
    LocalMux I__8221 (
            .O(N__39060),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ));
    InMux I__8220 (
            .O(N__39057),
            .I(N__39054));
    LocalMux I__8219 (
            .O(N__39054),
            .I(N__39051));
    Span4Mux_h I__8218 (
            .O(N__39051),
            .I(N__39048));
    Odrv4 I__8217 (
            .O(N__39048),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ));
    InMux I__8216 (
            .O(N__39045),
            .I(N__39041));
    InMux I__8215 (
            .O(N__39044),
            .I(N__39038));
    LocalMux I__8214 (
            .O(N__39041),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    LocalMux I__8213 (
            .O(N__39038),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ));
    CascadeMux I__8212 (
            .O(N__39033),
            .I(N__39030));
    InMux I__8211 (
            .O(N__39030),
            .I(N__39027));
    LocalMux I__8210 (
            .O(N__39027),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ));
    InMux I__8209 (
            .O(N__39024),
            .I(N__39020));
    InMux I__8208 (
            .O(N__39023),
            .I(N__39017));
    LocalMux I__8207 (
            .O(N__39020),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    LocalMux I__8206 (
            .O(N__39017),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ));
    CascadeMux I__8205 (
            .O(N__39012),
            .I(N__39009));
    InMux I__8204 (
            .O(N__39009),
            .I(N__39006));
    LocalMux I__8203 (
            .O(N__39006),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ));
    InMux I__8202 (
            .O(N__39003),
            .I(N__38999));
    InMux I__8201 (
            .O(N__39002),
            .I(N__38996));
    LocalMux I__8200 (
            .O(N__38999),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    LocalMux I__8199 (
            .O(N__38996),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ));
    InMux I__8198 (
            .O(N__38991),
            .I(N__38988));
    LocalMux I__8197 (
            .O(N__38988),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ));
    InMux I__8196 (
            .O(N__38985),
            .I(N__38981));
    InMux I__8195 (
            .O(N__38984),
            .I(N__38978));
    LocalMux I__8194 (
            .O(N__38981),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    LocalMux I__8193 (
            .O(N__38978),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ));
    CascadeMux I__8192 (
            .O(N__38973),
            .I(N__38970));
    InMux I__8191 (
            .O(N__38970),
            .I(N__38967));
    LocalMux I__8190 (
            .O(N__38967),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ));
    InMux I__8189 (
            .O(N__38964),
            .I(N__38960));
    InMux I__8188 (
            .O(N__38963),
            .I(N__38957));
    LocalMux I__8187 (
            .O(N__38960),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    LocalMux I__8186 (
            .O(N__38957),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ));
    CascadeMux I__8185 (
            .O(N__38952),
            .I(N__38949));
    InMux I__8184 (
            .O(N__38949),
            .I(N__38946));
    LocalMux I__8183 (
            .O(N__38946),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ));
    InMux I__8182 (
            .O(N__38943),
            .I(N__38940));
    LocalMux I__8181 (
            .O(N__38940),
            .I(N__38937));
    Span4Mux_v I__8180 (
            .O(N__38937),
            .I(N__38934));
    Odrv4 I__8179 (
            .O(N__38934),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ));
    InMux I__8178 (
            .O(N__38931),
            .I(N__38927));
    InMux I__8177 (
            .O(N__38930),
            .I(N__38924));
    LocalMux I__8176 (
            .O(N__38927),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    LocalMux I__8175 (
            .O(N__38924),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ));
    CascadeMux I__8174 (
            .O(N__38919),
            .I(N__38916));
    InMux I__8173 (
            .O(N__38916),
            .I(N__38913));
    LocalMux I__8172 (
            .O(N__38913),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ));
    InMux I__8171 (
            .O(N__38910),
            .I(N__38907));
    LocalMux I__8170 (
            .O(N__38907),
            .I(N__38904));
    Span4Mux_v I__8169 (
            .O(N__38904),
            .I(N__38901));
    Odrv4 I__8168 (
            .O(N__38901),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ));
    InMux I__8167 (
            .O(N__38898),
            .I(N__38894));
    InMux I__8166 (
            .O(N__38897),
            .I(N__38891));
    LocalMux I__8165 (
            .O(N__38894),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    LocalMux I__8164 (
            .O(N__38891),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ));
    CascadeMux I__8163 (
            .O(N__38886),
            .I(N__38883));
    InMux I__8162 (
            .O(N__38883),
            .I(N__38880));
    LocalMux I__8161 (
            .O(N__38880),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ));
    InMux I__8160 (
            .O(N__38877),
            .I(N__38873));
    InMux I__8159 (
            .O(N__38876),
            .I(N__38870));
    LocalMux I__8158 (
            .O(N__38873),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    LocalMux I__8157 (
            .O(N__38870),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ));
    CascadeMux I__8156 (
            .O(N__38865),
            .I(N__38862));
    InMux I__8155 (
            .O(N__38862),
            .I(N__38859));
    LocalMux I__8154 (
            .O(N__38859),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ));
    CascadeMux I__8153 (
            .O(N__38856),
            .I(N__38852));
    CascadeMux I__8152 (
            .O(N__38855),
            .I(N__38849));
    InMux I__8151 (
            .O(N__38852),
            .I(N__38846));
    InMux I__8150 (
            .O(N__38849),
            .I(N__38841));
    LocalMux I__8149 (
            .O(N__38846),
            .I(N__38838));
    CascadeMux I__8148 (
            .O(N__38845),
            .I(N__38835));
    InMux I__8147 (
            .O(N__38844),
            .I(N__38829));
    LocalMux I__8146 (
            .O(N__38841),
            .I(N__38824));
    Span4Mux_v I__8145 (
            .O(N__38838),
            .I(N__38824));
    InMux I__8144 (
            .O(N__38835),
            .I(N__38821));
    InMux I__8143 (
            .O(N__38834),
            .I(N__38817));
    InMux I__8142 (
            .O(N__38833),
            .I(N__38814));
    InMux I__8141 (
            .O(N__38832),
            .I(N__38811));
    LocalMux I__8140 (
            .O(N__38829),
            .I(N__38808));
    Sp12to4 I__8139 (
            .O(N__38824),
            .I(N__38803));
    LocalMux I__8138 (
            .O(N__38821),
            .I(N__38803));
    InMux I__8137 (
            .O(N__38820),
            .I(N__38800));
    LocalMux I__8136 (
            .O(N__38817),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__8135 (
            .O(N__38814),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__8134 (
            .O(N__38811),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv4 I__8133 (
            .O(N__38808),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    Odrv12 I__8132 (
            .O(N__38803),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    LocalMux I__8131 (
            .O(N__38800),
            .I(\phase_controller_inst1.stateZ0Z_3 ));
    InMux I__8130 (
            .O(N__38787),
            .I(N__38783));
    InMux I__8129 (
            .O(N__38786),
            .I(N__38780));
    LocalMux I__8128 (
            .O(N__38783),
            .I(\phase_controller_inst1.stoper_hc.N_8_0 ));
    LocalMux I__8127 (
            .O(N__38780),
            .I(\phase_controller_inst1.stoper_hc.N_8_0 ));
    InMux I__8126 (
            .O(N__38775),
            .I(N__38767));
    InMux I__8125 (
            .O(N__38774),
            .I(N__38764));
    InMux I__8124 (
            .O(N__38773),
            .I(N__38761));
    InMux I__8123 (
            .O(N__38772),
            .I(N__38754));
    InMux I__8122 (
            .O(N__38771),
            .I(N__38754));
    InMux I__8121 (
            .O(N__38770),
            .I(N__38754));
    LocalMux I__8120 (
            .O(N__38767),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__8119 (
            .O(N__38764),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__8118 (
            .O(N__38761),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__8117 (
            .O(N__38754),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    IoInMux I__8116 (
            .O(N__38745),
            .I(N__38742));
    LocalMux I__8115 (
            .O(N__38742),
            .I(N__38739));
    IoSpan4Mux I__8114 (
            .O(N__38739),
            .I(N__38736));
    Span4Mux_s2_v I__8113 (
            .O(N__38736),
            .I(N__38733));
    Sp12to4 I__8112 (
            .O(N__38733),
            .I(N__38730));
    Span12Mux_v I__8111 (
            .O(N__38730),
            .I(N__38727));
    Span12Mux_v I__8110 (
            .O(N__38727),
            .I(N__38723));
    InMux I__8109 (
            .O(N__38726),
            .I(N__38720));
    Odrv12 I__8108 (
            .O(N__38723),
            .I(test22_c));
    LocalMux I__8107 (
            .O(N__38720),
            .I(test22_c));
    InMux I__8106 (
            .O(N__38715),
            .I(N__38711));
    InMux I__8105 (
            .O(N__38714),
            .I(N__38708));
    LocalMux I__8104 (
            .O(N__38711),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__8103 (
            .O(N__38708),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    InMux I__8102 (
            .O(N__38703),
            .I(N__38699));
    InMux I__8101 (
            .O(N__38702),
            .I(N__38696));
    LocalMux I__8100 (
            .O(N__38699),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    LocalMux I__8099 (
            .O(N__38696),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    CascadeMux I__8098 (
            .O(N__38691),
            .I(N__38688));
    InMux I__8097 (
            .O(N__38688),
            .I(N__38685));
    LocalMux I__8096 (
            .O(N__38685),
            .I(N__38682));
    Odrv4 I__8095 (
            .O(N__38682),
            .I(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ));
    InMux I__8094 (
            .O(N__38679),
            .I(N__38675));
    InMux I__8093 (
            .O(N__38678),
            .I(N__38671));
    LocalMux I__8092 (
            .O(N__38675),
            .I(N__38668));
    InMux I__8091 (
            .O(N__38674),
            .I(N__38665));
    LocalMux I__8090 (
            .O(N__38671),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv12 I__8089 (
            .O(N__38668),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    LocalMux I__8088 (
            .O(N__38665),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    IoInMux I__8087 (
            .O(N__38658),
            .I(N__38655));
    LocalMux I__8086 (
            .O(N__38655),
            .I(N__38652));
    Span4Mux_s3_v I__8085 (
            .O(N__38652),
            .I(N__38649));
    Span4Mux_v I__8084 (
            .O(N__38649),
            .I(N__38646));
    Span4Mux_v I__8083 (
            .O(N__38646),
            .I(N__38643));
    Odrv4 I__8082 (
            .O(N__38643),
            .I(\current_shift_inst.timer_s1.N_339_i ));
    CascadeMux I__8081 (
            .O(N__38640),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ));
    InMux I__8080 (
            .O(N__38637),
            .I(N__38634));
    LocalMux I__8079 (
            .O(N__38634),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ));
    CascadeMux I__8078 (
            .O(N__38631),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ));
    InMux I__8077 (
            .O(N__38628),
            .I(N__38625));
    LocalMux I__8076 (
            .O(N__38625),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ));
    InMux I__8075 (
            .O(N__38622),
            .I(N__38619));
    LocalMux I__8074 (
            .O(N__38619),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ));
    CascadeMux I__8073 (
            .O(N__38616),
            .I(N__38613));
    InMux I__8072 (
            .O(N__38613),
            .I(N__38609));
    InMux I__8071 (
            .O(N__38612),
            .I(N__38606));
    LocalMux I__8070 (
            .O(N__38609),
            .I(N__38603));
    LocalMux I__8069 (
            .O(N__38606),
            .I(N__38599));
    Span4Mux_v I__8068 (
            .O(N__38603),
            .I(N__38596));
    InMux I__8067 (
            .O(N__38602),
            .I(N__38593));
    Span4Mux_v I__8066 (
            .O(N__38599),
            .I(N__38589));
    Span4Mux_h I__8065 (
            .O(N__38596),
            .I(N__38586));
    LocalMux I__8064 (
            .O(N__38593),
            .I(N__38583));
    InMux I__8063 (
            .O(N__38592),
            .I(N__38580));
    Odrv4 I__8062 (
            .O(N__38589),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__8061 (
            .O(N__38586),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__8060 (
            .O(N__38583),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    LocalMux I__8059 (
            .O(N__38580),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    InMux I__8058 (
            .O(N__38571),
            .I(N__38566));
    InMux I__8057 (
            .O(N__38570),
            .I(N__38563));
    InMux I__8056 (
            .O(N__38569),
            .I(N__38560));
    LocalMux I__8055 (
            .O(N__38566),
            .I(N__38555));
    LocalMux I__8054 (
            .O(N__38563),
            .I(N__38555));
    LocalMux I__8053 (
            .O(N__38560),
            .I(N__38552));
    Span4Mux_h I__8052 (
            .O(N__38555),
            .I(N__38547));
    Span4Mux_h I__8051 (
            .O(N__38552),
            .I(N__38547));
    Odrv4 I__8050 (
            .O(N__38547),
            .I(\current_shift_inst.un4_control_input1_8 ));
    CascadeMux I__8049 (
            .O(N__38544),
            .I(N__38541));
    InMux I__8048 (
            .O(N__38541),
            .I(N__38538));
    LocalMux I__8047 (
            .O(N__38538),
            .I(N__38535));
    Odrv12 I__8046 (
            .O(N__38535),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    InMux I__8045 (
            .O(N__38532),
            .I(N__38510));
    InMux I__8044 (
            .O(N__38531),
            .I(N__38510));
    InMux I__8043 (
            .O(N__38530),
            .I(N__38510));
    InMux I__8042 (
            .O(N__38529),
            .I(N__38501));
    InMux I__8041 (
            .O(N__38528),
            .I(N__38501));
    InMux I__8040 (
            .O(N__38527),
            .I(N__38501));
    InMux I__8039 (
            .O(N__38526),
            .I(N__38501));
    InMux I__8038 (
            .O(N__38525),
            .I(N__38494));
    InMux I__8037 (
            .O(N__38524),
            .I(N__38491));
    InMux I__8036 (
            .O(N__38523),
            .I(N__38486));
    InMux I__8035 (
            .O(N__38522),
            .I(N__38486));
    InMux I__8034 (
            .O(N__38521),
            .I(N__38483));
    InMux I__8033 (
            .O(N__38520),
            .I(N__38478));
    InMux I__8032 (
            .O(N__38519),
            .I(N__38478));
    InMux I__8031 (
            .O(N__38518),
            .I(N__38475));
    InMux I__8030 (
            .O(N__38517),
            .I(N__38472));
    LocalMux I__8029 (
            .O(N__38510),
            .I(N__38467));
    LocalMux I__8028 (
            .O(N__38501),
            .I(N__38467));
    InMux I__8027 (
            .O(N__38500),
            .I(N__38462));
    InMux I__8026 (
            .O(N__38499),
            .I(N__38462));
    InMux I__8025 (
            .O(N__38498),
            .I(N__38457));
    InMux I__8024 (
            .O(N__38497),
            .I(N__38457));
    LocalMux I__8023 (
            .O(N__38494),
            .I(N__38452));
    LocalMux I__8022 (
            .O(N__38491),
            .I(N__38452));
    LocalMux I__8021 (
            .O(N__38486),
            .I(N__38449));
    LocalMux I__8020 (
            .O(N__38483),
            .I(N__38440));
    LocalMux I__8019 (
            .O(N__38478),
            .I(N__38440));
    LocalMux I__8018 (
            .O(N__38475),
            .I(N__38440));
    LocalMux I__8017 (
            .O(N__38472),
            .I(N__38433));
    Span4Mux_v I__8016 (
            .O(N__38467),
            .I(N__38433));
    LocalMux I__8015 (
            .O(N__38462),
            .I(N__38433));
    LocalMux I__8014 (
            .O(N__38457),
            .I(N__38423));
    Span4Mux_v I__8013 (
            .O(N__38452),
            .I(N__38423));
    Span4Mux_v I__8012 (
            .O(N__38449),
            .I(N__38423));
    InMux I__8011 (
            .O(N__38448),
            .I(N__38418));
    InMux I__8010 (
            .O(N__38447),
            .I(N__38418));
    Span4Mux_v I__8009 (
            .O(N__38440),
            .I(N__38413));
    Span4Mux_v I__8008 (
            .O(N__38433),
            .I(N__38413));
    InMux I__8007 (
            .O(N__38432),
            .I(N__38410));
    InMux I__8006 (
            .O(N__38431),
            .I(N__38405));
    InMux I__8005 (
            .O(N__38430),
            .I(N__38405));
    Odrv4 I__8004 (
            .O(N__38423),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8003 (
            .O(N__38418),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__8002 (
            .O(N__38413),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8001 (
            .O(N__38410),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8000 (
            .O(N__38405),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__7999 (
            .O(N__38394),
            .I(N__38391));
    InMux I__7998 (
            .O(N__38391),
            .I(N__38388));
    LocalMux I__7997 (
            .O(N__38388),
            .I(N__38384));
    InMux I__7996 (
            .O(N__38387),
            .I(N__38381));
    Span4Mux_h I__7995 (
            .O(N__38384),
            .I(N__38378));
    LocalMux I__7994 (
            .O(N__38381),
            .I(N__38373));
    Span4Mux_h I__7993 (
            .O(N__38378),
            .I(N__38370));
    InMux I__7992 (
            .O(N__38377),
            .I(N__38367));
    InMux I__7991 (
            .O(N__38376),
            .I(N__38364));
    Odrv12 I__7990 (
            .O(N__38373),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__7989 (
            .O(N__38370),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__7988 (
            .O(N__38367),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__7987 (
            .O(N__38364),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    CascadeMux I__7986 (
            .O(N__38355),
            .I(N__38352));
    InMux I__7985 (
            .O(N__38352),
            .I(N__38348));
    InMux I__7984 (
            .O(N__38351),
            .I(N__38344));
    LocalMux I__7983 (
            .O(N__38348),
            .I(N__38341));
    InMux I__7982 (
            .O(N__38347),
            .I(N__38338));
    LocalMux I__7981 (
            .O(N__38344),
            .I(N__38335));
    Span4Mux_h I__7980 (
            .O(N__38341),
            .I(N__38332));
    LocalMux I__7979 (
            .O(N__38338),
            .I(N__38329));
    Span4Mux_h I__7978 (
            .O(N__38335),
            .I(N__38326));
    Odrv4 I__7977 (
            .O(N__38332),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv12 I__7976 (
            .O(N__38329),
            .I(\current_shift_inst.un4_control_input1_16 ));
    Odrv4 I__7975 (
            .O(N__38326),
            .I(\current_shift_inst.un4_control_input1_16 ));
    InMux I__7974 (
            .O(N__38319),
            .I(N__38316));
    LocalMux I__7973 (
            .O(N__38316),
            .I(N__38313));
    Span4Mux_v I__7972 (
            .O(N__38313),
            .I(N__38310));
    Span4Mux_h I__7971 (
            .O(N__38310),
            .I(N__38307));
    Odrv4 I__7970 (
            .O(N__38307),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    InMux I__7969 (
            .O(N__38304),
            .I(N__38300));
    InMux I__7968 (
            .O(N__38303),
            .I(N__38297));
    LocalMux I__7967 (
            .O(N__38300),
            .I(N__38291));
    LocalMux I__7966 (
            .O(N__38297),
            .I(N__38291));
    InMux I__7965 (
            .O(N__38296),
            .I(N__38288));
    Span4Mux_v I__7964 (
            .O(N__38291),
            .I(N__38283));
    LocalMux I__7963 (
            .O(N__38288),
            .I(N__38283));
    Odrv4 I__7962 (
            .O(N__38283),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    InMux I__7961 (
            .O(N__38280),
            .I(N__38276));
    InMux I__7960 (
            .O(N__38279),
            .I(N__38273));
    LocalMux I__7959 (
            .O(N__38276),
            .I(N__38266));
    LocalMux I__7958 (
            .O(N__38273),
            .I(N__38266));
    InMux I__7957 (
            .O(N__38272),
            .I(N__38261));
    InMux I__7956 (
            .O(N__38271),
            .I(N__38261));
    Span4Mux_v I__7955 (
            .O(N__38266),
            .I(N__38258));
    LocalMux I__7954 (
            .O(N__38261),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__7953 (
            .O(N__38258),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__7952 (
            .O(N__38253),
            .I(N__38245));
    InMux I__7951 (
            .O(N__38252),
            .I(N__38245));
    InMux I__7950 (
            .O(N__38251),
            .I(N__38242));
    InMux I__7949 (
            .O(N__38250),
            .I(N__38239));
    LocalMux I__7948 (
            .O(N__38245),
            .I(N__38236));
    LocalMux I__7947 (
            .O(N__38242),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    LocalMux I__7946 (
            .O(N__38239),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv12 I__7945 (
            .O(N__38236),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__7944 (
            .O(N__38229),
            .I(N__38226));
    LocalMux I__7943 (
            .O(N__38226),
            .I(N__38223));
    Span4Mux_s3_h I__7942 (
            .O(N__38223),
            .I(N__38219));
    InMux I__7941 (
            .O(N__38222),
            .I(N__38216));
    Sp12to4 I__7940 (
            .O(N__38219),
            .I(N__38213));
    LocalMux I__7939 (
            .O(N__38216),
            .I(N__38210));
    Span12Mux_s11_v I__7938 (
            .O(N__38213),
            .I(N__38207));
    Odrv4 I__7937 (
            .O(N__38210),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv12 I__7936 (
            .O(N__38207),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__7935 (
            .O(N__38202),
            .I(N__38199));
    LocalMux I__7934 (
            .O(N__38199),
            .I(N__38196));
    Span4Mux_v I__7933 (
            .O(N__38196),
            .I(N__38193));
    Sp12to4 I__7932 (
            .O(N__38193),
            .I(N__38190));
    Odrv12 I__7931 (
            .O(N__38190),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__7930 (
            .O(N__38187),
            .I(N__38182));
    InMux I__7929 (
            .O(N__38186),
            .I(N__38179));
    InMux I__7928 (
            .O(N__38185),
            .I(N__38175));
    LocalMux I__7927 (
            .O(N__38182),
            .I(N__38170));
    LocalMux I__7926 (
            .O(N__38179),
            .I(N__38170));
    InMux I__7925 (
            .O(N__38178),
            .I(N__38167));
    LocalMux I__7924 (
            .O(N__38175),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv4 I__7923 (
            .O(N__38170),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    LocalMux I__7922 (
            .O(N__38167),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    CEMux I__7921 (
            .O(N__38160),
            .I(N__38157));
    LocalMux I__7920 (
            .O(N__38157),
            .I(N__38154));
    Span4Mux_v I__7919 (
            .O(N__38154),
            .I(N__38150));
    InMux I__7918 (
            .O(N__38153),
            .I(N__38147));
    Sp12to4 I__7917 (
            .O(N__38150),
            .I(N__38142));
    LocalMux I__7916 (
            .O(N__38147),
            .I(N__38142));
    Span12Mux_v I__7915 (
            .O(N__38142),
            .I(N__38139));
    Odrv12 I__7914 (
            .O(N__38139),
            .I(S1_RNI9RLH));
    CascadeMux I__7913 (
            .O(N__38136),
            .I(\current_shift_inst.PI_CTRL.N_77_cascade_ ));
    InMux I__7912 (
            .O(N__38133),
            .I(N__38130));
    LocalMux I__7911 (
            .O(N__38130),
            .I(N__38127));
    Span4Mux_h I__7910 (
            .O(N__38127),
            .I(N__38124));
    Odrv4 I__7909 (
            .O(N__38124),
            .I(\current_shift_inst.PI_CTRL.N_286 ));
    InMux I__7908 (
            .O(N__38121),
            .I(N__38118));
    LocalMux I__7907 (
            .O(N__38118),
            .I(N__38115));
    Odrv12 I__7906 (
            .O(N__38115),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__7905 (
            .O(N__38112),
            .I(N__38108));
    InMux I__7904 (
            .O(N__38111),
            .I(N__38105));
    LocalMux I__7903 (
            .O(N__38108),
            .I(N__38102));
    LocalMux I__7902 (
            .O(N__38105),
            .I(N__38098));
    Span4Mux_h I__7901 (
            .O(N__38102),
            .I(N__38095));
    InMux I__7900 (
            .O(N__38101),
            .I(N__38092));
    Span4Mux_v I__7899 (
            .O(N__38098),
            .I(N__38085));
    Span4Mux_v I__7898 (
            .O(N__38095),
            .I(N__38085));
    LocalMux I__7897 (
            .O(N__38092),
            .I(N__38085));
    Span4Mux_h I__7896 (
            .O(N__38085),
            .I(N__38081));
    InMux I__7895 (
            .O(N__38084),
            .I(N__38078));
    Odrv4 I__7894 (
            .O(N__38081),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__7893 (
            .O(N__38078),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    InMux I__7892 (
            .O(N__38073),
            .I(N__38070));
    LocalMux I__7891 (
            .O(N__38070),
            .I(N__38067));
    Odrv4 I__7890 (
            .O(N__38067),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__7889 (
            .O(N__38064),
            .I(N__38061));
    LocalMux I__7888 (
            .O(N__38061),
            .I(N__38057));
    InMux I__7887 (
            .O(N__38060),
            .I(N__38054));
    Span4Mux_h I__7886 (
            .O(N__38057),
            .I(N__38049));
    LocalMux I__7885 (
            .O(N__38054),
            .I(N__38049));
    Span4Mux_h I__7884 (
            .O(N__38049),
            .I(N__38044));
    InMux I__7883 (
            .O(N__38048),
            .I(N__38041));
    InMux I__7882 (
            .O(N__38047),
            .I(N__38038));
    Odrv4 I__7881 (
            .O(N__38044),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__7880 (
            .O(N__38041),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__7879 (
            .O(N__38038),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__7878 (
            .O(N__38031),
            .I(N__38026));
    InMux I__7877 (
            .O(N__38030),
            .I(N__38023));
    InMux I__7876 (
            .O(N__38029),
            .I(N__38020));
    LocalMux I__7875 (
            .O(N__38026),
            .I(N__38017));
    LocalMux I__7874 (
            .O(N__38023),
            .I(N__38014));
    LocalMux I__7873 (
            .O(N__38020),
            .I(N__38011));
    Span4Mux_v I__7872 (
            .O(N__38017),
            .I(N__38008));
    Span4Mux_h I__7871 (
            .O(N__38014),
            .I(N__38005));
    Span4Mux_h I__7870 (
            .O(N__38011),
            .I(N__38002));
    Odrv4 I__7869 (
            .O(N__38008),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__7868 (
            .O(N__38005),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv4 I__7867 (
            .O(N__38002),
            .I(\current_shift_inst.un4_control_input1_12 ));
    InMux I__7866 (
            .O(N__37995),
            .I(N__37992));
    LocalMux I__7865 (
            .O(N__37992),
            .I(N__37989));
    Span4Mux_v I__7864 (
            .O(N__37989),
            .I(N__37986));
    Odrv4 I__7863 (
            .O(N__37986),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__7862 (
            .O(N__37983),
            .I(N__37979));
    InMux I__7861 (
            .O(N__37982),
            .I(N__37976));
    InMux I__7860 (
            .O(N__37979),
            .I(N__37973));
    LocalMux I__7859 (
            .O(N__37976),
            .I(N__37970));
    LocalMux I__7858 (
            .O(N__37973),
            .I(N__37967));
    Span4Mux_v I__7857 (
            .O(N__37970),
            .I(N__37962));
    Span4Mux_h I__7856 (
            .O(N__37967),
            .I(N__37962));
    Span4Mux_h I__7855 (
            .O(N__37962),
            .I(N__37957));
    InMux I__7854 (
            .O(N__37961),
            .I(N__37954));
    InMux I__7853 (
            .O(N__37960),
            .I(N__37951));
    Odrv4 I__7852 (
            .O(N__37957),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__7851 (
            .O(N__37954),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__7850 (
            .O(N__37951),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__7849 (
            .O(N__37944),
            .I(N__37941));
    LocalMux I__7848 (
            .O(N__37941),
            .I(N__37937));
    InMux I__7847 (
            .O(N__37940),
            .I(N__37934));
    Span4Mux_v I__7846 (
            .O(N__37937),
            .I(N__37930));
    LocalMux I__7845 (
            .O(N__37934),
            .I(N__37927));
    InMux I__7844 (
            .O(N__37933),
            .I(N__37924));
    Span4Mux_h I__7843 (
            .O(N__37930),
            .I(N__37921));
    Span4Mux_h I__7842 (
            .O(N__37927),
            .I(N__37918));
    LocalMux I__7841 (
            .O(N__37924),
            .I(N__37915));
    Odrv4 I__7840 (
            .O(N__37921),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__7839 (
            .O(N__37918),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__7838 (
            .O(N__37915),
            .I(\current_shift_inst.un4_control_input1_18 ));
    CascadeMux I__7837 (
            .O(N__37908),
            .I(N__37905));
    InMux I__7836 (
            .O(N__37905),
            .I(N__37902));
    LocalMux I__7835 (
            .O(N__37902),
            .I(N__37899));
    Span4Mux_h I__7834 (
            .O(N__37899),
            .I(N__37896));
    Odrv4 I__7833 (
            .O(N__37896),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__7832 (
            .O(N__37893),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__7831 (
            .O(N__37890),
            .I(N__37884));
    InMux I__7830 (
            .O(N__37889),
            .I(N__37884));
    LocalMux I__7829 (
            .O(N__37884),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ));
    InMux I__7828 (
            .O(N__37881),
            .I(N__37874));
    InMux I__7827 (
            .O(N__37880),
            .I(N__37874));
    InMux I__7826 (
            .O(N__37879),
            .I(N__37871));
    LocalMux I__7825 (
            .O(N__37874),
            .I(N__37868));
    LocalMux I__7824 (
            .O(N__37871),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    Odrv4 I__7823 (
            .O(N__37868),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ));
    CascadeMux I__7822 (
            .O(N__37863),
            .I(N__37859));
    InMux I__7821 (
            .O(N__37862),
            .I(N__37853));
    InMux I__7820 (
            .O(N__37859),
            .I(N__37853));
    InMux I__7819 (
            .O(N__37858),
            .I(N__37850));
    LocalMux I__7818 (
            .O(N__37853),
            .I(N__37847));
    LocalMux I__7817 (
            .O(N__37850),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    Odrv4 I__7816 (
            .O(N__37847),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ));
    CascadeMux I__7815 (
            .O(N__37842),
            .I(N__37838));
    InMux I__7814 (
            .O(N__37841),
            .I(N__37833));
    InMux I__7813 (
            .O(N__37838),
            .I(N__37833));
    LocalMux I__7812 (
            .O(N__37833),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ));
    CascadeMux I__7811 (
            .O(N__37830),
            .I(N__37827));
    InMux I__7810 (
            .O(N__37827),
            .I(N__37823));
    CascadeMux I__7809 (
            .O(N__37826),
            .I(N__37820));
    LocalMux I__7808 (
            .O(N__37823),
            .I(N__37817));
    InMux I__7807 (
            .O(N__37820),
            .I(N__37814));
    Span4Mux_h I__7806 (
            .O(N__37817),
            .I(N__37811));
    LocalMux I__7805 (
            .O(N__37814),
            .I(N__37808));
    Odrv4 I__7804 (
            .O(N__37811),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    Odrv4 I__7803 (
            .O(N__37808),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ));
    InMux I__7802 (
            .O(N__37803),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ));
    InMux I__7801 (
            .O(N__37800),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ));
    InMux I__7800 (
            .O(N__37797),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ));
    InMux I__7799 (
            .O(N__37794),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ));
    InMux I__7798 (
            .O(N__37791),
            .I(N__37786));
    InMux I__7797 (
            .O(N__37790),
            .I(N__37781));
    InMux I__7796 (
            .O(N__37789),
            .I(N__37781));
    LocalMux I__7795 (
            .O(N__37786),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    LocalMux I__7794 (
            .O(N__37781),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ));
    CascadeMux I__7793 (
            .O(N__37776),
            .I(N__37771));
    InMux I__7792 (
            .O(N__37775),
            .I(N__37768));
    InMux I__7791 (
            .O(N__37774),
            .I(N__37763));
    InMux I__7790 (
            .O(N__37771),
            .I(N__37763));
    LocalMux I__7789 (
            .O(N__37768),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    LocalMux I__7788 (
            .O(N__37763),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ));
    CascadeMux I__7787 (
            .O(N__37758),
            .I(N__37755));
    InMux I__7786 (
            .O(N__37755),
            .I(N__37749));
    InMux I__7785 (
            .O(N__37754),
            .I(N__37749));
    LocalMux I__7784 (
            .O(N__37749),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ));
    InMux I__7783 (
            .O(N__37746),
            .I(N__37740));
    InMux I__7782 (
            .O(N__37745),
            .I(N__37740));
    LocalMux I__7781 (
            .O(N__37740),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ));
    InMux I__7780 (
            .O(N__37737),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ));
    InMux I__7779 (
            .O(N__37734),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ));
    InMux I__7778 (
            .O(N__37731),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ));
    InMux I__7777 (
            .O(N__37728),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ));
    InMux I__7776 (
            .O(N__37725),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ));
    InMux I__7775 (
            .O(N__37722),
            .I(N__37717));
    InMux I__7774 (
            .O(N__37721),
            .I(N__37714));
    InMux I__7773 (
            .O(N__37720),
            .I(N__37711));
    LocalMux I__7772 (
            .O(N__37717),
            .I(N__37708));
    LocalMux I__7771 (
            .O(N__37714),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    LocalMux I__7770 (
            .O(N__37711),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    Odrv4 I__7769 (
            .O(N__37708),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ));
    InMux I__7768 (
            .O(N__37701),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ));
    InMux I__7767 (
            .O(N__37698),
            .I(N__37693));
    InMux I__7766 (
            .O(N__37697),
            .I(N__37690));
    InMux I__7765 (
            .O(N__37696),
            .I(N__37687));
    LocalMux I__7764 (
            .O(N__37693),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__7763 (
            .O(N__37690),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    LocalMux I__7762 (
            .O(N__37687),
            .I(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ));
    InMux I__7761 (
            .O(N__37680),
            .I(bfn_15_8_0_));
    InMux I__7760 (
            .O(N__37677),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ));
    InMux I__7759 (
            .O(N__37674),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ));
    InMux I__7758 (
            .O(N__37671),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ));
    InMux I__7757 (
            .O(N__37668),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ));
    InMux I__7756 (
            .O(N__37665),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ));
    InMux I__7755 (
            .O(N__37662),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ));
    InMux I__7754 (
            .O(N__37659),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ));
    InMux I__7753 (
            .O(N__37656),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ));
    InMux I__7752 (
            .O(N__37653),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ));
    InMux I__7751 (
            .O(N__37650),
            .I(bfn_15_7_0_));
    InMux I__7750 (
            .O(N__37647),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ));
    InMux I__7749 (
            .O(N__37644),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ));
    CascadeMux I__7748 (
            .O(N__37641),
            .I(N__37637));
    CascadeMux I__7747 (
            .O(N__37640),
            .I(N__37634));
    InMux I__7746 (
            .O(N__37637),
            .I(N__37629));
    InMux I__7745 (
            .O(N__37634),
            .I(N__37629));
    LocalMux I__7744 (
            .O(N__37629),
            .I(\phase_controller_inst1.stoper_hc.N_45_i ));
    InMux I__7743 (
            .O(N__37626),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ));
    InMux I__7742 (
            .O(N__37623),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ));
    InMux I__7741 (
            .O(N__37620),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ));
    InMux I__7740 (
            .O(N__37617),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ));
    InMux I__7739 (
            .O(N__37614),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ));
    InMux I__7738 (
            .O(N__37611),
            .I(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ));
    InMux I__7737 (
            .O(N__37608),
            .I(bfn_15_6_0_));
    InMux I__7736 (
            .O(N__37605),
            .I(N__37602));
    LocalMux I__7735 (
            .O(N__37602),
            .I(\phase_controller_inst1.stoper_hc.N_27 ));
    InMux I__7734 (
            .O(N__37599),
            .I(N__37596));
    LocalMux I__7733 (
            .O(N__37596),
            .I(N__37593));
    Span4Mux_h I__7732 (
            .O(N__37593),
            .I(N__37590));
    Span4Mux_h I__7731 (
            .O(N__37590),
            .I(N__37587));
    Odrv4 I__7730 (
            .O(N__37587),
            .I(il_max_comp1_c));
    InMux I__7729 (
            .O(N__37584),
            .I(N__37581));
    LocalMux I__7728 (
            .O(N__37581),
            .I(N__37576));
    InMux I__7727 (
            .O(N__37580),
            .I(N__37569));
    InMux I__7726 (
            .O(N__37579),
            .I(N__37569));
    Span4Mux_h I__7725 (
            .O(N__37576),
            .I(N__37566));
    InMux I__7724 (
            .O(N__37575),
            .I(N__37563));
    InMux I__7723 (
            .O(N__37574),
            .I(N__37560));
    LocalMux I__7722 (
            .O(N__37569),
            .I(\phase_controller_inst1.N_175_1 ));
    Odrv4 I__7721 (
            .O(N__37566),
            .I(\phase_controller_inst1.N_175_1 ));
    LocalMux I__7720 (
            .O(N__37563),
            .I(\phase_controller_inst1.N_175_1 ));
    LocalMux I__7719 (
            .O(N__37560),
            .I(\phase_controller_inst1.N_175_1 ));
    CascadeMux I__7718 (
            .O(N__37551),
            .I(\phase_controller_inst1.stoper_hc.N_8_0_cascade_ ));
    InMux I__7717 (
            .O(N__37548),
            .I(N__37545));
    LocalMux I__7716 (
            .O(N__37545),
            .I(\phase_controller_inst1.stoper_hc.m12_ns_1 ));
    InMux I__7715 (
            .O(N__37542),
            .I(N__37535));
    InMux I__7714 (
            .O(N__37541),
            .I(N__37535));
    InMux I__7713 (
            .O(N__37540),
            .I(N__37530));
    LocalMux I__7712 (
            .O(N__37535),
            .I(N__37527));
    InMux I__7711 (
            .O(N__37534),
            .I(N__37524));
    InMux I__7710 (
            .O(N__37533),
            .I(N__37521));
    LocalMux I__7709 (
            .O(N__37530),
            .I(N__37518));
    Span4Mux_h I__7708 (
            .O(N__37527),
            .I(N__37515));
    LocalMux I__7707 (
            .O(N__37524),
            .I(N__37510));
    LocalMux I__7706 (
            .O(N__37521),
            .I(N__37510));
    Span12Mux_h I__7705 (
            .O(N__37518),
            .I(N__37507));
    IoSpan4Mux I__7704 (
            .O(N__37515),
            .I(N__37502));
    IoSpan4Mux I__7703 (
            .O(N__37510),
            .I(N__37502));
    Odrv12 I__7702 (
            .O(N__37507),
            .I(il_min_comp1_c));
    Odrv4 I__7701 (
            .O(N__37502),
            .I(il_min_comp1_c));
    InMux I__7700 (
            .O(N__37497),
            .I(N__37494));
    LocalMux I__7699 (
            .O(N__37494),
            .I(\phase_controller_inst1.N_14_0 ));
    CascadeMux I__7698 (
            .O(N__37491),
            .I(N__37488));
    InMux I__7697 (
            .O(N__37488),
            .I(N__37485));
    LocalMux I__7696 (
            .O(N__37485),
            .I(N__37482));
    Odrv4 I__7695 (
            .O(N__37482),
            .I(\phase_controller_inst1.N_13_0 ));
    InMux I__7694 (
            .O(N__37479),
            .I(N__37476));
    LocalMux I__7693 (
            .O(N__37476),
            .I(N__37473));
    Span4Mux_v I__7692 (
            .O(N__37473),
            .I(N__37467));
    InMux I__7691 (
            .O(N__37472),
            .I(N__37464));
    CascadeMux I__7690 (
            .O(N__37471),
            .I(N__37459));
    InMux I__7689 (
            .O(N__37470),
            .I(N__37456));
    Sp12to4 I__7688 (
            .O(N__37467),
            .I(N__37453));
    LocalMux I__7687 (
            .O(N__37464),
            .I(N__37450));
    InMux I__7686 (
            .O(N__37463),
            .I(N__37447));
    InMux I__7685 (
            .O(N__37462),
            .I(N__37442));
    InMux I__7684 (
            .O(N__37459),
            .I(N__37442));
    LocalMux I__7683 (
            .O(N__37456),
            .I(N__37437));
    Span12Mux_v I__7682 (
            .O(N__37453),
            .I(N__37437));
    Span4Mux_h I__7681 (
            .O(N__37450),
            .I(N__37434));
    LocalMux I__7680 (
            .O(N__37447),
            .I(N__37431));
    LocalMux I__7679 (
            .O(N__37442),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv12 I__7678 (
            .O(N__37437),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__7677 (
            .O(N__37434),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__7676 (
            .O(N__37431),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    InMux I__7675 (
            .O(N__37422),
            .I(N__37419));
    LocalMux I__7674 (
            .O(N__37419),
            .I(\phase_controller_inst2.m21 ));
    InMux I__7673 (
            .O(N__37416),
            .I(N__37412));
    CascadeMux I__7672 (
            .O(N__37415),
            .I(N__37409));
    LocalMux I__7671 (
            .O(N__37412),
            .I(N__37406));
    InMux I__7670 (
            .O(N__37409),
            .I(N__37403));
    Sp12to4 I__7669 (
            .O(N__37406),
            .I(N__37398));
    LocalMux I__7668 (
            .O(N__37403),
            .I(N__37395));
    InMux I__7667 (
            .O(N__37402),
            .I(N__37392));
    CascadeMux I__7666 (
            .O(N__37401),
            .I(N__37389));
    Span12Mux_s8_v I__7665 (
            .O(N__37398),
            .I(N__37384));
    Span4Mux_v I__7664 (
            .O(N__37395),
            .I(N__37379));
    LocalMux I__7663 (
            .O(N__37392),
            .I(N__37379));
    InMux I__7662 (
            .O(N__37389),
            .I(N__37376));
    InMux I__7661 (
            .O(N__37388),
            .I(N__37373));
    InMux I__7660 (
            .O(N__37387),
            .I(N__37370));
    Span12Mux_v I__7659 (
            .O(N__37384),
            .I(N__37367));
    Span4Mux_h I__7658 (
            .O(N__37379),
            .I(N__37364));
    LocalMux I__7657 (
            .O(N__37376),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__7656 (
            .O(N__37373),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__7655 (
            .O(N__37370),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv12 I__7654 (
            .O(N__37367),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    Odrv4 I__7653 (
            .O(N__37364),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    InMux I__7652 (
            .O(N__37353),
            .I(N__37350));
    LocalMux I__7651 (
            .O(N__37350),
            .I(\phase_controller_inst2.time_passed_er_RNI23UO1 ));
    IoInMux I__7650 (
            .O(N__37347),
            .I(N__37344));
    LocalMux I__7649 (
            .O(N__37344),
            .I(N__37341));
    Span4Mux_s2_v I__7648 (
            .O(N__37341),
            .I(N__37338));
    Sp12to4 I__7647 (
            .O(N__37338),
            .I(N__37335));
    Span12Mux_h I__7646 (
            .O(N__37335),
            .I(N__37332));
    Span12Mux_v I__7645 (
            .O(N__37332),
            .I(N__37329));
    Span12Mux_v I__7644 (
            .O(N__37329),
            .I(N__37325));
    InMux I__7643 (
            .O(N__37328),
            .I(N__37322));
    Odrv12 I__7642 (
            .O(N__37325),
            .I(s1_phy_c));
    LocalMux I__7641 (
            .O(N__37322),
            .I(s1_phy_c));
    InMux I__7640 (
            .O(N__37317),
            .I(N__37313));
    InMux I__7639 (
            .O(N__37316),
            .I(N__37310));
    LocalMux I__7638 (
            .O(N__37313),
            .I(N__37307));
    LocalMux I__7637 (
            .O(N__37310),
            .I(N__37304));
    Span4Mux_v I__7636 (
            .O(N__37307),
            .I(N__37301));
    Span4Mux_h I__7635 (
            .O(N__37304),
            .I(N__37298));
    Sp12to4 I__7634 (
            .O(N__37301),
            .I(N__37295));
    Span4Mux_h I__7633 (
            .O(N__37298),
            .I(N__37292));
    Span12Mux_h I__7632 (
            .O(N__37295),
            .I(N__37289));
    Odrv4 I__7631 (
            .O(N__37292),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    Odrv12 I__7630 (
            .O(N__37289),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__7629 (
            .O(N__37284),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__7628 (
            .O(N__37281),
            .I(N__37278));
    LocalMux I__7627 (
            .O(N__37278),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__7626 (
            .O(N__37275),
            .I(N__37271));
    InMux I__7625 (
            .O(N__37274),
            .I(N__37268));
    LocalMux I__7624 (
            .O(N__37271),
            .I(N__37265));
    LocalMux I__7623 (
            .O(N__37268),
            .I(N__37262));
    Span4Mux_v I__7622 (
            .O(N__37265),
            .I(N__37259));
    Span4Mux_s3_h I__7621 (
            .O(N__37262),
            .I(N__37256));
    Sp12to4 I__7620 (
            .O(N__37259),
            .I(N__37253));
    Span4Mux_h I__7619 (
            .O(N__37256),
            .I(N__37250));
    Span12Mux_s7_h I__7618 (
            .O(N__37253),
            .I(N__37245));
    Sp12to4 I__7617 (
            .O(N__37250),
            .I(N__37245));
    Span12Mux_v I__7616 (
            .O(N__37245),
            .I(N__37242));
    Odrv12 I__7615 (
            .O(N__37242),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__7614 (
            .O(N__37239),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__7613 (
            .O(N__37236),
            .I(N__37233));
    LocalMux I__7612 (
            .O(N__37233),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__7611 (
            .O(N__37230),
            .I(N__37227));
    LocalMux I__7610 (
            .O(N__37227),
            .I(N__37223));
    InMux I__7609 (
            .O(N__37226),
            .I(N__37220));
    Span4Mux_v I__7608 (
            .O(N__37223),
            .I(N__37217));
    LocalMux I__7607 (
            .O(N__37220),
            .I(N__37214));
    Sp12to4 I__7606 (
            .O(N__37217),
            .I(N__37211));
    Span4Mux_v I__7605 (
            .O(N__37214),
            .I(N__37208));
    Span12Mux_s6_h I__7604 (
            .O(N__37211),
            .I(N__37205));
    Sp12to4 I__7603 (
            .O(N__37208),
            .I(N__37200));
    Span12Mux_v I__7602 (
            .O(N__37205),
            .I(N__37200));
    Odrv12 I__7601 (
            .O(N__37200),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__7600 (
            .O(N__37197),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__7599 (
            .O(N__37194),
            .I(N__37191));
    LocalMux I__7598 (
            .O(N__37191),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__7597 (
            .O(N__37188),
            .I(N__37185));
    LocalMux I__7596 (
            .O(N__37185),
            .I(N__37181));
    InMux I__7595 (
            .O(N__37184),
            .I(N__37178));
    Sp12to4 I__7594 (
            .O(N__37181),
            .I(N__37175));
    LocalMux I__7593 (
            .O(N__37178),
            .I(N__37172));
    Span12Mux_v I__7592 (
            .O(N__37175),
            .I(N__37169));
    Span12Mux_v I__7591 (
            .O(N__37172),
            .I(N__37166));
    Span12Mux_h I__7590 (
            .O(N__37169),
            .I(N__37163));
    Odrv12 I__7589 (
            .O(N__37166),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    Odrv12 I__7588 (
            .O(N__37163),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__7587 (
            .O(N__37158),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__7586 (
            .O(N__37155),
            .I(N__37152));
    LocalMux I__7585 (
            .O(N__37152),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    InMux I__7584 (
            .O(N__37149),
            .I(N__37145));
    InMux I__7583 (
            .O(N__37148),
            .I(N__37142));
    LocalMux I__7582 (
            .O(N__37145),
            .I(N__37139));
    LocalMux I__7581 (
            .O(N__37142),
            .I(N__37136));
    Span4Mux_h I__7580 (
            .O(N__37139),
            .I(N__37133));
    Span12Mux_v I__7579 (
            .O(N__37136),
            .I(N__37130));
    Span4Mux_h I__7578 (
            .O(N__37133),
            .I(N__37127));
    Span12Mux_h I__7577 (
            .O(N__37130),
            .I(N__37124));
    Odrv4 I__7576 (
            .O(N__37127),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    Odrv12 I__7575 (
            .O(N__37124),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__7574 (
            .O(N__37119),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__7573 (
            .O(N__37116),
            .I(N__37112));
    InMux I__7572 (
            .O(N__37115),
            .I(N__37109));
    LocalMux I__7571 (
            .O(N__37112),
            .I(\current_shift_inst.control_input_31 ));
    LocalMux I__7570 (
            .O(N__37109),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__7569 (
            .O(N__37104),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__7568 (
            .O(N__37101),
            .I(N__37098));
    LocalMux I__7567 (
            .O(N__37098),
            .I(N__37095));
    Span4Mux_h I__7566 (
            .O(N__37095),
            .I(N__37092));
    Span4Mux_h I__7565 (
            .O(N__37092),
            .I(N__37089));
    Odrv4 I__7564 (
            .O(N__37089),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    IoInMux I__7563 (
            .O(N__37086),
            .I(N__37083));
    LocalMux I__7562 (
            .O(N__37083),
            .I(N__37080));
    Span12Mux_s5_v I__7561 (
            .O(N__37080),
            .I(N__37077));
    Odrv12 I__7560 (
            .O(N__37077),
            .I(s2_phy_c));
    InMux I__7559 (
            .O(N__37074),
            .I(N__37071));
    LocalMux I__7558 (
            .O(N__37071),
            .I(N__37068));
    Odrv4 I__7557 (
            .O(N__37068),
            .I(\phase_controller_inst1.stoper_hc.m19_ns_1 ));
    InMux I__7556 (
            .O(N__37065),
            .I(N__37062));
    LocalMux I__7555 (
            .O(N__37062),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__7554 (
            .O(N__37059),
            .I(N__37056));
    LocalMux I__7553 (
            .O(N__37056),
            .I(N__37053));
    Span4Mux_s2_h I__7552 (
            .O(N__37053),
            .I(N__37049));
    InMux I__7551 (
            .O(N__37052),
            .I(N__37046));
    Sp12to4 I__7550 (
            .O(N__37049),
            .I(N__37043));
    LocalMux I__7549 (
            .O(N__37046),
            .I(N__37038));
    Span12Mux_v I__7548 (
            .O(N__37043),
            .I(N__37038));
    Span12Mux_h I__7547 (
            .O(N__37038),
            .I(N__37035));
    Odrv12 I__7546 (
            .O(N__37035),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__7545 (
            .O(N__37032),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__7544 (
            .O(N__37029),
            .I(N__37026));
    LocalMux I__7543 (
            .O(N__37026),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__7542 (
            .O(N__37023),
            .I(N__37019));
    InMux I__7541 (
            .O(N__37022),
            .I(N__37016));
    LocalMux I__7540 (
            .O(N__37019),
            .I(N__37013));
    LocalMux I__7539 (
            .O(N__37016),
            .I(N__37010));
    Span4Mux_h I__7538 (
            .O(N__37013),
            .I(N__37007));
    Span12Mux_s2_h I__7537 (
            .O(N__37010),
            .I(N__37004));
    Span4Mux_h I__7536 (
            .O(N__37007),
            .I(N__37001));
    Span12Mux_h I__7535 (
            .O(N__37004),
            .I(N__36998));
    Odrv4 I__7534 (
            .O(N__37001),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    Odrv12 I__7533 (
            .O(N__36998),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__7532 (
            .O(N__36993),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__7531 (
            .O(N__36990),
            .I(N__36987));
    LocalMux I__7530 (
            .O(N__36987),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__7529 (
            .O(N__36984),
            .I(N__36980));
    InMux I__7528 (
            .O(N__36983),
            .I(N__36977));
    LocalMux I__7527 (
            .O(N__36980),
            .I(N__36974));
    LocalMux I__7526 (
            .O(N__36977),
            .I(N__36971));
    Sp12to4 I__7525 (
            .O(N__36974),
            .I(N__36968));
    Span4Mux_v I__7524 (
            .O(N__36971),
            .I(N__36965));
    Span12Mux_v I__7523 (
            .O(N__36968),
            .I(N__36962));
    Span4Mux_h I__7522 (
            .O(N__36965),
            .I(N__36959));
    Span12Mux_h I__7521 (
            .O(N__36962),
            .I(N__36956));
    Odrv4 I__7520 (
            .O(N__36959),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv12 I__7519 (
            .O(N__36956),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__7518 (
            .O(N__36951),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__7517 (
            .O(N__36948),
            .I(N__36945));
    LocalMux I__7516 (
            .O(N__36945),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__7515 (
            .O(N__36942),
            .I(N__36939));
    LocalMux I__7514 (
            .O(N__36939),
            .I(N__36935));
    InMux I__7513 (
            .O(N__36938),
            .I(N__36932));
    Span4Mux_v I__7512 (
            .O(N__36935),
            .I(N__36929));
    LocalMux I__7511 (
            .O(N__36932),
            .I(N__36926));
    Sp12to4 I__7510 (
            .O(N__36929),
            .I(N__36921));
    Span12Mux_v I__7509 (
            .O(N__36926),
            .I(N__36921));
    Span12Mux_h I__7508 (
            .O(N__36921),
            .I(N__36918));
    Odrv12 I__7507 (
            .O(N__36918),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    InMux I__7506 (
            .O(N__36915),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__7505 (
            .O(N__36912),
            .I(N__36909));
    LocalMux I__7504 (
            .O(N__36909),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__7503 (
            .O(N__36906),
            .I(N__36903));
    LocalMux I__7502 (
            .O(N__36903),
            .I(N__36900));
    Span4Mux_s3_h I__7501 (
            .O(N__36900),
            .I(N__36896));
    InMux I__7500 (
            .O(N__36899),
            .I(N__36893));
    Span4Mux_v I__7499 (
            .O(N__36896),
            .I(N__36890));
    LocalMux I__7498 (
            .O(N__36893),
            .I(N__36885));
    Span4Mux_v I__7497 (
            .O(N__36890),
            .I(N__36885));
    Sp12to4 I__7496 (
            .O(N__36885),
            .I(N__36882));
    Odrv12 I__7495 (
            .O(N__36882),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__7494 (
            .O(N__36879),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__7493 (
            .O(N__36876),
            .I(N__36873));
    LocalMux I__7492 (
            .O(N__36873),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__7491 (
            .O(N__36870),
            .I(N__36866));
    InMux I__7490 (
            .O(N__36869),
            .I(N__36863));
    LocalMux I__7489 (
            .O(N__36866),
            .I(N__36860));
    LocalMux I__7488 (
            .O(N__36863),
            .I(N__36857));
    Span4Mux_v I__7487 (
            .O(N__36860),
            .I(N__36854));
    Span4Mux_h I__7486 (
            .O(N__36857),
            .I(N__36851));
    Span4Mux_s1_h I__7485 (
            .O(N__36854),
            .I(N__36848));
    Span4Mux_h I__7484 (
            .O(N__36851),
            .I(N__36845));
    Sp12to4 I__7483 (
            .O(N__36848),
            .I(N__36842));
    Span4Mux_h I__7482 (
            .O(N__36845),
            .I(N__36839));
    Span12Mux_h I__7481 (
            .O(N__36842),
            .I(N__36836));
    Odrv4 I__7480 (
            .O(N__36839),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    Odrv12 I__7479 (
            .O(N__36836),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__7478 (
            .O(N__36831),
            .I(bfn_14_21_0_));
    InMux I__7477 (
            .O(N__36828),
            .I(N__36825));
    LocalMux I__7476 (
            .O(N__36825),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__7475 (
            .O(N__36822),
            .I(N__36818));
    InMux I__7474 (
            .O(N__36821),
            .I(N__36815));
    LocalMux I__7473 (
            .O(N__36818),
            .I(N__36812));
    LocalMux I__7472 (
            .O(N__36815),
            .I(N__36809));
    Span4Mux_v I__7471 (
            .O(N__36812),
            .I(N__36806));
    Span4Mux_v I__7470 (
            .O(N__36809),
            .I(N__36803));
    Sp12to4 I__7469 (
            .O(N__36806),
            .I(N__36800));
    Span4Mux_h I__7468 (
            .O(N__36803),
            .I(N__36797));
    Span12Mux_s2_h I__7467 (
            .O(N__36800),
            .I(N__36794));
    Span4Mux_h I__7466 (
            .O(N__36797),
            .I(N__36791));
    Span12Mux_h I__7465 (
            .O(N__36794),
            .I(N__36788));
    Odrv4 I__7464 (
            .O(N__36791),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    Odrv12 I__7463 (
            .O(N__36788),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__7462 (
            .O(N__36783),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__7461 (
            .O(N__36780),
            .I(N__36777));
    LocalMux I__7460 (
            .O(N__36777),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__7459 (
            .O(N__36774),
            .I(N__36771));
    LocalMux I__7458 (
            .O(N__36771),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__7457 (
            .O(N__36768),
            .I(N__36765));
    LocalMux I__7456 (
            .O(N__36765),
            .I(N__36762));
    Span4Mux_v I__7455 (
            .O(N__36762),
            .I(N__36758));
    InMux I__7454 (
            .O(N__36761),
            .I(N__36755));
    Span4Mux_h I__7453 (
            .O(N__36758),
            .I(N__36752));
    LocalMux I__7452 (
            .O(N__36755),
            .I(N__36749));
    Span4Mux_h I__7451 (
            .O(N__36752),
            .I(N__36746));
    Span12Mux_s11_v I__7450 (
            .O(N__36749),
            .I(N__36743));
    Span4Mux_v I__7449 (
            .O(N__36746),
            .I(N__36740));
    Odrv12 I__7448 (
            .O(N__36743),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv4 I__7447 (
            .O(N__36740),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__7446 (
            .O(N__36735),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__7445 (
            .O(N__36732),
            .I(N__36729));
    LocalMux I__7444 (
            .O(N__36729),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__7443 (
            .O(N__36726),
            .I(N__36722));
    InMux I__7442 (
            .O(N__36725),
            .I(N__36719));
    LocalMux I__7441 (
            .O(N__36722),
            .I(N__36716));
    LocalMux I__7440 (
            .O(N__36719),
            .I(N__36713));
    Span4Mux_v I__7439 (
            .O(N__36716),
            .I(N__36710));
    Span4Mux_v I__7438 (
            .O(N__36713),
            .I(N__36707));
    Span4Mux_v I__7437 (
            .O(N__36710),
            .I(N__36704));
    Span4Mux_h I__7436 (
            .O(N__36707),
            .I(N__36701));
    Sp12to4 I__7435 (
            .O(N__36704),
            .I(N__36698));
    Odrv4 I__7434 (
            .O(N__36701),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__7433 (
            .O(N__36698),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__7432 (
            .O(N__36693),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__7431 (
            .O(N__36690),
            .I(N__36687));
    LocalMux I__7430 (
            .O(N__36687),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__7429 (
            .O(N__36684),
            .I(N__36681));
    LocalMux I__7428 (
            .O(N__36681),
            .I(N__36677));
    InMux I__7427 (
            .O(N__36680),
            .I(N__36674));
    Span4Mux_v I__7426 (
            .O(N__36677),
            .I(N__36671));
    LocalMux I__7425 (
            .O(N__36674),
            .I(N__36668));
    Span4Mux_h I__7424 (
            .O(N__36671),
            .I(N__36665));
    Span12Mux_s11_v I__7423 (
            .O(N__36668),
            .I(N__36662));
    Odrv4 I__7422 (
            .O(N__36665),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv12 I__7421 (
            .O(N__36662),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__7420 (
            .O(N__36657),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__7419 (
            .O(N__36654),
            .I(N__36651));
    LocalMux I__7418 (
            .O(N__36651),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__7417 (
            .O(N__36648),
            .I(N__36645));
    LocalMux I__7416 (
            .O(N__36645),
            .I(N__36641));
    InMux I__7415 (
            .O(N__36644),
            .I(N__36638));
    Span4Mux_h I__7414 (
            .O(N__36641),
            .I(N__36635));
    LocalMux I__7413 (
            .O(N__36638),
            .I(N__36632));
    Span4Mux_h I__7412 (
            .O(N__36635),
            .I(N__36629));
    Span12Mux_s11_h I__7411 (
            .O(N__36632),
            .I(N__36626));
    Odrv4 I__7410 (
            .O(N__36629),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv12 I__7409 (
            .O(N__36626),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__7408 (
            .O(N__36621),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__7407 (
            .O(N__36618),
            .I(N__36615));
    LocalMux I__7406 (
            .O(N__36615),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__7405 (
            .O(N__36612),
            .I(N__36609));
    LocalMux I__7404 (
            .O(N__36609),
            .I(N__36606));
    Span4Mux_s3_h I__7403 (
            .O(N__36606),
            .I(N__36602));
    InMux I__7402 (
            .O(N__36605),
            .I(N__36599));
    Sp12to4 I__7401 (
            .O(N__36602),
            .I(N__36596));
    LocalMux I__7400 (
            .O(N__36599),
            .I(N__36591));
    Span12Mux_v I__7399 (
            .O(N__36596),
            .I(N__36591));
    Odrv12 I__7398 (
            .O(N__36591),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__7397 (
            .O(N__36588),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__7396 (
            .O(N__36585),
            .I(N__36582));
    LocalMux I__7395 (
            .O(N__36582),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__7394 (
            .O(N__36579),
            .I(N__36575));
    InMux I__7393 (
            .O(N__36578),
            .I(N__36572));
    LocalMux I__7392 (
            .O(N__36575),
            .I(N__36569));
    LocalMux I__7391 (
            .O(N__36572),
            .I(N__36566));
    Span4Mux_v I__7390 (
            .O(N__36569),
            .I(N__36563));
    Span4Mux_v I__7389 (
            .O(N__36566),
            .I(N__36560));
    Sp12to4 I__7388 (
            .O(N__36563),
            .I(N__36557));
    Span4Mux_h I__7387 (
            .O(N__36560),
            .I(N__36554));
    Span12Mux_s10_h I__7386 (
            .O(N__36557),
            .I(N__36551));
    Span4Mux_h I__7385 (
            .O(N__36554),
            .I(N__36548));
    Span12Mux_v I__7384 (
            .O(N__36551),
            .I(N__36545));
    Odrv4 I__7383 (
            .O(N__36548),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv12 I__7382 (
            .O(N__36545),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__7381 (
            .O(N__36540),
            .I(bfn_14_20_0_));
    InMux I__7380 (
            .O(N__36537),
            .I(N__36534));
    LocalMux I__7379 (
            .O(N__36534),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__7378 (
            .O(N__36531),
            .I(N__36528));
    LocalMux I__7377 (
            .O(N__36528),
            .I(N__36525));
    Span4Mux_s2_h I__7376 (
            .O(N__36525),
            .I(N__36521));
    InMux I__7375 (
            .O(N__36524),
            .I(N__36518));
    Sp12to4 I__7374 (
            .O(N__36521),
            .I(N__36515));
    LocalMux I__7373 (
            .O(N__36518),
            .I(N__36510));
    Span12Mux_v I__7372 (
            .O(N__36515),
            .I(N__36510));
    Span12Mux_h I__7371 (
            .O(N__36510),
            .I(N__36507));
    Odrv12 I__7370 (
            .O(N__36507),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__7369 (
            .O(N__36504),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__7368 (
            .O(N__36501),
            .I(N__36498));
    LocalMux I__7367 (
            .O(N__36498),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__7366 (
            .O(N__36495),
            .I(N__36491));
    InMux I__7365 (
            .O(N__36494),
            .I(N__36488));
    LocalMux I__7364 (
            .O(N__36491),
            .I(N__36485));
    LocalMux I__7363 (
            .O(N__36488),
            .I(N__36482));
    Span4Mux_h I__7362 (
            .O(N__36485),
            .I(N__36479));
    Span4Mux_v I__7361 (
            .O(N__36482),
            .I(N__36476));
    Span4Mux_h I__7360 (
            .O(N__36479),
            .I(N__36473));
    Sp12to4 I__7359 (
            .O(N__36476),
            .I(N__36470));
    Span4Mux_h I__7358 (
            .O(N__36473),
            .I(N__36467));
    Span12Mux_h I__7357 (
            .O(N__36470),
            .I(N__36464));
    Odrv4 I__7356 (
            .O(N__36467),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    Odrv12 I__7355 (
            .O(N__36464),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__7354 (
            .O(N__36459),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__7353 (
            .O(N__36456),
            .I(N__36453));
    LocalMux I__7352 (
            .O(N__36453),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__7351 (
            .O(N__36450),
            .I(N__36447));
    LocalMux I__7350 (
            .O(N__36447),
            .I(N__36444));
    Span4Mux_s2_h I__7349 (
            .O(N__36444),
            .I(N__36440));
    InMux I__7348 (
            .O(N__36443),
            .I(N__36437));
    Span4Mux_h I__7347 (
            .O(N__36440),
            .I(N__36434));
    LocalMux I__7346 (
            .O(N__36437),
            .I(N__36431));
    Span4Mux_h I__7345 (
            .O(N__36434),
            .I(N__36428));
    Span12Mux_v I__7344 (
            .O(N__36431),
            .I(N__36425));
    Span4Mux_v I__7343 (
            .O(N__36428),
            .I(N__36422));
    Odrv12 I__7342 (
            .O(N__36425),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv4 I__7341 (
            .O(N__36422),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__7340 (
            .O(N__36417),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__7339 (
            .O(N__36414),
            .I(N__36411));
    LocalMux I__7338 (
            .O(N__36411),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__7337 (
            .O(N__36408),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__7336 (
            .O(N__36405),
            .I(N__36402));
    LocalMux I__7335 (
            .O(N__36402),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__7334 (
            .O(N__36399),
            .I(N__36396));
    LocalMux I__7333 (
            .O(N__36396),
            .I(N__36392));
    InMux I__7332 (
            .O(N__36395),
            .I(N__36389));
    Span4Mux_h I__7331 (
            .O(N__36392),
            .I(N__36386));
    LocalMux I__7330 (
            .O(N__36389),
            .I(N__36383));
    Span4Mux_h I__7329 (
            .O(N__36386),
            .I(N__36380));
    Span12Mux_v I__7328 (
            .O(N__36383),
            .I(N__36377));
    Odrv4 I__7327 (
            .O(N__36380),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv12 I__7326 (
            .O(N__36377),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__7325 (
            .O(N__36372),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__7324 (
            .O(N__36369),
            .I(N__36366));
    LocalMux I__7323 (
            .O(N__36366),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__7322 (
            .O(N__36363),
            .I(N__36359));
    InMux I__7321 (
            .O(N__36362),
            .I(N__36356));
    LocalMux I__7320 (
            .O(N__36359),
            .I(N__36353));
    LocalMux I__7319 (
            .O(N__36356),
            .I(N__36350));
    Span4Mux_v I__7318 (
            .O(N__36353),
            .I(N__36347));
    Span4Mux_h I__7317 (
            .O(N__36350),
            .I(N__36344));
    Span4Mux_v I__7316 (
            .O(N__36347),
            .I(N__36341));
    Span4Mux_h I__7315 (
            .O(N__36344),
            .I(N__36338));
    Sp12to4 I__7314 (
            .O(N__36341),
            .I(N__36335));
    Odrv4 I__7313 (
            .O(N__36338),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv12 I__7312 (
            .O(N__36335),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__7311 (
            .O(N__36330),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__7310 (
            .O(N__36327),
            .I(N__36324));
    LocalMux I__7309 (
            .O(N__36324),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__7308 (
            .O(N__36321),
            .I(N__36317));
    InMux I__7307 (
            .O(N__36320),
            .I(N__36314));
    LocalMux I__7306 (
            .O(N__36317),
            .I(N__36311));
    LocalMux I__7305 (
            .O(N__36314),
            .I(N__36308));
    Span12Mux_s11_h I__7304 (
            .O(N__36311),
            .I(N__36305));
    Odrv12 I__7303 (
            .O(N__36308),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv12 I__7302 (
            .O(N__36305),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__7301 (
            .O(N__36300),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__7300 (
            .O(N__36297),
            .I(N__36294));
    LocalMux I__7299 (
            .O(N__36294),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__7298 (
            .O(N__36291),
            .I(bfn_14_19_0_));
    InMux I__7297 (
            .O(N__36288),
            .I(N__36285));
    LocalMux I__7296 (
            .O(N__36285),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__7295 (
            .O(N__36282),
            .I(N__36279));
    LocalMux I__7294 (
            .O(N__36279),
            .I(N__36276));
    Span4Mux_s2_h I__7293 (
            .O(N__36276),
            .I(N__36272));
    InMux I__7292 (
            .O(N__36275),
            .I(N__36269));
    Span4Mux_h I__7291 (
            .O(N__36272),
            .I(N__36266));
    LocalMux I__7290 (
            .O(N__36269),
            .I(N__36263));
    Span4Mux_h I__7289 (
            .O(N__36266),
            .I(N__36260));
    Span12Mux_s9_h I__7288 (
            .O(N__36263),
            .I(N__36257));
    Span4Mux_v I__7287 (
            .O(N__36260),
            .I(N__36254));
    Odrv12 I__7286 (
            .O(N__36257),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv4 I__7285 (
            .O(N__36254),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__7284 (
            .O(N__36249),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__7283 (
            .O(N__36246),
            .I(N__36243));
    LocalMux I__7282 (
            .O(N__36243),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__7281 (
            .O(N__36240),
            .I(N__36237));
    LocalMux I__7280 (
            .O(N__36237),
            .I(N__36234));
    Span4Mux_s3_h I__7279 (
            .O(N__36234),
            .I(N__36230));
    InMux I__7278 (
            .O(N__36233),
            .I(N__36227));
    Span4Mux_h I__7277 (
            .O(N__36230),
            .I(N__36224));
    LocalMux I__7276 (
            .O(N__36227),
            .I(N__36221));
    Span4Mux_h I__7275 (
            .O(N__36224),
            .I(N__36218));
    Span12Mux_s8_h I__7274 (
            .O(N__36221),
            .I(N__36215));
    Sp12to4 I__7273 (
            .O(N__36218),
            .I(N__36212));
    Odrv12 I__7272 (
            .O(N__36215),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv12 I__7271 (
            .O(N__36212),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__7270 (
            .O(N__36207),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__7269 (
            .O(N__36204),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__7268 (
            .O(N__36201),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    CEMux I__7267 (
            .O(N__36198),
            .I(N__36174));
    CEMux I__7266 (
            .O(N__36197),
            .I(N__36174));
    CEMux I__7265 (
            .O(N__36196),
            .I(N__36174));
    CEMux I__7264 (
            .O(N__36195),
            .I(N__36174));
    CEMux I__7263 (
            .O(N__36194),
            .I(N__36174));
    CEMux I__7262 (
            .O(N__36193),
            .I(N__36174));
    CEMux I__7261 (
            .O(N__36192),
            .I(N__36174));
    CEMux I__7260 (
            .O(N__36191),
            .I(N__36174));
    GlobalMux I__7259 (
            .O(N__36174),
            .I(N__36171));
    gio2CtrlBuf I__7258 (
            .O(N__36171),
            .I(\current_shift_inst.timer_s1.N_339_i_g ));
    InMux I__7257 (
            .O(N__36168),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    InMux I__7256 (
            .O(N__36165),
            .I(N__36161));
    InMux I__7255 (
            .O(N__36164),
            .I(N__36157));
    LocalMux I__7254 (
            .O(N__36161),
            .I(N__36154));
    InMux I__7253 (
            .O(N__36160),
            .I(N__36151));
    LocalMux I__7252 (
            .O(N__36157),
            .I(N__36148));
    Span4Mux_h I__7251 (
            .O(N__36154),
            .I(N__36145));
    LocalMux I__7250 (
            .O(N__36151),
            .I(N__36142));
    Span4Mux_v I__7249 (
            .O(N__36148),
            .I(N__36139));
    Span4Mux_h I__7248 (
            .O(N__36145),
            .I(N__36134));
    Span4Mux_v I__7247 (
            .O(N__36142),
            .I(N__36134));
    Span4Mux_h I__7246 (
            .O(N__36139),
            .I(N__36131));
    Odrv4 I__7245 (
            .O(N__36134),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__7244 (
            .O(N__36131),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CascadeMux I__7243 (
            .O(N__36126),
            .I(N__36122));
    InMux I__7242 (
            .O(N__36125),
            .I(N__36118));
    InMux I__7241 (
            .O(N__36122),
            .I(N__36115));
    InMux I__7240 (
            .O(N__36121),
            .I(N__36112));
    LocalMux I__7239 (
            .O(N__36118),
            .I(N__36109));
    LocalMux I__7238 (
            .O(N__36115),
            .I(N__36104));
    LocalMux I__7237 (
            .O(N__36112),
            .I(N__36104));
    Span4Mux_h I__7236 (
            .O(N__36109),
            .I(N__36098));
    Span4Mux_h I__7235 (
            .O(N__36104),
            .I(N__36098));
    InMux I__7234 (
            .O(N__36103),
            .I(N__36095));
    Odrv4 I__7233 (
            .O(N__36098),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__7232 (
            .O(N__36095),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__7231 (
            .O(N__36090),
            .I(N__36087));
    LocalMux I__7230 (
            .O(N__36087),
            .I(N__36084));
    Span4Mux_h I__7229 (
            .O(N__36084),
            .I(N__36081));
    Odrv4 I__7228 (
            .O(N__36081),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__7227 (
            .O(N__36078),
            .I(N__36074));
    InMux I__7226 (
            .O(N__36077),
            .I(N__36071));
    LocalMux I__7225 (
            .O(N__36074),
            .I(N__36068));
    LocalMux I__7224 (
            .O(N__36071),
            .I(N__36062));
    Span4Mux_h I__7223 (
            .O(N__36068),
            .I(N__36062));
    InMux I__7222 (
            .O(N__36067),
            .I(N__36059));
    Span4Mux_v I__7221 (
            .O(N__36062),
            .I(N__36053));
    LocalMux I__7220 (
            .O(N__36059),
            .I(N__36053));
    InMux I__7219 (
            .O(N__36058),
            .I(N__36050));
    Odrv4 I__7218 (
            .O(N__36053),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    LocalMux I__7217 (
            .O(N__36050),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__7216 (
            .O(N__36045),
            .I(N__36042));
    LocalMux I__7215 (
            .O(N__36042),
            .I(N__36039));
    Span4Mux_h I__7214 (
            .O(N__36039),
            .I(N__36036));
    Odrv4 I__7213 (
            .O(N__36036),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__7212 (
            .O(N__36033),
            .I(N__36030));
    LocalMux I__7211 (
            .O(N__36030),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__7210 (
            .O(N__36027),
            .I(N__36024));
    LocalMux I__7209 (
            .O(N__36024),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__7208 (
            .O(N__36021),
            .I(N__36018));
    LocalMux I__7207 (
            .O(N__36018),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__7206 (
            .O(N__36015),
            .I(N__36011));
    InMux I__7205 (
            .O(N__36014),
            .I(N__36008));
    LocalMux I__7204 (
            .O(N__36011),
            .I(N__36005));
    LocalMux I__7203 (
            .O(N__36008),
            .I(N__36002));
    Span4Mux_v I__7202 (
            .O(N__36005),
            .I(N__35999));
    Span4Mux_v I__7201 (
            .O(N__36002),
            .I(N__35996));
    Span4Mux_h I__7200 (
            .O(N__35999),
            .I(N__35993));
    Span4Mux_h I__7199 (
            .O(N__35996),
            .I(N__35990));
    Span4Mux_h I__7198 (
            .O(N__35993),
            .I(N__35987));
    Span4Mux_h I__7197 (
            .O(N__35990),
            .I(N__35982));
    Span4Mux_v I__7196 (
            .O(N__35987),
            .I(N__35982));
    Odrv4 I__7195 (
            .O(N__35982),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__7194 (
            .O(N__35979),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__7193 (
            .O(N__35976),
            .I(N__35973));
    LocalMux I__7192 (
            .O(N__35973),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__7191 (
            .O(N__35970),
            .I(N__35967));
    LocalMux I__7190 (
            .O(N__35967),
            .I(N__35963));
    InMux I__7189 (
            .O(N__35966),
            .I(N__35960));
    Span4Mux_v I__7188 (
            .O(N__35963),
            .I(N__35957));
    LocalMux I__7187 (
            .O(N__35960),
            .I(N__35954));
    Sp12to4 I__7186 (
            .O(N__35957),
            .I(N__35951));
    Span4Mux_h I__7185 (
            .O(N__35954),
            .I(N__35948));
    Span12Mux_s11_h I__7184 (
            .O(N__35951),
            .I(N__35945));
    Odrv4 I__7183 (
            .O(N__35948),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv12 I__7182 (
            .O(N__35945),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__7181 (
            .O(N__35940),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    CascadeMux I__7180 (
            .O(N__35937),
            .I(N__35933));
    CascadeMux I__7179 (
            .O(N__35936),
            .I(N__35930));
    InMux I__7178 (
            .O(N__35933),
            .I(N__35927));
    InMux I__7177 (
            .O(N__35930),
            .I(N__35924));
    LocalMux I__7176 (
            .O(N__35927),
            .I(N__35921));
    LocalMux I__7175 (
            .O(N__35924),
            .I(N__35918));
    Span4Mux_v I__7174 (
            .O(N__35921),
            .I(N__35914));
    Span4Mux_v I__7173 (
            .O(N__35918),
            .I(N__35911));
    InMux I__7172 (
            .O(N__35917),
            .I(N__35908));
    Span4Mux_h I__7171 (
            .O(N__35914),
            .I(N__35904));
    Span4Mux_h I__7170 (
            .O(N__35911),
            .I(N__35899));
    LocalMux I__7169 (
            .O(N__35908),
            .I(N__35899));
    InMux I__7168 (
            .O(N__35907),
            .I(N__35896));
    Odrv4 I__7167 (
            .O(N__35904),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__7166 (
            .O(N__35899),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    LocalMux I__7165 (
            .O(N__35896),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    InMux I__7164 (
            .O(N__35889),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__7163 (
            .O(N__35886),
            .I(N__35883));
    InMux I__7162 (
            .O(N__35883),
            .I(N__35879));
    CascadeMux I__7161 (
            .O(N__35882),
            .I(N__35876));
    LocalMux I__7160 (
            .O(N__35879),
            .I(N__35873));
    InMux I__7159 (
            .O(N__35876),
            .I(N__35870));
    Span4Mux_h I__7158 (
            .O(N__35873),
            .I(N__35865));
    LocalMux I__7157 (
            .O(N__35870),
            .I(N__35865));
    Span4Mux_h I__7156 (
            .O(N__35865),
            .I(N__35860));
    InMux I__7155 (
            .O(N__35864),
            .I(N__35857));
    InMux I__7154 (
            .O(N__35863),
            .I(N__35854));
    Odrv4 I__7153 (
            .O(N__35860),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__7152 (
            .O(N__35857),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__7151 (
            .O(N__35854),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__7150 (
            .O(N__35847),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__7149 (
            .O(N__35844),
            .I(N__35840));
    InMux I__7148 (
            .O(N__35843),
            .I(N__35837));
    InMux I__7147 (
            .O(N__35840),
            .I(N__35834));
    LocalMux I__7146 (
            .O(N__35837),
            .I(N__35830));
    LocalMux I__7145 (
            .O(N__35834),
            .I(N__35827));
    InMux I__7144 (
            .O(N__35833),
            .I(N__35824));
    Span4Mux_h I__7143 (
            .O(N__35830),
            .I(N__35818));
    Span4Mux_h I__7142 (
            .O(N__35827),
            .I(N__35818));
    LocalMux I__7141 (
            .O(N__35824),
            .I(N__35815));
    InMux I__7140 (
            .O(N__35823),
            .I(N__35812));
    Odrv4 I__7139 (
            .O(N__35818),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    Odrv4 I__7138 (
            .O(N__35815),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__7137 (
            .O(N__35812),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    InMux I__7136 (
            .O(N__35805),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__7135 (
            .O(N__35802),
            .I(N__35798));
    InMux I__7134 (
            .O(N__35801),
            .I(N__35795));
    InMux I__7133 (
            .O(N__35798),
            .I(N__35792));
    LocalMux I__7132 (
            .O(N__35795),
            .I(N__35788));
    LocalMux I__7131 (
            .O(N__35792),
            .I(N__35785));
    InMux I__7130 (
            .O(N__35791),
            .I(N__35782));
    Span4Mux_v I__7129 (
            .O(N__35788),
            .I(N__35779));
    Span4Mux_h I__7128 (
            .O(N__35785),
            .I(N__35774));
    LocalMux I__7127 (
            .O(N__35782),
            .I(N__35774));
    Span4Mux_h I__7126 (
            .O(N__35779),
            .I(N__35771));
    Span4Mux_v I__7125 (
            .O(N__35774),
            .I(N__35768));
    Span4Mux_v I__7124 (
            .O(N__35771),
            .I(N__35764));
    Span4Mux_h I__7123 (
            .O(N__35768),
            .I(N__35761));
    InMux I__7122 (
            .O(N__35767),
            .I(N__35758));
    Odrv4 I__7121 (
            .O(N__35764),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    Odrv4 I__7120 (
            .O(N__35761),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__7119 (
            .O(N__35758),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    InMux I__7118 (
            .O(N__35751),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__7117 (
            .O(N__35748),
            .I(N__35745));
    InMux I__7116 (
            .O(N__35745),
            .I(N__35741));
    InMux I__7115 (
            .O(N__35744),
            .I(N__35738));
    LocalMux I__7114 (
            .O(N__35741),
            .I(N__35734));
    LocalMux I__7113 (
            .O(N__35738),
            .I(N__35731));
    InMux I__7112 (
            .O(N__35737),
            .I(N__35728));
    Span4Mux_v I__7111 (
            .O(N__35734),
            .I(N__35725));
    Span4Mux_h I__7110 (
            .O(N__35731),
            .I(N__35722));
    LocalMux I__7109 (
            .O(N__35728),
            .I(N__35719));
    Sp12to4 I__7108 (
            .O(N__35725),
            .I(N__35715));
    Span4Mux_h I__7107 (
            .O(N__35722),
            .I(N__35712));
    Span4Mux_v I__7106 (
            .O(N__35719),
            .I(N__35709));
    InMux I__7105 (
            .O(N__35718),
            .I(N__35706));
    Odrv12 I__7104 (
            .O(N__35715),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__7103 (
            .O(N__35712),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__7102 (
            .O(N__35709),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__7101 (
            .O(N__35706),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__7100 (
            .O(N__35697),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__7099 (
            .O(N__35694),
            .I(N__35691));
    LocalMux I__7098 (
            .O(N__35691),
            .I(N__35687));
    InMux I__7097 (
            .O(N__35690),
            .I(N__35684));
    Span4Mux_v I__7096 (
            .O(N__35687),
            .I(N__35678));
    LocalMux I__7095 (
            .O(N__35684),
            .I(N__35678));
    InMux I__7094 (
            .O(N__35683),
            .I(N__35674));
    Span4Mux_h I__7093 (
            .O(N__35678),
            .I(N__35671));
    InMux I__7092 (
            .O(N__35677),
            .I(N__35668));
    LocalMux I__7091 (
            .O(N__35674),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__7090 (
            .O(N__35671),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    LocalMux I__7089 (
            .O(N__35668),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__7088 (
            .O(N__35661),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__7087 (
            .O(N__35658),
            .I(N__35655));
    InMux I__7086 (
            .O(N__35655),
            .I(N__35651));
    CascadeMux I__7085 (
            .O(N__35654),
            .I(N__35648));
    LocalMux I__7084 (
            .O(N__35651),
            .I(N__35645));
    InMux I__7083 (
            .O(N__35648),
            .I(N__35642));
    Span4Mux_v I__7082 (
            .O(N__35645),
            .I(N__35636));
    LocalMux I__7081 (
            .O(N__35642),
            .I(N__35636));
    InMux I__7080 (
            .O(N__35641),
            .I(N__35633));
    Span4Mux_h I__7079 (
            .O(N__35636),
            .I(N__35629));
    LocalMux I__7078 (
            .O(N__35633),
            .I(N__35626));
    InMux I__7077 (
            .O(N__35632),
            .I(N__35623));
    Odrv4 I__7076 (
            .O(N__35629),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__7075 (
            .O(N__35626),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    LocalMux I__7074 (
            .O(N__35623),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__7073 (
            .O(N__35616),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7072 (
            .O(N__35613),
            .I(N__35609));
    InMux I__7071 (
            .O(N__35612),
            .I(N__35606));
    InMux I__7070 (
            .O(N__35609),
            .I(N__35603));
    LocalMux I__7069 (
            .O(N__35606),
            .I(N__35597));
    LocalMux I__7068 (
            .O(N__35603),
            .I(N__35597));
    InMux I__7067 (
            .O(N__35602),
            .I(N__35594));
    Span4Mux_v I__7066 (
            .O(N__35597),
            .I(N__35589));
    LocalMux I__7065 (
            .O(N__35594),
            .I(N__35589));
    Span4Mux_h I__7064 (
            .O(N__35589),
            .I(N__35585));
    InMux I__7063 (
            .O(N__35588),
            .I(N__35582));
    Odrv4 I__7062 (
            .O(N__35585),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    LocalMux I__7061 (
            .O(N__35582),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__7060 (
            .O(N__35577),
            .I(bfn_14_17_0_));
    InMux I__7059 (
            .O(N__35574),
            .I(N__35568));
    InMux I__7058 (
            .O(N__35573),
            .I(N__35568));
    LocalMux I__7057 (
            .O(N__35568),
            .I(N__35564));
    InMux I__7056 (
            .O(N__35567),
            .I(N__35561));
    Span4Mux_v I__7055 (
            .O(N__35564),
            .I(N__35556));
    LocalMux I__7054 (
            .O(N__35561),
            .I(N__35556));
    Span4Mux_h I__7053 (
            .O(N__35556),
            .I(N__35552));
    InMux I__7052 (
            .O(N__35555),
            .I(N__35549));
    Odrv4 I__7051 (
            .O(N__35552),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__7050 (
            .O(N__35549),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__7049 (
            .O(N__35544),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__7048 (
            .O(N__35541),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__7047 (
            .O(N__35538),
            .I(N__35535));
    InMux I__7046 (
            .O(N__35535),
            .I(N__35531));
    InMux I__7045 (
            .O(N__35534),
            .I(N__35528));
    LocalMux I__7044 (
            .O(N__35531),
            .I(N__35524));
    LocalMux I__7043 (
            .O(N__35528),
            .I(N__35521));
    InMux I__7042 (
            .O(N__35527),
            .I(N__35518));
    Span4Mux_h I__7041 (
            .O(N__35524),
            .I(N__35515));
    Span4Mux_v I__7040 (
            .O(N__35521),
            .I(N__35512));
    LocalMux I__7039 (
            .O(N__35518),
            .I(N__35509));
    Span4Mux_h I__7038 (
            .O(N__35515),
            .I(N__35505));
    Span4Mux_h I__7037 (
            .O(N__35512),
            .I(N__35500));
    Span4Mux_v I__7036 (
            .O(N__35509),
            .I(N__35500));
    InMux I__7035 (
            .O(N__35508),
            .I(N__35497));
    Odrv4 I__7034 (
            .O(N__35505),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    Odrv4 I__7033 (
            .O(N__35500),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__7032 (
            .O(N__35497),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__7031 (
            .O(N__35490),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__7030 (
            .O(N__35487),
            .I(N__35484));
    LocalMux I__7029 (
            .O(N__35484),
            .I(N__35479));
    InMux I__7028 (
            .O(N__35483),
            .I(N__35476));
    InMux I__7027 (
            .O(N__35482),
            .I(N__35473));
    Span4Mux_v I__7026 (
            .O(N__35479),
            .I(N__35468));
    LocalMux I__7025 (
            .O(N__35476),
            .I(N__35468));
    LocalMux I__7024 (
            .O(N__35473),
            .I(N__35465));
    Span4Mux_h I__7023 (
            .O(N__35468),
            .I(N__35461));
    Span4Mux_v I__7022 (
            .O(N__35465),
            .I(N__35458));
    InMux I__7021 (
            .O(N__35464),
            .I(N__35455));
    Odrv4 I__7020 (
            .O(N__35461),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv4 I__7019 (
            .O(N__35458),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__7018 (
            .O(N__35455),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__7017 (
            .O(N__35448),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__7016 (
            .O(N__35445),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__7015 (
            .O(N__35442),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7014 (
            .O(N__35439),
            .I(N__35435));
    InMux I__7013 (
            .O(N__35438),
            .I(N__35432));
    InMux I__7012 (
            .O(N__35435),
            .I(N__35428));
    LocalMux I__7011 (
            .O(N__35432),
            .I(N__35425));
    InMux I__7010 (
            .O(N__35431),
            .I(N__35422));
    LocalMux I__7009 (
            .O(N__35428),
            .I(N__35417));
    Span4Mux_h I__7008 (
            .O(N__35425),
            .I(N__35417));
    LocalMux I__7007 (
            .O(N__35422),
            .I(N__35414));
    Span4Mux_h I__7006 (
            .O(N__35417),
            .I(N__35408));
    Span4Mux_h I__7005 (
            .O(N__35414),
            .I(N__35408));
    InMux I__7004 (
            .O(N__35413),
            .I(N__35405));
    Odrv4 I__7003 (
            .O(N__35408),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__7002 (
            .O(N__35405),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    InMux I__7001 (
            .O(N__35400),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    InMux I__7000 (
            .O(N__35397),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    InMux I__6999 (
            .O(N__35394),
            .I(N__35390));
    InMux I__6998 (
            .O(N__35393),
            .I(N__35387));
    LocalMux I__6997 (
            .O(N__35390),
            .I(N__35383));
    LocalMux I__6996 (
            .O(N__35387),
            .I(N__35380));
    InMux I__6995 (
            .O(N__35386),
            .I(N__35377));
    Span12Mux_v I__6994 (
            .O(N__35383),
            .I(N__35371));
    Span12Mux_v I__6993 (
            .O(N__35380),
            .I(N__35371));
    LocalMux I__6992 (
            .O(N__35377),
            .I(N__35368));
    InMux I__6991 (
            .O(N__35376),
            .I(N__35365));
    Odrv12 I__6990 (
            .O(N__35371),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__6989 (
            .O(N__35368),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    LocalMux I__6988 (
            .O(N__35365),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    InMux I__6987 (
            .O(N__35358),
            .I(bfn_14_16_0_));
    CascadeMux I__6986 (
            .O(N__35355),
            .I(N__35352));
    InMux I__6985 (
            .O(N__35352),
            .I(N__35348));
    InMux I__6984 (
            .O(N__35351),
            .I(N__35345));
    LocalMux I__6983 (
            .O(N__35348),
            .I(N__35341));
    LocalMux I__6982 (
            .O(N__35345),
            .I(N__35338));
    InMux I__6981 (
            .O(N__35344),
            .I(N__35335));
    Span4Mux_v I__6980 (
            .O(N__35341),
            .I(N__35328));
    Span4Mux_v I__6979 (
            .O(N__35338),
            .I(N__35328));
    LocalMux I__6978 (
            .O(N__35335),
            .I(N__35328));
    Span4Mux_h I__6977 (
            .O(N__35328),
            .I(N__35324));
    InMux I__6976 (
            .O(N__35327),
            .I(N__35321));
    Odrv4 I__6975 (
            .O(N__35324),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__6974 (
            .O(N__35321),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__6973 (
            .O(N__35316),
            .I(N__35312));
    InMux I__6972 (
            .O(N__35315),
            .I(N__35309));
    LocalMux I__6971 (
            .O(N__35312),
            .I(N__35306));
    LocalMux I__6970 (
            .O(N__35309),
            .I(N__35303));
    Span4Mux_v I__6969 (
            .O(N__35306),
            .I(N__35300));
    Span4Mux_h I__6968 (
            .O(N__35303),
            .I(N__35297));
    Span4Mux_h I__6967 (
            .O(N__35300),
            .I(N__35292));
    Span4Mux_h I__6966 (
            .O(N__35297),
            .I(N__35289));
    InMux I__6965 (
            .O(N__35296),
            .I(N__35284));
    InMux I__6964 (
            .O(N__35295),
            .I(N__35284));
    Odrv4 I__6963 (
            .O(N__35292),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    Odrv4 I__6962 (
            .O(N__35289),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__6961 (
            .O(N__35284),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__6960 (
            .O(N__35277),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    InMux I__6959 (
            .O(N__35274),
            .I(N__35270));
    InMux I__6958 (
            .O(N__35273),
            .I(N__35267));
    LocalMux I__6957 (
            .O(N__35270),
            .I(N__35264));
    LocalMux I__6956 (
            .O(N__35267),
            .I(N__35261));
    Span4Mux_v I__6955 (
            .O(N__35264),
            .I(N__35256));
    Span4Mux_h I__6954 (
            .O(N__35261),
            .I(N__35253));
    InMux I__6953 (
            .O(N__35260),
            .I(N__35248));
    InMux I__6952 (
            .O(N__35259),
            .I(N__35248));
    Odrv4 I__6951 (
            .O(N__35256),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__6950 (
            .O(N__35253),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__6949 (
            .O(N__35248),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__6948 (
            .O(N__35241),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    InMux I__6947 (
            .O(N__35238),
            .I(N__35234));
    CascadeMux I__6946 (
            .O(N__35237),
            .I(N__35231));
    LocalMux I__6945 (
            .O(N__35234),
            .I(N__35228));
    InMux I__6944 (
            .O(N__35231),
            .I(N__35225));
    Span4Mux_v I__6943 (
            .O(N__35228),
            .I(N__35219));
    LocalMux I__6942 (
            .O(N__35225),
            .I(N__35219));
    InMux I__6941 (
            .O(N__35224),
            .I(N__35216));
    Span4Mux_h I__6940 (
            .O(N__35219),
            .I(N__35211));
    LocalMux I__6939 (
            .O(N__35216),
            .I(N__35211));
    Span4Mux_h I__6938 (
            .O(N__35211),
            .I(N__35207));
    InMux I__6937 (
            .O(N__35210),
            .I(N__35204));
    Odrv4 I__6936 (
            .O(N__35207),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__6935 (
            .O(N__35204),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__6934 (
            .O(N__35199),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__6933 (
            .O(N__35196),
            .I(N__35192));
    CascadeMux I__6932 (
            .O(N__35195),
            .I(N__35189));
    InMux I__6931 (
            .O(N__35192),
            .I(N__35186));
    InMux I__6930 (
            .O(N__35189),
            .I(N__35183));
    LocalMux I__6929 (
            .O(N__35186),
            .I(N__35179));
    LocalMux I__6928 (
            .O(N__35183),
            .I(N__35176));
    InMux I__6927 (
            .O(N__35182),
            .I(N__35173));
    Span4Mux_h I__6926 (
            .O(N__35179),
            .I(N__35170));
    Span4Mux_v I__6925 (
            .O(N__35176),
            .I(N__35165));
    LocalMux I__6924 (
            .O(N__35173),
            .I(N__35165));
    Span4Mux_h I__6923 (
            .O(N__35170),
            .I(N__35161));
    Span4Mux_h I__6922 (
            .O(N__35165),
            .I(N__35158));
    InMux I__6921 (
            .O(N__35164),
            .I(N__35155));
    Odrv4 I__6920 (
            .O(N__35161),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__6919 (
            .O(N__35158),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__6918 (
            .O(N__35155),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__6917 (
            .O(N__35148),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    InMux I__6916 (
            .O(N__35145),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__6915 (
            .O(N__35142),
            .I(N__35139));
    InMux I__6914 (
            .O(N__35139),
            .I(N__35135));
    CascadeMux I__6913 (
            .O(N__35138),
            .I(N__35132));
    LocalMux I__6912 (
            .O(N__35135),
            .I(N__35128));
    InMux I__6911 (
            .O(N__35132),
            .I(N__35125));
    InMux I__6910 (
            .O(N__35131),
            .I(N__35122));
    Span4Mux_h I__6909 (
            .O(N__35128),
            .I(N__35119));
    LocalMux I__6908 (
            .O(N__35125),
            .I(N__35114));
    LocalMux I__6907 (
            .O(N__35122),
            .I(N__35114));
    Span4Mux_h I__6906 (
            .O(N__35119),
            .I(N__35110));
    Span4Mux_v I__6905 (
            .O(N__35114),
            .I(N__35107));
    InMux I__6904 (
            .O(N__35113),
            .I(N__35104));
    Odrv4 I__6903 (
            .O(N__35110),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    Odrv4 I__6902 (
            .O(N__35107),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__6901 (
            .O(N__35104),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__6900 (
            .O(N__35097),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    InMux I__6899 (
            .O(N__35094),
            .I(N__35090));
    InMux I__6898 (
            .O(N__35093),
            .I(N__35087));
    LocalMux I__6897 (
            .O(N__35090),
            .I(N__35081));
    LocalMux I__6896 (
            .O(N__35087),
            .I(N__35081));
    InMux I__6895 (
            .O(N__35086),
            .I(N__35078));
    Span4Mux_v I__6894 (
            .O(N__35081),
            .I(N__35073));
    LocalMux I__6893 (
            .O(N__35078),
            .I(N__35073));
    Span4Mux_h I__6892 (
            .O(N__35073),
            .I(N__35069));
    InMux I__6891 (
            .O(N__35072),
            .I(N__35066));
    Odrv4 I__6890 (
            .O(N__35069),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__6889 (
            .O(N__35066),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    InMux I__6888 (
            .O(N__35061),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__6887 (
            .O(N__35058),
            .I(N__35055));
    InMux I__6886 (
            .O(N__35055),
            .I(N__35052));
    LocalMux I__6885 (
            .O(N__35052),
            .I(N__35047));
    InMux I__6884 (
            .O(N__35051),
            .I(N__35042));
    InMux I__6883 (
            .O(N__35050),
            .I(N__35042));
    Span4Mux_h I__6882 (
            .O(N__35047),
            .I(N__35039));
    LocalMux I__6881 (
            .O(N__35042),
            .I(N__35036));
    Span4Mux_h I__6880 (
            .O(N__35039),
            .I(N__35032));
    Span12Mux_v I__6879 (
            .O(N__35036),
            .I(N__35029));
    InMux I__6878 (
            .O(N__35035),
            .I(N__35026));
    Odrv4 I__6877 (
            .O(N__35032),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv12 I__6876 (
            .O(N__35029),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__6875 (
            .O(N__35026),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__6874 (
            .O(N__35019),
            .I(bfn_14_15_0_));
    InMux I__6873 (
            .O(N__35016),
            .I(N__35012));
    InMux I__6872 (
            .O(N__35015),
            .I(N__35009));
    LocalMux I__6871 (
            .O(N__35012),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    LocalMux I__6870 (
            .O(N__35009),
            .I(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ));
    CEMux I__6869 (
            .O(N__35004),
            .I(N__35001));
    LocalMux I__6868 (
            .O(N__35001),
            .I(N__34998));
    Odrv4 I__6867 (
            .O(N__34998),
            .I(\phase_controller_inst2.stoper_hc.N_266_0 ));
    InMux I__6866 (
            .O(N__34995),
            .I(N__34991));
    InMux I__6865 (
            .O(N__34994),
            .I(N__34987));
    LocalMux I__6864 (
            .O(N__34991),
            .I(N__34984));
    InMux I__6863 (
            .O(N__34990),
            .I(N__34981));
    LocalMux I__6862 (
            .O(N__34987),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    Odrv4 I__6861 (
            .O(N__34984),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    LocalMux I__6860 (
            .O(N__34981),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    InMux I__6859 (
            .O(N__34974),
            .I(N__34969));
    InMux I__6858 (
            .O(N__34973),
            .I(N__34966));
    InMux I__6857 (
            .O(N__34972),
            .I(N__34963));
    LocalMux I__6856 (
            .O(N__34969),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__6855 (
            .O(N__34966),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    LocalMux I__6854 (
            .O(N__34963),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    ClkMux I__6853 (
            .O(N__34956),
            .I(N__34953));
    GlobalMux I__6852 (
            .O(N__34953),
            .I(N__34950));
    gio2CtrlBuf I__6851 (
            .O(N__34950),
            .I(delay_hc_input_c_g));
    InMux I__6850 (
            .O(N__34947),
            .I(N__34944));
    LocalMux I__6849 (
            .O(N__34944),
            .I(N__34941));
    Odrv12 I__6848 (
            .O(N__34941),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    CascadeMux I__6847 (
            .O(N__34938),
            .I(N__34934));
    InMux I__6846 (
            .O(N__34937),
            .I(N__34930));
    InMux I__6845 (
            .O(N__34934),
            .I(N__34927));
    InMux I__6844 (
            .O(N__34933),
            .I(N__34924));
    LocalMux I__6843 (
            .O(N__34930),
            .I(N__34919));
    LocalMux I__6842 (
            .O(N__34927),
            .I(N__34919));
    LocalMux I__6841 (
            .O(N__34924),
            .I(N__34914));
    Span4Mux_s3_v I__6840 (
            .O(N__34919),
            .I(N__34914));
    Odrv4 I__6839 (
            .O(N__34914),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__6838 (
            .O(N__34911),
            .I(N__34908));
    LocalMux I__6837 (
            .O(N__34908),
            .I(N__34901));
    InMux I__6836 (
            .O(N__34907),
            .I(N__34896));
    InMux I__6835 (
            .O(N__34906),
            .I(N__34896));
    InMux I__6834 (
            .O(N__34905),
            .I(N__34893));
    InMux I__6833 (
            .O(N__34904),
            .I(N__34890));
    Span12Mux_v I__6832 (
            .O(N__34901),
            .I(N__34887));
    LocalMux I__6831 (
            .O(N__34896),
            .I(\phase_controller_inst2.N_139_1 ));
    LocalMux I__6830 (
            .O(N__34893),
            .I(\phase_controller_inst2.N_139_1 ));
    LocalMux I__6829 (
            .O(N__34890),
            .I(\phase_controller_inst2.N_139_1 ));
    Odrv12 I__6828 (
            .O(N__34887),
            .I(\phase_controller_inst2.N_139_1 ));
    InMux I__6827 (
            .O(N__34878),
            .I(N__34875));
    LocalMux I__6826 (
            .O(N__34875),
            .I(\phase_controller_inst2.stoper_hc.N_34 ));
    InMux I__6825 (
            .O(N__34872),
            .I(N__34869));
    LocalMux I__6824 (
            .O(N__34869),
            .I(\phase_controller_inst2.stoper_hc.m20_nsZ0Z_1 ));
    InMux I__6823 (
            .O(N__34866),
            .I(N__34860));
    InMux I__6822 (
            .O(N__34865),
            .I(N__34856));
    InMux I__6821 (
            .O(N__34864),
            .I(N__34853));
    InMux I__6820 (
            .O(N__34863),
            .I(N__34850));
    LocalMux I__6819 (
            .O(N__34860),
            .I(N__34847));
    InMux I__6818 (
            .O(N__34859),
            .I(N__34844));
    LocalMux I__6817 (
            .O(N__34856),
            .I(N__34839));
    LocalMux I__6816 (
            .O(N__34853),
            .I(N__34839));
    LocalMux I__6815 (
            .O(N__34850),
            .I(N__34836));
    Span4Mux_v I__6814 (
            .O(N__34847),
            .I(N__34831));
    LocalMux I__6813 (
            .O(N__34844),
            .I(N__34831));
    Span4Mux_h I__6812 (
            .O(N__34839),
            .I(N__34826));
    Span4Mux_h I__6811 (
            .O(N__34836),
            .I(N__34826));
    Span4Mux_h I__6810 (
            .O(N__34831),
            .I(N__34823));
    Span4Mux_h I__6809 (
            .O(N__34826),
            .I(N__34820));
    Span4Mux_h I__6808 (
            .O(N__34823),
            .I(N__34817));
    Odrv4 I__6807 (
            .O(N__34820),
            .I(il_min_comp2_c));
    Odrv4 I__6806 (
            .O(N__34817),
            .I(il_min_comp2_c));
    CascadeMux I__6805 (
            .O(N__34812),
            .I(N__34809));
    InMux I__6804 (
            .O(N__34809),
            .I(N__34805));
    InMux I__6803 (
            .O(N__34808),
            .I(N__34800));
    LocalMux I__6802 (
            .O(N__34805),
            .I(N__34796));
    InMux I__6801 (
            .O(N__34804),
            .I(N__34791));
    InMux I__6800 (
            .O(N__34803),
            .I(N__34791));
    LocalMux I__6799 (
            .O(N__34800),
            .I(N__34788));
    InMux I__6798 (
            .O(N__34799),
            .I(N__34785));
    Span4Mux_h I__6797 (
            .O(N__34796),
            .I(N__34780));
    LocalMux I__6796 (
            .O(N__34791),
            .I(N__34780));
    Odrv12 I__6795 (
            .O(N__34788),
            .I(\phase_controller_inst2.stoper_hc.hc_time_passed ));
    LocalMux I__6794 (
            .O(N__34785),
            .I(\phase_controller_inst2.stoper_hc.hc_time_passed ));
    Odrv4 I__6793 (
            .O(N__34780),
            .I(\phase_controller_inst2.stoper_hc.hc_time_passed ));
    InMux I__6792 (
            .O(N__34773),
            .I(N__34770));
    LocalMux I__6791 (
            .O(N__34770),
            .I(N__34767));
    Odrv12 I__6790 (
            .O(N__34767),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__6789 (
            .O(N__34764),
            .I(\current_shift_inst.control_input_cry_27 ));
    InMux I__6788 (
            .O(N__34761),
            .I(N__34758));
    LocalMux I__6787 (
            .O(N__34758),
            .I(\current_shift_inst.control_input_axb_29 ));
    InMux I__6786 (
            .O(N__34755),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__6785 (
            .O(N__34752),
            .I(N__34747));
    InMux I__6784 (
            .O(N__34751),
            .I(N__34744));
    CascadeMux I__6783 (
            .O(N__34750),
            .I(N__34741));
    LocalMux I__6782 (
            .O(N__34747),
            .I(N__34737));
    LocalMux I__6781 (
            .O(N__34744),
            .I(N__34734));
    InMux I__6780 (
            .O(N__34741),
            .I(N__34731));
    InMux I__6779 (
            .O(N__34740),
            .I(N__34723));
    Span4Mux_h I__6778 (
            .O(N__34737),
            .I(N__34713));
    Span4Mux_h I__6777 (
            .O(N__34734),
            .I(N__34692));
    LocalMux I__6776 (
            .O(N__34731),
            .I(N__34692));
    InMux I__6775 (
            .O(N__34730),
            .I(N__34681));
    InMux I__6774 (
            .O(N__34729),
            .I(N__34681));
    InMux I__6773 (
            .O(N__34728),
            .I(N__34681));
    InMux I__6772 (
            .O(N__34727),
            .I(N__34681));
    InMux I__6771 (
            .O(N__34726),
            .I(N__34681));
    LocalMux I__6770 (
            .O(N__34723),
            .I(N__34678));
    InMux I__6769 (
            .O(N__34722),
            .I(N__34667));
    InMux I__6768 (
            .O(N__34721),
            .I(N__34667));
    InMux I__6767 (
            .O(N__34720),
            .I(N__34667));
    InMux I__6766 (
            .O(N__34719),
            .I(N__34667));
    InMux I__6765 (
            .O(N__34718),
            .I(N__34667));
    InMux I__6764 (
            .O(N__34717),
            .I(N__34662));
    InMux I__6763 (
            .O(N__34716),
            .I(N__34662));
    Span4Mux_v I__6762 (
            .O(N__34713),
            .I(N__34659));
    InMux I__6761 (
            .O(N__34712),
            .I(N__34644));
    InMux I__6760 (
            .O(N__34711),
            .I(N__34644));
    InMux I__6759 (
            .O(N__34710),
            .I(N__34644));
    InMux I__6758 (
            .O(N__34709),
            .I(N__34644));
    InMux I__6757 (
            .O(N__34708),
            .I(N__34644));
    InMux I__6756 (
            .O(N__34707),
            .I(N__34644));
    InMux I__6755 (
            .O(N__34706),
            .I(N__34644));
    InMux I__6754 (
            .O(N__34705),
            .I(N__34635));
    InMux I__6753 (
            .O(N__34704),
            .I(N__34635));
    InMux I__6752 (
            .O(N__34703),
            .I(N__34635));
    InMux I__6751 (
            .O(N__34702),
            .I(N__34635));
    InMux I__6750 (
            .O(N__34701),
            .I(N__34624));
    InMux I__6749 (
            .O(N__34700),
            .I(N__34624));
    InMux I__6748 (
            .O(N__34699),
            .I(N__34624));
    InMux I__6747 (
            .O(N__34698),
            .I(N__34624));
    InMux I__6746 (
            .O(N__34697),
            .I(N__34624));
    Span4Mux_h I__6745 (
            .O(N__34692),
            .I(N__34619));
    LocalMux I__6744 (
            .O(N__34681),
            .I(N__34619));
    Odrv4 I__6743 (
            .O(N__34678),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__6742 (
            .O(N__34667),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__6741 (
            .O(N__34662),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__6740 (
            .O(N__34659),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__6739 (
            .O(N__34644),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__6738 (
            .O(N__34635),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__6737 (
            .O(N__34624),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__6736 (
            .O(N__34619),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__6735 (
            .O(N__34602),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__6734 (
            .O(N__34599),
            .I(N__34596));
    LocalMux I__6733 (
            .O(N__34596),
            .I(N__34593));
    Odrv4 I__6732 (
            .O(N__34593),
            .I(\current_shift_inst.control_input_axb_19 ));
    InMux I__6731 (
            .O(N__34590),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__6730 (
            .O(N__34587),
            .I(N__34584));
    LocalMux I__6729 (
            .O(N__34584),
            .I(\current_shift_inst.control_input_axb_20 ));
    InMux I__6728 (
            .O(N__34581),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__6727 (
            .O(N__34578),
            .I(N__34575));
    LocalMux I__6726 (
            .O(N__34575),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__6725 (
            .O(N__34572),
            .I(\current_shift_inst.control_input_cry_20 ));
    InMux I__6724 (
            .O(N__34569),
            .I(N__34566));
    LocalMux I__6723 (
            .O(N__34566),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__6722 (
            .O(N__34563),
            .I(\current_shift_inst.control_input_cry_21 ));
    InMux I__6721 (
            .O(N__34560),
            .I(N__34557));
    LocalMux I__6720 (
            .O(N__34557),
            .I(\current_shift_inst.control_input_axb_23 ));
    InMux I__6719 (
            .O(N__34554),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__6718 (
            .O(N__34551),
            .I(N__34548));
    LocalMux I__6717 (
            .O(N__34548),
            .I(N__34545));
    Odrv12 I__6716 (
            .O(N__34545),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__6715 (
            .O(N__34542),
            .I(bfn_13_20_0_));
    InMux I__6714 (
            .O(N__34539),
            .I(N__34536));
    LocalMux I__6713 (
            .O(N__34536),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__6712 (
            .O(N__34533),
            .I(\current_shift_inst.control_input_cry_24 ));
    InMux I__6711 (
            .O(N__34530),
            .I(N__34527));
    LocalMux I__6710 (
            .O(N__34527),
            .I(N__34524));
    Odrv4 I__6709 (
            .O(N__34524),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__6708 (
            .O(N__34521),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__6707 (
            .O(N__34518),
            .I(N__34515));
    LocalMux I__6706 (
            .O(N__34515),
            .I(N__34512));
    Odrv4 I__6705 (
            .O(N__34512),
            .I(\current_shift_inst.control_input_axb_27 ));
    InMux I__6704 (
            .O(N__34509),
            .I(\current_shift_inst.control_input_cry_26 ));
    InMux I__6703 (
            .O(N__34506),
            .I(N__34503));
    LocalMux I__6702 (
            .O(N__34503),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__6701 (
            .O(N__34500),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__6700 (
            .O(N__34497),
            .I(N__34494));
    LocalMux I__6699 (
            .O(N__34494),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__6698 (
            .O(N__34491),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__6697 (
            .O(N__34488),
            .I(N__34485));
    LocalMux I__6696 (
            .O(N__34485),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__6695 (
            .O(N__34482),
            .I(\current_shift_inst.control_input_cry_12 ));
    InMux I__6694 (
            .O(N__34479),
            .I(N__34476));
    LocalMux I__6693 (
            .O(N__34476),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__6692 (
            .O(N__34473),
            .I(\current_shift_inst.control_input_cry_13 ));
    InMux I__6691 (
            .O(N__34470),
            .I(N__34467));
    LocalMux I__6690 (
            .O(N__34467),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__6689 (
            .O(N__34464),
            .I(\current_shift_inst.control_input_cry_14 ));
    InMux I__6688 (
            .O(N__34461),
            .I(N__34458));
    LocalMux I__6687 (
            .O(N__34458),
            .I(N__34455));
    Odrv12 I__6686 (
            .O(N__34455),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__6685 (
            .O(N__34452),
            .I(bfn_13_19_0_));
    InMux I__6684 (
            .O(N__34449),
            .I(N__34446));
    LocalMux I__6683 (
            .O(N__34446),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__6682 (
            .O(N__34443),
            .I(\current_shift_inst.control_input_cry_16 ));
    CascadeMux I__6681 (
            .O(N__34440),
            .I(N__34437));
    InMux I__6680 (
            .O(N__34437),
            .I(N__34434));
    LocalMux I__6679 (
            .O(N__34434),
            .I(N__34431));
    Odrv4 I__6678 (
            .O(N__34431),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__6677 (
            .O(N__34428),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__6676 (
            .O(N__34425),
            .I(N__34422));
    LocalMux I__6675 (
            .O(N__34422),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__6674 (
            .O(N__34419),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__6673 (
            .O(N__34416),
            .I(N__34413));
    LocalMux I__6672 (
            .O(N__34413),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__6671 (
            .O(N__34410),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__6670 (
            .O(N__34407),
            .I(N__34404));
    LocalMux I__6669 (
            .O(N__34404),
            .I(N__34401));
    Span4Mux_v I__6668 (
            .O(N__34401),
            .I(N__34398));
    Odrv4 I__6667 (
            .O(N__34398),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__6666 (
            .O(N__34395),
            .I(\current_shift_inst.control_input_cry_4 ));
    InMux I__6665 (
            .O(N__34392),
            .I(N__34389));
    LocalMux I__6664 (
            .O(N__34389),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__6663 (
            .O(N__34386),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__6662 (
            .O(N__34383),
            .I(N__34380));
    LocalMux I__6661 (
            .O(N__34380),
            .I(N__34377));
    Span4Mux_h I__6660 (
            .O(N__34377),
            .I(N__34374));
    Odrv4 I__6659 (
            .O(N__34374),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__6658 (
            .O(N__34371),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__6657 (
            .O(N__34368),
            .I(N__34365));
    LocalMux I__6656 (
            .O(N__34365),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__6655 (
            .O(N__34362),
            .I(bfn_13_18_0_));
    InMux I__6654 (
            .O(N__34359),
            .I(N__34356));
    LocalMux I__6653 (
            .O(N__34356),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__6652 (
            .O(N__34353),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__6651 (
            .O(N__34350),
            .I(N__34347));
    LocalMux I__6650 (
            .O(N__34347),
            .I(\current_shift_inst.control_input_axb_10 ));
    InMux I__6649 (
            .O(N__34344),
            .I(\current_shift_inst.control_input_cry_9 ));
    CascadeMux I__6648 (
            .O(N__34341),
            .I(N__34321));
    InMux I__6647 (
            .O(N__34340),
            .I(N__34308));
    InMux I__6646 (
            .O(N__34339),
            .I(N__34303));
    InMux I__6645 (
            .O(N__34338),
            .I(N__34303));
    InMux I__6644 (
            .O(N__34337),
            .I(N__34300));
    InMux I__6643 (
            .O(N__34336),
            .I(N__34297));
    InMux I__6642 (
            .O(N__34335),
            .I(N__34290));
    InMux I__6641 (
            .O(N__34334),
            .I(N__34290));
    InMux I__6640 (
            .O(N__34333),
            .I(N__34290));
    InMux I__6639 (
            .O(N__34332),
            .I(N__34279));
    InMux I__6638 (
            .O(N__34331),
            .I(N__34274));
    InMux I__6637 (
            .O(N__34330),
            .I(N__34274));
    InMux I__6636 (
            .O(N__34329),
            .I(N__34269));
    InMux I__6635 (
            .O(N__34328),
            .I(N__34269));
    InMux I__6634 (
            .O(N__34327),
            .I(N__34262));
    InMux I__6633 (
            .O(N__34326),
            .I(N__34262));
    InMux I__6632 (
            .O(N__34325),
            .I(N__34262));
    InMux I__6631 (
            .O(N__34324),
            .I(N__34249));
    InMux I__6630 (
            .O(N__34321),
            .I(N__34249));
    InMux I__6629 (
            .O(N__34320),
            .I(N__34249));
    InMux I__6628 (
            .O(N__34319),
            .I(N__34249));
    InMux I__6627 (
            .O(N__34318),
            .I(N__34249));
    InMux I__6626 (
            .O(N__34317),
            .I(N__34249));
    InMux I__6625 (
            .O(N__34316),
            .I(N__34235));
    InMux I__6624 (
            .O(N__34315),
            .I(N__34235));
    InMux I__6623 (
            .O(N__34314),
            .I(N__34232));
    InMux I__6622 (
            .O(N__34313),
            .I(N__34229));
    InMux I__6621 (
            .O(N__34312),
            .I(N__34226));
    InMux I__6620 (
            .O(N__34311),
            .I(N__34222));
    LocalMux I__6619 (
            .O(N__34308),
            .I(N__34219));
    LocalMux I__6618 (
            .O(N__34303),
            .I(N__34216));
    LocalMux I__6617 (
            .O(N__34300),
            .I(N__34209));
    LocalMux I__6616 (
            .O(N__34297),
            .I(N__34204));
    LocalMux I__6615 (
            .O(N__34290),
            .I(N__34204));
    InMux I__6614 (
            .O(N__34289),
            .I(N__34199));
    InMux I__6613 (
            .O(N__34288),
            .I(N__34199));
    CascadeMux I__6612 (
            .O(N__34287),
            .I(N__34187));
    CascadeMux I__6611 (
            .O(N__34286),
            .I(N__34184));
    InMux I__6610 (
            .O(N__34285),
            .I(N__34169));
    InMux I__6609 (
            .O(N__34284),
            .I(N__34169));
    InMux I__6608 (
            .O(N__34283),
            .I(N__34169));
    InMux I__6607 (
            .O(N__34282),
            .I(N__34166));
    LocalMux I__6606 (
            .O(N__34279),
            .I(N__34161));
    LocalMux I__6605 (
            .O(N__34274),
            .I(N__34161));
    LocalMux I__6604 (
            .O(N__34269),
            .I(N__34154));
    LocalMux I__6603 (
            .O(N__34262),
            .I(N__34154));
    LocalMux I__6602 (
            .O(N__34249),
            .I(N__34154));
    InMux I__6601 (
            .O(N__34248),
            .I(N__34145));
    InMux I__6600 (
            .O(N__34247),
            .I(N__34145));
    InMux I__6599 (
            .O(N__34246),
            .I(N__34145));
    InMux I__6598 (
            .O(N__34245),
            .I(N__34145));
    InMux I__6597 (
            .O(N__34244),
            .I(N__34134));
    InMux I__6596 (
            .O(N__34243),
            .I(N__34134));
    InMux I__6595 (
            .O(N__34242),
            .I(N__34134));
    InMux I__6594 (
            .O(N__34241),
            .I(N__34134));
    InMux I__6593 (
            .O(N__34240),
            .I(N__34134));
    LocalMux I__6592 (
            .O(N__34235),
            .I(N__34127));
    LocalMux I__6591 (
            .O(N__34232),
            .I(N__34124));
    LocalMux I__6590 (
            .O(N__34229),
            .I(N__34119));
    LocalMux I__6589 (
            .O(N__34226),
            .I(N__34119));
    InMux I__6588 (
            .O(N__34225),
            .I(N__34116));
    LocalMux I__6587 (
            .O(N__34222),
            .I(N__34113));
    Span4Mux_v I__6586 (
            .O(N__34219),
            .I(N__34108));
    Span4Mux_v I__6585 (
            .O(N__34216),
            .I(N__34108));
    InMux I__6584 (
            .O(N__34215),
            .I(N__34099));
    InMux I__6583 (
            .O(N__34214),
            .I(N__34099));
    InMux I__6582 (
            .O(N__34213),
            .I(N__34099));
    InMux I__6581 (
            .O(N__34212),
            .I(N__34099));
    Span12Mux_h I__6580 (
            .O(N__34209),
            .I(N__34092));
    Sp12to4 I__6579 (
            .O(N__34204),
            .I(N__34092));
    LocalMux I__6578 (
            .O(N__34199),
            .I(N__34092));
    InMux I__6577 (
            .O(N__34198),
            .I(N__34087));
    InMux I__6576 (
            .O(N__34197),
            .I(N__34087));
    InMux I__6575 (
            .O(N__34196),
            .I(N__34076));
    InMux I__6574 (
            .O(N__34195),
            .I(N__34076));
    InMux I__6573 (
            .O(N__34194),
            .I(N__34076));
    InMux I__6572 (
            .O(N__34193),
            .I(N__34076));
    InMux I__6571 (
            .O(N__34192),
            .I(N__34076));
    InMux I__6570 (
            .O(N__34191),
            .I(N__34059));
    InMux I__6569 (
            .O(N__34190),
            .I(N__34059));
    InMux I__6568 (
            .O(N__34187),
            .I(N__34059));
    InMux I__6567 (
            .O(N__34184),
            .I(N__34059));
    InMux I__6566 (
            .O(N__34183),
            .I(N__34059));
    InMux I__6565 (
            .O(N__34182),
            .I(N__34059));
    InMux I__6564 (
            .O(N__34181),
            .I(N__34059));
    InMux I__6563 (
            .O(N__34180),
            .I(N__34059));
    InMux I__6562 (
            .O(N__34179),
            .I(N__34054));
    InMux I__6561 (
            .O(N__34178),
            .I(N__34054));
    InMux I__6560 (
            .O(N__34177),
            .I(N__34049));
    InMux I__6559 (
            .O(N__34176),
            .I(N__34049));
    LocalMux I__6558 (
            .O(N__34169),
            .I(N__34042));
    LocalMux I__6557 (
            .O(N__34166),
            .I(N__34042));
    Span4Mux_h I__6556 (
            .O(N__34161),
            .I(N__34042));
    Span4Mux_v I__6555 (
            .O(N__34154),
            .I(N__34035));
    LocalMux I__6554 (
            .O(N__34145),
            .I(N__34035));
    LocalMux I__6553 (
            .O(N__34134),
            .I(N__34035));
    InMux I__6552 (
            .O(N__34133),
            .I(N__34026));
    InMux I__6551 (
            .O(N__34132),
            .I(N__34026));
    InMux I__6550 (
            .O(N__34131),
            .I(N__34026));
    InMux I__6549 (
            .O(N__34130),
            .I(N__34026));
    Span4Mux_v I__6548 (
            .O(N__34127),
            .I(N__34017));
    Span4Mux_v I__6547 (
            .O(N__34124),
            .I(N__34017));
    Span4Mux_v I__6546 (
            .O(N__34119),
            .I(N__34017));
    LocalMux I__6545 (
            .O(N__34116),
            .I(N__34017));
    Odrv12 I__6544 (
            .O(N__34113),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6543 (
            .O(N__34108),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6542 (
            .O(N__34099),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv12 I__6541 (
            .O(N__34092),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6540 (
            .O(N__34087),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6539 (
            .O(N__34076),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6538 (
            .O(N__34059),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6537 (
            .O(N__34054),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6536 (
            .O(N__34049),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6535 (
            .O(N__34042),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6534 (
            .O(N__34035),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__6533 (
            .O(N__34026),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__6532 (
            .O(N__34017),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    CascadeMux I__6531 (
            .O(N__33990),
            .I(N__33972));
    CascadeMux I__6530 (
            .O(N__33989),
            .I(N__33964));
    InMux I__6529 (
            .O(N__33988),
            .I(N__33954));
    InMux I__6528 (
            .O(N__33987),
            .I(N__33954));
    CascadeMux I__6527 (
            .O(N__33986),
            .I(N__33949));
    CascadeMux I__6526 (
            .O(N__33985),
            .I(N__33942));
    CascadeMux I__6525 (
            .O(N__33984),
            .I(N__33938));
    CascadeMux I__6524 (
            .O(N__33983),
            .I(N__33932));
    CascadeMux I__6523 (
            .O(N__33982),
            .I(N__33928));
    CascadeMux I__6522 (
            .O(N__33981),
            .I(N__33924));
    CascadeMux I__6521 (
            .O(N__33980),
            .I(N__33921));
    CascadeMux I__6520 (
            .O(N__33979),
            .I(N__33917));
    CascadeMux I__6519 (
            .O(N__33978),
            .I(N__33912));
    CascadeMux I__6518 (
            .O(N__33977),
            .I(N__33908));
    CascadeMux I__6517 (
            .O(N__33976),
            .I(N__33905));
    InMux I__6516 (
            .O(N__33975),
            .I(N__33902));
    InMux I__6515 (
            .O(N__33972),
            .I(N__33899));
    CascadeMux I__6514 (
            .O(N__33971),
            .I(N__33892));
    CascadeMux I__6513 (
            .O(N__33970),
            .I(N__33889));
    CascadeMux I__6512 (
            .O(N__33969),
            .I(N__33884));
    CascadeMux I__6511 (
            .O(N__33968),
            .I(N__33880));
    CascadeMux I__6510 (
            .O(N__33967),
            .I(N__33876));
    InMux I__6509 (
            .O(N__33964),
            .I(N__33860));
    CascadeMux I__6508 (
            .O(N__33963),
            .I(N__33856));
    InMux I__6507 (
            .O(N__33962),
            .I(N__33846));
    InMux I__6506 (
            .O(N__33961),
            .I(N__33846));
    InMux I__6505 (
            .O(N__33960),
            .I(N__33846));
    InMux I__6504 (
            .O(N__33959),
            .I(N__33846));
    LocalMux I__6503 (
            .O(N__33954),
            .I(N__33843));
    InMux I__6502 (
            .O(N__33953),
            .I(N__33838));
    InMux I__6501 (
            .O(N__33952),
            .I(N__33838));
    InMux I__6500 (
            .O(N__33949),
            .I(N__33835));
    InMux I__6499 (
            .O(N__33948),
            .I(N__33828));
    InMux I__6498 (
            .O(N__33947),
            .I(N__33828));
    InMux I__6497 (
            .O(N__33946),
            .I(N__33828));
    InMux I__6496 (
            .O(N__33945),
            .I(N__33825));
    InMux I__6495 (
            .O(N__33942),
            .I(N__33814));
    InMux I__6494 (
            .O(N__33941),
            .I(N__33814));
    InMux I__6493 (
            .O(N__33938),
            .I(N__33814));
    InMux I__6492 (
            .O(N__33937),
            .I(N__33814));
    InMux I__6491 (
            .O(N__33936),
            .I(N__33814));
    InMux I__6490 (
            .O(N__33935),
            .I(N__33805));
    InMux I__6489 (
            .O(N__33932),
            .I(N__33805));
    InMux I__6488 (
            .O(N__33931),
            .I(N__33805));
    InMux I__6487 (
            .O(N__33928),
            .I(N__33805));
    InMux I__6486 (
            .O(N__33927),
            .I(N__33794));
    InMux I__6485 (
            .O(N__33924),
            .I(N__33794));
    InMux I__6484 (
            .O(N__33921),
            .I(N__33794));
    InMux I__6483 (
            .O(N__33920),
            .I(N__33794));
    InMux I__6482 (
            .O(N__33917),
            .I(N__33794));
    CascadeMux I__6481 (
            .O(N__33916),
            .I(N__33790));
    InMux I__6480 (
            .O(N__33915),
            .I(N__33774));
    InMux I__6479 (
            .O(N__33912),
            .I(N__33774));
    InMux I__6478 (
            .O(N__33911),
            .I(N__33774));
    InMux I__6477 (
            .O(N__33908),
            .I(N__33769));
    InMux I__6476 (
            .O(N__33905),
            .I(N__33769));
    LocalMux I__6475 (
            .O(N__33902),
            .I(N__33766));
    LocalMux I__6474 (
            .O(N__33899),
            .I(N__33759));
    CascadeMux I__6473 (
            .O(N__33898),
            .I(N__33755));
    CascadeMux I__6472 (
            .O(N__33897),
            .I(N__33751));
    CascadeMux I__6471 (
            .O(N__33896),
            .I(N__33747));
    InMux I__6470 (
            .O(N__33895),
            .I(N__33739));
    InMux I__6469 (
            .O(N__33892),
            .I(N__33739));
    InMux I__6468 (
            .O(N__33889),
            .I(N__33739));
    InMux I__6467 (
            .O(N__33888),
            .I(N__33722));
    InMux I__6466 (
            .O(N__33887),
            .I(N__33722));
    InMux I__6465 (
            .O(N__33884),
            .I(N__33722));
    InMux I__6464 (
            .O(N__33883),
            .I(N__33722));
    InMux I__6463 (
            .O(N__33880),
            .I(N__33722));
    InMux I__6462 (
            .O(N__33879),
            .I(N__33722));
    InMux I__6461 (
            .O(N__33876),
            .I(N__33722));
    InMux I__6460 (
            .O(N__33875),
            .I(N__33722));
    CascadeMux I__6459 (
            .O(N__33874),
            .I(N__33719));
    CascadeMux I__6458 (
            .O(N__33873),
            .I(N__33715));
    CascadeMux I__6457 (
            .O(N__33872),
            .I(N__33711));
    CascadeMux I__6456 (
            .O(N__33871),
            .I(N__33707));
    CascadeMux I__6455 (
            .O(N__33870),
            .I(N__33703));
    CascadeMux I__6454 (
            .O(N__33869),
            .I(N__33699));
    CascadeMux I__6453 (
            .O(N__33868),
            .I(N__33695));
    CascadeMux I__6452 (
            .O(N__33867),
            .I(N__33691));
    CascadeMux I__6451 (
            .O(N__33866),
            .I(N__33687));
    CascadeMux I__6450 (
            .O(N__33865),
            .I(N__33683));
    CascadeMux I__6449 (
            .O(N__33864),
            .I(N__33679));
    CascadeMux I__6448 (
            .O(N__33863),
            .I(N__33675));
    LocalMux I__6447 (
            .O(N__33860),
            .I(N__33667));
    InMux I__6446 (
            .O(N__33859),
            .I(N__33662));
    InMux I__6445 (
            .O(N__33856),
            .I(N__33662));
    CascadeMux I__6444 (
            .O(N__33855),
            .I(N__33658));
    LocalMux I__6443 (
            .O(N__33846),
            .I(N__33655));
    Span4Mux_h I__6442 (
            .O(N__33843),
            .I(N__33650));
    LocalMux I__6441 (
            .O(N__33838),
            .I(N__33650));
    LocalMux I__6440 (
            .O(N__33835),
            .I(N__33639));
    LocalMux I__6439 (
            .O(N__33828),
            .I(N__33639));
    LocalMux I__6438 (
            .O(N__33825),
            .I(N__33639));
    LocalMux I__6437 (
            .O(N__33814),
            .I(N__33639));
    LocalMux I__6436 (
            .O(N__33805),
            .I(N__33639));
    LocalMux I__6435 (
            .O(N__33794),
            .I(N__33636));
    InMux I__6434 (
            .O(N__33793),
            .I(N__33633));
    InMux I__6433 (
            .O(N__33790),
            .I(N__33630));
    CascadeMux I__6432 (
            .O(N__33789),
            .I(N__33623));
    CascadeMux I__6431 (
            .O(N__33788),
            .I(N__33618));
    InMux I__6430 (
            .O(N__33787),
            .I(N__33611));
    InMux I__6429 (
            .O(N__33786),
            .I(N__33611));
    InMux I__6428 (
            .O(N__33785),
            .I(N__33611));
    InMux I__6427 (
            .O(N__33784),
            .I(N__33606));
    InMux I__6426 (
            .O(N__33783),
            .I(N__33606));
    InMux I__6425 (
            .O(N__33782),
            .I(N__33601));
    InMux I__6424 (
            .O(N__33781),
            .I(N__33601));
    LocalMux I__6423 (
            .O(N__33774),
            .I(N__33594));
    LocalMux I__6422 (
            .O(N__33769),
            .I(N__33594));
    Span4Mux_v I__6421 (
            .O(N__33766),
            .I(N__33594));
    CascadeMux I__6420 (
            .O(N__33765),
            .I(N__33590));
    CascadeMux I__6419 (
            .O(N__33764),
            .I(N__33586));
    CascadeMux I__6418 (
            .O(N__33763),
            .I(N__33582));
    CascadeMux I__6417 (
            .O(N__33762),
            .I(N__33578));
    Span4Mux_h I__6416 (
            .O(N__33759),
            .I(N__33575));
    InMux I__6415 (
            .O(N__33758),
            .I(N__33560));
    InMux I__6414 (
            .O(N__33755),
            .I(N__33560));
    InMux I__6413 (
            .O(N__33754),
            .I(N__33560));
    InMux I__6412 (
            .O(N__33751),
            .I(N__33560));
    InMux I__6411 (
            .O(N__33750),
            .I(N__33560));
    InMux I__6410 (
            .O(N__33747),
            .I(N__33560));
    InMux I__6409 (
            .O(N__33746),
            .I(N__33560));
    LocalMux I__6408 (
            .O(N__33739),
            .I(N__33555));
    LocalMux I__6407 (
            .O(N__33722),
            .I(N__33555));
    InMux I__6406 (
            .O(N__33719),
            .I(N__33538));
    InMux I__6405 (
            .O(N__33718),
            .I(N__33538));
    InMux I__6404 (
            .O(N__33715),
            .I(N__33538));
    InMux I__6403 (
            .O(N__33714),
            .I(N__33538));
    InMux I__6402 (
            .O(N__33711),
            .I(N__33538));
    InMux I__6401 (
            .O(N__33710),
            .I(N__33538));
    InMux I__6400 (
            .O(N__33707),
            .I(N__33538));
    InMux I__6399 (
            .O(N__33706),
            .I(N__33538));
    InMux I__6398 (
            .O(N__33703),
            .I(N__33521));
    InMux I__6397 (
            .O(N__33702),
            .I(N__33521));
    InMux I__6396 (
            .O(N__33699),
            .I(N__33521));
    InMux I__6395 (
            .O(N__33698),
            .I(N__33521));
    InMux I__6394 (
            .O(N__33695),
            .I(N__33521));
    InMux I__6393 (
            .O(N__33694),
            .I(N__33521));
    InMux I__6392 (
            .O(N__33691),
            .I(N__33521));
    InMux I__6391 (
            .O(N__33690),
            .I(N__33521));
    InMux I__6390 (
            .O(N__33687),
            .I(N__33504));
    InMux I__6389 (
            .O(N__33686),
            .I(N__33504));
    InMux I__6388 (
            .O(N__33683),
            .I(N__33504));
    InMux I__6387 (
            .O(N__33682),
            .I(N__33504));
    InMux I__6386 (
            .O(N__33679),
            .I(N__33504));
    InMux I__6385 (
            .O(N__33678),
            .I(N__33504));
    InMux I__6384 (
            .O(N__33675),
            .I(N__33504));
    InMux I__6383 (
            .O(N__33674),
            .I(N__33504));
    CascadeMux I__6382 (
            .O(N__33673),
            .I(N__33499));
    CascadeMux I__6381 (
            .O(N__33672),
            .I(N__33495));
    CascadeMux I__6380 (
            .O(N__33671),
            .I(N__33491));
    CascadeMux I__6379 (
            .O(N__33670),
            .I(N__33485));
    Span4Mux_h I__6378 (
            .O(N__33667),
            .I(N__33479));
    LocalMux I__6377 (
            .O(N__33662),
            .I(N__33479));
    InMux I__6376 (
            .O(N__33661),
            .I(N__33474));
    InMux I__6375 (
            .O(N__33658),
            .I(N__33474));
    Span4Mux_v I__6374 (
            .O(N__33655),
            .I(N__33461));
    Span4Mux_v I__6373 (
            .O(N__33650),
            .I(N__33461));
    Span4Mux_v I__6372 (
            .O(N__33639),
            .I(N__33461));
    Span4Mux_v I__6371 (
            .O(N__33636),
            .I(N__33461));
    LocalMux I__6370 (
            .O(N__33633),
            .I(N__33461));
    LocalMux I__6369 (
            .O(N__33630),
            .I(N__33461));
    InMux I__6368 (
            .O(N__33629),
            .I(N__33444));
    InMux I__6367 (
            .O(N__33628),
            .I(N__33444));
    InMux I__6366 (
            .O(N__33627),
            .I(N__33444));
    InMux I__6365 (
            .O(N__33626),
            .I(N__33444));
    InMux I__6364 (
            .O(N__33623),
            .I(N__33444));
    InMux I__6363 (
            .O(N__33622),
            .I(N__33444));
    InMux I__6362 (
            .O(N__33621),
            .I(N__33444));
    InMux I__6361 (
            .O(N__33618),
            .I(N__33444));
    LocalMux I__6360 (
            .O(N__33611),
            .I(N__33435));
    LocalMux I__6359 (
            .O(N__33606),
            .I(N__33435));
    LocalMux I__6358 (
            .O(N__33601),
            .I(N__33435));
    Span4Mux_h I__6357 (
            .O(N__33594),
            .I(N__33435));
    InMux I__6356 (
            .O(N__33593),
            .I(N__33418));
    InMux I__6355 (
            .O(N__33590),
            .I(N__33418));
    InMux I__6354 (
            .O(N__33589),
            .I(N__33418));
    InMux I__6353 (
            .O(N__33586),
            .I(N__33418));
    InMux I__6352 (
            .O(N__33585),
            .I(N__33418));
    InMux I__6351 (
            .O(N__33582),
            .I(N__33418));
    InMux I__6350 (
            .O(N__33581),
            .I(N__33418));
    InMux I__6349 (
            .O(N__33578),
            .I(N__33418));
    Span4Mux_h I__6348 (
            .O(N__33575),
            .I(N__33405));
    LocalMux I__6347 (
            .O(N__33560),
            .I(N__33405));
    Span4Mux_v I__6346 (
            .O(N__33555),
            .I(N__33405));
    LocalMux I__6345 (
            .O(N__33538),
            .I(N__33405));
    LocalMux I__6344 (
            .O(N__33521),
            .I(N__33405));
    LocalMux I__6343 (
            .O(N__33504),
            .I(N__33405));
    InMux I__6342 (
            .O(N__33503),
            .I(N__33400));
    InMux I__6341 (
            .O(N__33502),
            .I(N__33400));
    InMux I__6340 (
            .O(N__33499),
            .I(N__33387));
    InMux I__6339 (
            .O(N__33498),
            .I(N__33387));
    InMux I__6338 (
            .O(N__33495),
            .I(N__33387));
    InMux I__6337 (
            .O(N__33494),
            .I(N__33387));
    InMux I__6336 (
            .O(N__33491),
            .I(N__33387));
    InMux I__6335 (
            .O(N__33490),
            .I(N__33387));
    InMux I__6334 (
            .O(N__33489),
            .I(N__33378));
    InMux I__6333 (
            .O(N__33488),
            .I(N__33378));
    InMux I__6332 (
            .O(N__33485),
            .I(N__33378));
    InMux I__6331 (
            .O(N__33484),
            .I(N__33378));
    Odrv4 I__6330 (
            .O(N__33479),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6329 (
            .O(N__33474),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6328 (
            .O(N__33461),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6327 (
            .O(N__33444),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6326 (
            .O(N__33435),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6325 (
            .O(N__33418),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__6324 (
            .O(N__33405),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6323 (
            .O(N__33400),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6322 (
            .O(N__33387),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__6321 (
            .O(N__33378),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    CascadeMux I__6320 (
            .O(N__33357),
            .I(N__33354));
    InMux I__6319 (
            .O(N__33354),
            .I(N__33351));
    LocalMux I__6318 (
            .O(N__33351),
            .I(N__33347));
    InMux I__6317 (
            .O(N__33350),
            .I(N__33344));
    Span4Mux_h I__6316 (
            .O(N__33347),
            .I(N__33340));
    LocalMux I__6315 (
            .O(N__33344),
            .I(N__33337));
    InMux I__6314 (
            .O(N__33343),
            .I(N__33334));
    Sp12to4 I__6313 (
            .O(N__33340),
            .I(N__33331));
    Span4Mux_h I__6312 (
            .O(N__33337),
            .I(N__33328));
    LocalMux I__6311 (
            .O(N__33334),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv12 I__6310 (
            .O(N__33331),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__6309 (
            .O(N__33328),
            .I(\current_shift_inst.un4_control_input1_25 ));
    CascadeMux I__6308 (
            .O(N__33321),
            .I(N__33318));
    InMux I__6307 (
            .O(N__33318),
            .I(N__33315));
    LocalMux I__6306 (
            .O(N__33315),
            .I(N__33312));
    Span4Mux_h I__6305 (
            .O(N__33312),
            .I(N__33309));
    Span4Mux_v I__6304 (
            .O(N__33309),
            .I(N__33306));
    Odrv4 I__6303 (
            .O(N__33306),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__6302 (
            .O(N__33303),
            .I(N__33300));
    LocalMux I__6301 (
            .O(N__33300),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__6300 (
            .O(N__33297),
            .I(N__33294));
    LocalMux I__6299 (
            .O(N__33294),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    InMux I__6298 (
            .O(N__33291),
            .I(N__33288));
    LocalMux I__6297 (
            .O(N__33288),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__6296 (
            .O(N__33285),
            .I(N__33281));
    InMux I__6295 (
            .O(N__33284),
            .I(N__33278));
    LocalMux I__6294 (
            .O(N__33281),
            .I(N__33273));
    LocalMux I__6293 (
            .O(N__33278),
            .I(N__33273));
    Span4Mux_h I__6292 (
            .O(N__33273),
            .I(N__33270));
    Span4Mux_v I__6291 (
            .O(N__33270),
            .I(N__33266));
    InMux I__6290 (
            .O(N__33269),
            .I(N__33263));
    Odrv4 I__6289 (
            .O(N__33266),
            .I(\current_shift_inst.un4_control_input1_21 ));
    LocalMux I__6288 (
            .O(N__33263),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__6287 (
            .O(N__33258),
            .I(N__33255));
    LocalMux I__6286 (
            .O(N__33255),
            .I(N__33252));
    Span4Mux_h I__6285 (
            .O(N__33252),
            .I(N__33249));
    Odrv4 I__6284 (
            .O(N__33249),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__6283 (
            .O(N__33246),
            .I(N__33243));
    LocalMux I__6282 (
            .O(N__33243),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__6281 (
            .O(N__33240),
            .I(N__33237));
    LocalMux I__6280 (
            .O(N__33237),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__6279 (
            .O(N__33234),
            .I(N__33229));
    InMux I__6278 (
            .O(N__33233),
            .I(N__33226));
    InMux I__6277 (
            .O(N__33232),
            .I(N__33223));
    InMux I__6276 (
            .O(N__33229),
            .I(N__33220));
    LocalMux I__6275 (
            .O(N__33226),
            .I(\current_shift_inst.N_1275_i ));
    LocalMux I__6274 (
            .O(N__33223),
            .I(\current_shift_inst.N_1275_i ));
    LocalMux I__6273 (
            .O(N__33220),
            .I(\current_shift_inst.N_1275_i ));
    InMux I__6272 (
            .O(N__33213),
            .I(N__33210));
    LocalMux I__6271 (
            .O(N__33210),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__6270 (
            .O(N__33207),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__6269 (
            .O(N__33204),
            .I(N__33201));
    LocalMux I__6268 (
            .O(N__33201),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__6267 (
            .O(N__33198),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__6266 (
            .O(N__33195),
            .I(N__33192));
    LocalMux I__6265 (
            .O(N__33192),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__6264 (
            .O(N__33189),
            .I(N__33186));
    LocalMux I__6263 (
            .O(N__33186),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    CascadeMux I__6262 (
            .O(N__33183),
            .I(N__33180));
    InMux I__6261 (
            .O(N__33180),
            .I(N__33177));
    LocalMux I__6260 (
            .O(N__33177),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__6259 (
            .O(N__33174),
            .I(N__33171));
    LocalMux I__6258 (
            .O(N__33171),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__6257 (
            .O(N__33168),
            .I(N__33165));
    LocalMux I__6256 (
            .O(N__33165),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__6255 (
            .O(N__33162),
            .I(N__33159));
    LocalMux I__6254 (
            .O(N__33159),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__6253 (
            .O(N__33156),
            .I(N__33153));
    LocalMux I__6252 (
            .O(N__33153),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__6251 (
            .O(N__33150),
            .I(N__33147));
    LocalMux I__6250 (
            .O(N__33147),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__6249 (
            .O(N__33144),
            .I(N__33141));
    LocalMux I__6248 (
            .O(N__33141),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__6247 (
            .O(N__33138),
            .I(N__33134));
    InMux I__6246 (
            .O(N__33137),
            .I(N__33131));
    LocalMux I__6245 (
            .O(N__33134),
            .I(N__33127));
    LocalMux I__6244 (
            .O(N__33131),
            .I(N__33124));
    InMux I__6243 (
            .O(N__33130),
            .I(N__33121));
    Odrv12 I__6242 (
            .O(N__33127),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__6241 (
            .O(N__33124),
            .I(\current_shift_inst.un4_control_input1_20 ));
    LocalMux I__6240 (
            .O(N__33121),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__6239 (
            .O(N__33114),
            .I(N__33111));
    InMux I__6238 (
            .O(N__33111),
            .I(N__33108));
    LocalMux I__6237 (
            .O(N__33108),
            .I(N__33105));
    Span4Mux_v I__6236 (
            .O(N__33105),
            .I(N__33102));
    Odrv4 I__6235 (
            .O(N__33102),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__6234 (
            .O(N__33099),
            .I(N__33096));
    LocalMux I__6233 (
            .O(N__33096),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__6232 (
            .O(N__33093),
            .I(N__33090));
    LocalMux I__6231 (
            .O(N__33090),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__6230 (
            .O(N__33087),
            .I(N__33084));
    LocalMux I__6229 (
            .O(N__33084),
            .I(N__33080));
    InMux I__6228 (
            .O(N__33083),
            .I(N__33077));
    Span12Mux_h I__6227 (
            .O(N__33080),
            .I(N__33073));
    LocalMux I__6226 (
            .O(N__33077),
            .I(N__33070));
    InMux I__6225 (
            .O(N__33076),
            .I(N__33067));
    Odrv12 I__6224 (
            .O(N__33073),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__6223 (
            .O(N__33070),
            .I(\current_shift_inst.un4_control_input1_22 ));
    LocalMux I__6222 (
            .O(N__33067),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__6221 (
            .O(N__33060),
            .I(N__33057));
    InMux I__6220 (
            .O(N__33057),
            .I(N__33054));
    LocalMux I__6219 (
            .O(N__33054),
            .I(N__33051));
    Span4Mux_v I__6218 (
            .O(N__33051),
            .I(N__33048));
    Odrv4 I__6217 (
            .O(N__33048),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    InMux I__6216 (
            .O(N__33045),
            .I(N__33042));
    LocalMux I__6215 (
            .O(N__33042),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__6214 (
            .O(N__33039),
            .I(N__33036));
    LocalMux I__6213 (
            .O(N__33036),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    CascadeMux I__6212 (
            .O(N__33033),
            .I(N__33030));
    InMux I__6211 (
            .O(N__33030),
            .I(N__33027));
    LocalMux I__6210 (
            .O(N__33027),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__6209 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__6208 (
            .O(N__33021),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__6207 (
            .O(N__33018),
            .I(N__33014));
    InMux I__6206 (
            .O(N__33017),
            .I(N__33011));
    LocalMux I__6205 (
            .O(N__33014),
            .I(N__33006));
    LocalMux I__6204 (
            .O(N__33011),
            .I(N__33006));
    Span4Mux_h I__6203 (
            .O(N__33006),
            .I(N__33003));
    Span4Mux_v I__6202 (
            .O(N__33003),
            .I(N__32998));
    InMux I__6201 (
            .O(N__33002),
            .I(N__32993));
    InMux I__6200 (
            .O(N__33001),
            .I(N__32993));
    Odrv4 I__6199 (
            .O(N__32998),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__6198 (
            .O(N__32993),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    InMux I__6197 (
            .O(N__32988),
            .I(N__32985));
    LocalMux I__6196 (
            .O(N__32985),
            .I(N__32982));
    Span4Mux_h I__6195 (
            .O(N__32982),
            .I(N__32978));
    InMux I__6194 (
            .O(N__32981),
            .I(N__32975));
    Span4Mux_v I__6193 (
            .O(N__32978),
            .I(N__32972));
    LocalMux I__6192 (
            .O(N__32975),
            .I(N__32969));
    Span4Mux_h I__6191 (
            .O(N__32972),
            .I(N__32965));
    Span4Mux_h I__6190 (
            .O(N__32969),
            .I(N__32962));
    InMux I__6189 (
            .O(N__32968),
            .I(N__32959));
    Odrv4 I__6188 (
            .O(N__32965),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__6187 (
            .O(N__32962),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__6186 (
            .O(N__32959),
            .I(\current_shift_inst.un4_control_input1_4 ));
    CascadeMux I__6185 (
            .O(N__32952),
            .I(N__32949));
    InMux I__6184 (
            .O(N__32949),
            .I(N__32946));
    LocalMux I__6183 (
            .O(N__32946),
            .I(N__32943));
    Span4Mux_v I__6182 (
            .O(N__32943),
            .I(N__32940));
    Odrv4 I__6181 (
            .O(N__32940),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__6180 (
            .O(N__32937),
            .I(N__32934));
    LocalMux I__6179 (
            .O(N__32934),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__6178 (
            .O(N__32931),
            .I(N__32928));
    LocalMux I__6177 (
            .O(N__32928),
            .I(N__32925));
    Span4Mux_h I__6176 (
            .O(N__32925),
            .I(N__32921));
    InMux I__6175 (
            .O(N__32924),
            .I(N__32918));
    Span4Mux_v I__6174 (
            .O(N__32921),
            .I(N__32914));
    LocalMux I__6173 (
            .O(N__32918),
            .I(N__32911));
    InMux I__6172 (
            .O(N__32917),
            .I(N__32908));
    Odrv4 I__6171 (
            .O(N__32914),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__6170 (
            .O(N__32911),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__6169 (
            .O(N__32908),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__6168 (
            .O(N__32901),
            .I(N__32898));
    LocalMux I__6167 (
            .O(N__32898),
            .I(N__32895));
    Span4Mux_h I__6166 (
            .O(N__32895),
            .I(N__32892));
    Odrv4 I__6165 (
            .O(N__32892),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    InMux I__6164 (
            .O(N__32889),
            .I(N__32886));
    LocalMux I__6163 (
            .O(N__32886),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    CascadeMux I__6162 (
            .O(N__32883),
            .I(N__32880));
    InMux I__6161 (
            .O(N__32880),
            .I(N__32877));
    LocalMux I__6160 (
            .O(N__32877),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__6159 (
            .O(N__32874),
            .I(N__32871));
    LocalMux I__6158 (
            .O(N__32871),
            .I(N__32868));
    Span12Mux_v I__6157 (
            .O(N__32868),
            .I(N__32865));
    Odrv12 I__6156 (
            .O(N__32865),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__6155 (
            .O(N__32862),
            .I(N__32859));
    LocalMux I__6154 (
            .O(N__32859),
            .I(N__32856));
    Span4Mux_v I__6153 (
            .O(N__32856),
            .I(N__32853));
    Span4Mux_h I__6152 (
            .O(N__32853),
            .I(N__32850));
    Odrv4 I__6151 (
            .O(N__32850),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__6150 (
            .O(N__32847),
            .I(N__32844));
    LocalMux I__6149 (
            .O(N__32844),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__6148 (
            .O(N__32841),
            .I(N__32838));
    LocalMux I__6147 (
            .O(N__32838),
            .I(N__32834));
    InMux I__6146 (
            .O(N__32837),
            .I(N__32831));
    Odrv4 I__6145 (
            .O(N__32834),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    LocalMux I__6144 (
            .O(N__32831),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    CascadeMux I__6143 (
            .O(N__32826),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_));
    InMux I__6142 (
            .O(N__32823),
            .I(N__32816));
    InMux I__6141 (
            .O(N__32822),
            .I(N__32816));
    InMux I__6140 (
            .O(N__32821),
            .I(N__32813));
    LocalMux I__6139 (
            .O(N__32816),
            .I(N__32809));
    LocalMux I__6138 (
            .O(N__32813),
            .I(N__32806));
    InMux I__6137 (
            .O(N__32812),
            .I(N__32803));
    Span4Mux_v I__6136 (
            .O(N__32809),
            .I(N__32800));
    Span4Mux_h I__6135 (
            .O(N__32806),
            .I(N__32795));
    LocalMux I__6134 (
            .O(N__32803),
            .I(N__32795));
    Span4Mux_h I__6133 (
            .O(N__32800),
            .I(N__32792));
    Span4Mux_h I__6132 (
            .O(N__32795),
            .I(N__32789));
    Odrv4 I__6131 (
            .O(N__32792),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    Odrv4 I__6130 (
            .O(N__32789),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    CascadeMux I__6129 (
            .O(N__32784),
            .I(N__32781));
    InMux I__6128 (
            .O(N__32781),
            .I(N__32775));
    InMux I__6127 (
            .O(N__32780),
            .I(N__32775));
    LocalMux I__6126 (
            .O(N__32775),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ));
    InMux I__6125 (
            .O(N__32772),
            .I(N__32769));
    LocalMux I__6124 (
            .O(N__32769),
            .I(N__32764));
    InMux I__6123 (
            .O(N__32768),
            .I(N__32761));
    InMux I__6122 (
            .O(N__32767),
            .I(N__32758));
    Span4Mux_v I__6121 (
            .O(N__32764),
            .I(N__32753));
    LocalMux I__6120 (
            .O(N__32761),
            .I(N__32753));
    LocalMux I__6119 (
            .O(N__32758),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    Odrv4 I__6118 (
            .O(N__32753),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__6117 (
            .O(N__32748),
            .I(N__32742));
    CascadeMux I__6116 (
            .O(N__32747),
            .I(N__32739));
    InMux I__6115 (
            .O(N__32746),
            .I(N__32736));
    InMux I__6114 (
            .O(N__32745),
            .I(N__32733));
    LocalMux I__6113 (
            .O(N__32742),
            .I(N__32730));
    InMux I__6112 (
            .O(N__32739),
            .I(N__32727));
    LocalMux I__6111 (
            .O(N__32736),
            .I(N__32724));
    LocalMux I__6110 (
            .O(N__32733),
            .I(N__32717));
    Span4Mux_h I__6109 (
            .O(N__32730),
            .I(N__32717));
    LocalMux I__6108 (
            .O(N__32727),
            .I(N__32717));
    Span4Mux_h I__6107 (
            .O(N__32724),
            .I(N__32714));
    Span4Mux_h I__6106 (
            .O(N__32717),
            .I(N__32711));
    Odrv4 I__6105 (
            .O(N__32714),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    Odrv4 I__6104 (
            .O(N__32711),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    InMux I__6103 (
            .O(N__32706),
            .I(N__32703));
    LocalMux I__6102 (
            .O(N__32703),
            .I(N__32700));
    Span4Mux_h I__6101 (
            .O(N__32700),
            .I(N__32697));
    Odrv4 I__6100 (
            .O(N__32697),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__6099 (
            .O(N__32694),
            .I(N__32645));
    InMux I__6098 (
            .O(N__32693),
            .I(N__32641));
    InMux I__6097 (
            .O(N__32692),
            .I(N__32634));
    InMux I__6096 (
            .O(N__32691),
            .I(N__32634));
    InMux I__6095 (
            .O(N__32690),
            .I(N__32627));
    InMux I__6094 (
            .O(N__32689),
            .I(N__32627));
    InMux I__6093 (
            .O(N__32688),
            .I(N__32627));
    InMux I__6092 (
            .O(N__32687),
            .I(N__32613));
    InMux I__6091 (
            .O(N__32686),
            .I(N__32613));
    InMux I__6090 (
            .O(N__32685),
            .I(N__32613));
    InMux I__6089 (
            .O(N__32684),
            .I(N__32613));
    InMux I__6088 (
            .O(N__32683),
            .I(N__32596));
    InMux I__6087 (
            .O(N__32682),
            .I(N__32596));
    InMux I__6086 (
            .O(N__32681),
            .I(N__32596));
    InMux I__6085 (
            .O(N__32680),
            .I(N__32589));
    InMux I__6084 (
            .O(N__32679),
            .I(N__32589));
    InMux I__6083 (
            .O(N__32678),
            .I(N__32589));
    InMux I__6082 (
            .O(N__32677),
            .I(N__32578));
    InMux I__6081 (
            .O(N__32676),
            .I(N__32578));
    InMux I__6080 (
            .O(N__32675),
            .I(N__32578));
    InMux I__6079 (
            .O(N__32674),
            .I(N__32578));
    InMux I__6078 (
            .O(N__32673),
            .I(N__32578));
    InMux I__6077 (
            .O(N__32672),
            .I(N__32571));
    InMux I__6076 (
            .O(N__32671),
            .I(N__32571));
    InMux I__6075 (
            .O(N__32670),
            .I(N__32571));
    InMux I__6074 (
            .O(N__32669),
            .I(N__32566));
    InMux I__6073 (
            .O(N__32668),
            .I(N__32566));
    InMux I__6072 (
            .O(N__32667),
            .I(N__32558));
    InMux I__6071 (
            .O(N__32666),
            .I(N__32551));
    InMux I__6070 (
            .O(N__32665),
            .I(N__32551));
    InMux I__6069 (
            .O(N__32664),
            .I(N__32551));
    InMux I__6068 (
            .O(N__32663),
            .I(N__32542));
    InMux I__6067 (
            .O(N__32662),
            .I(N__32542));
    InMux I__6066 (
            .O(N__32661),
            .I(N__32542));
    InMux I__6065 (
            .O(N__32660),
            .I(N__32542));
    InMux I__6064 (
            .O(N__32659),
            .I(N__32539));
    InMux I__6063 (
            .O(N__32658),
            .I(N__32534));
    InMux I__6062 (
            .O(N__32657),
            .I(N__32534));
    InMux I__6061 (
            .O(N__32656),
            .I(N__32521));
    InMux I__6060 (
            .O(N__32655),
            .I(N__32521));
    InMux I__6059 (
            .O(N__32654),
            .I(N__32521));
    InMux I__6058 (
            .O(N__32653),
            .I(N__32521));
    InMux I__6057 (
            .O(N__32652),
            .I(N__32521));
    InMux I__6056 (
            .O(N__32651),
            .I(N__32521));
    InMux I__6055 (
            .O(N__32650),
            .I(N__32510));
    InMux I__6054 (
            .O(N__32649),
            .I(N__32510));
    InMux I__6053 (
            .O(N__32648),
            .I(N__32510));
    InMux I__6052 (
            .O(N__32645),
            .I(N__32510));
    InMux I__6051 (
            .O(N__32644),
            .I(N__32510));
    LocalMux I__6050 (
            .O(N__32641),
            .I(N__32507));
    InMux I__6049 (
            .O(N__32640),
            .I(N__32504));
    InMux I__6048 (
            .O(N__32639),
            .I(N__32501));
    LocalMux I__6047 (
            .O(N__32634),
            .I(N__32498));
    LocalMux I__6046 (
            .O(N__32627),
            .I(N__32495));
    InMux I__6045 (
            .O(N__32626),
            .I(N__32478));
    InMux I__6044 (
            .O(N__32625),
            .I(N__32478));
    InMux I__6043 (
            .O(N__32624),
            .I(N__32478));
    InMux I__6042 (
            .O(N__32623),
            .I(N__32473));
    InMux I__6041 (
            .O(N__32622),
            .I(N__32473));
    LocalMux I__6040 (
            .O(N__32613),
            .I(N__32470));
    InMux I__6039 (
            .O(N__32612),
            .I(N__32465));
    InMux I__6038 (
            .O(N__32611),
            .I(N__32465));
    InMux I__6037 (
            .O(N__32610),
            .I(N__32460));
    InMux I__6036 (
            .O(N__32609),
            .I(N__32460));
    InMux I__6035 (
            .O(N__32608),
            .I(N__32447));
    InMux I__6034 (
            .O(N__32607),
            .I(N__32447));
    InMux I__6033 (
            .O(N__32606),
            .I(N__32447));
    InMux I__6032 (
            .O(N__32605),
            .I(N__32447));
    InMux I__6031 (
            .O(N__32604),
            .I(N__32447));
    InMux I__6030 (
            .O(N__32603),
            .I(N__32447));
    LocalMux I__6029 (
            .O(N__32596),
            .I(N__32442));
    LocalMux I__6028 (
            .O(N__32589),
            .I(N__32442));
    LocalMux I__6027 (
            .O(N__32578),
            .I(N__32437));
    LocalMux I__6026 (
            .O(N__32571),
            .I(N__32437));
    LocalMux I__6025 (
            .O(N__32566),
            .I(N__32434));
    InMux I__6024 (
            .O(N__32565),
            .I(N__32427));
    InMux I__6023 (
            .O(N__32564),
            .I(N__32427));
    InMux I__6022 (
            .O(N__32563),
            .I(N__32422));
    InMux I__6021 (
            .O(N__32562),
            .I(N__32422));
    InMux I__6020 (
            .O(N__32561),
            .I(N__32419));
    LocalMux I__6019 (
            .O(N__32558),
            .I(N__32416));
    LocalMux I__6018 (
            .O(N__32551),
            .I(N__32411));
    LocalMux I__6017 (
            .O(N__32542),
            .I(N__32411));
    LocalMux I__6016 (
            .O(N__32539),
            .I(N__32400));
    LocalMux I__6015 (
            .O(N__32534),
            .I(N__32400));
    LocalMux I__6014 (
            .O(N__32521),
            .I(N__32400));
    LocalMux I__6013 (
            .O(N__32510),
            .I(N__32400));
    Span4Mux_v I__6012 (
            .O(N__32507),
            .I(N__32400));
    LocalMux I__6011 (
            .O(N__32504),
            .I(N__32391));
    LocalMux I__6010 (
            .O(N__32501),
            .I(N__32391));
    Span4Mux_v I__6009 (
            .O(N__32498),
            .I(N__32391));
    Span4Mux_v I__6008 (
            .O(N__32495),
            .I(N__32391));
    InMux I__6007 (
            .O(N__32494),
            .I(N__32377));
    InMux I__6006 (
            .O(N__32493),
            .I(N__32377));
    InMux I__6005 (
            .O(N__32492),
            .I(N__32374));
    InMux I__6004 (
            .O(N__32491),
            .I(N__32365));
    InMux I__6003 (
            .O(N__32490),
            .I(N__32365));
    InMux I__6002 (
            .O(N__32489),
            .I(N__32365));
    InMux I__6001 (
            .O(N__32488),
            .I(N__32365));
    InMux I__6000 (
            .O(N__32487),
            .I(N__32359));
    InMux I__5999 (
            .O(N__32486),
            .I(N__32359));
    InMux I__5998 (
            .O(N__32485),
            .I(N__32356));
    LocalMux I__5997 (
            .O(N__32478),
            .I(N__32353));
    LocalMux I__5996 (
            .O(N__32473),
            .I(N__32346));
    Span4Mux_h I__5995 (
            .O(N__32470),
            .I(N__32346));
    LocalMux I__5994 (
            .O(N__32465),
            .I(N__32346));
    LocalMux I__5993 (
            .O(N__32460),
            .I(N__32335));
    LocalMux I__5992 (
            .O(N__32447),
            .I(N__32335));
    Span4Mux_v I__5991 (
            .O(N__32442),
            .I(N__32335));
    Span4Mux_v I__5990 (
            .O(N__32437),
            .I(N__32335));
    Span4Mux_h I__5989 (
            .O(N__32434),
            .I(N__32335));
    InMux I__5988 (
            .O(N__32433),
            .I(N__32330));
    InMux I__5987 (
            .O(N__32432),
            .I(N__32330));
    LocalMux I__5986 (
            .O(N__32427),
            .I(N__32325));
    LocalMux I__5985 (
            .O(N__32422),
            .I(N__32325));
    LocalMux I__5984 (
            .O(N__32419),
            .I(N__32314));
    Span4Mux_v I__5983 (
            .O(N__32416),
            .I(N__32314));
    Span4Mux_v I__5982 (
            .O(N__32411),
            .I(N__32314));
    Span4Mux_v I__5981 (
            .O(N__32400),
            .I(N__32314));
    Span4Mux_h I__5980 (
            .O(N__32391),
            .I(N__32314));
    InMux I__5979 (
            .O(N__32390),
            .I(N__32303));
    InMux I__5978 (
            .O(N__32389),
            .I(N__32303));
    InMux I__5977 (
            .O(N__32388),
            .I(N__32303));
    InMux I__5976 (
            .O(N__32387),
            .I(N__32303));
    InMux I__5975 (
            .O(N__32386),
            .I(N__32303));
    InMux I__5974 (
            .O(N__32385),
            .I(N__32294));
    InMux I__5973 (
            .O(N__32384),
            .I(N__32294));
    InMux I__5972 (
            .O(N__32383),
            .I(N__32294));
    InMux I__5971 (
            .O(N__32382),
            .I(N__32294));
    LocalMux I__5970 (
            .O(N__32377),
            .I(N__32287));
    LocalMux I__5969 (
            .O(N__32374),
            .I(N__32287));
    LocalMux I__5968 (
            .O(N__32365),
            .I(N__32287));
    InMux I__5967 (
            .O(N__32364),
            .I(N__32284));
    LocalMux I__5966 (
            .O(N__32359),
            .I(N__32277));
    LocalMux I__5965 (
            .O(N__32356),
            .I(N__32277));
    Span12Mux_h I__5964 (
            .O(N__32353),
            .I(N__32277));
    Span4Mux_h I__5963 (
            .O(N__32346),
            .I(N__32272));
    Span4Mux_h I__5962 (
            .O(N__32335),
            .I(N__32272));
    LocalMux I__5961 (
            .O(N__32330),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__5960 (
            .O(N__32325),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5959 (
            .O(N__32314),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5958 (
            .O(N__32303),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5957 (
            .O(N__32294),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5956 (
            .O(N__32287),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5955 (
            .O(N__32284),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__5954 (
            .O(N__32277),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5953 (
            .O(N__32272),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__5952 (
            .O(N__32253),
            .I(N__32249));
    InMux I__5951 (
            .O(N__32252),
            .I(N__32245));
    LocalMux I__5950 (
            .O(N__32249),
            .I(N__32242));
    InMux I__5949 (
            .O(N__32248),
            .I(N__32239));
    LocalMux I__5948 (
            .O(N__32245),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    Odrv12 I__5947 (
            .O(N__32242),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__5946 (
            .O(N__32239),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    InMux I__5945 (
            .O(N__32232),
            .I(N__32227));
    InMux I__5944 (
            .O(N__32231),
            .I(N__32224));
    InMux I__5943 (
            .O(N__32230),
            .I(N__32220));
    LocalMux I__5942 (
            .O(N__32227),
            .I(N__32217));
    LocalMux I__5941 (
            .O(N__32224),
            .I(N__32214));
    InMux I__5940 (
            .O(N__32223),
            .I(N__32211));
    LocalMux I__5939 (
            .O(N__32220),
            .I(N__32208));
    Span4Mux_h I__5938 (
            .O(N__32217),
            .I(N__32205));
    Span4Mux_h I__5937 (
            .O(N__32214),
            .I(N__32200));
    LocalMux I__5936 (
            .O(N__32211),
            .I(N__32200));
    Span4Mux_h I__5935 (
            .O(N__32208),
            .I(N__32195));
    Span4Mux_v I__5934 (
            .O(N__32205),
            .I(N__32195));
    Span4Mux_h I__5933 (
            .O(N__32200),
            .I(N__32192));
    Odrv4 I__5932 (
            .O(N__32195),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    Odrv4 I__5931 (
            .O(N__32192),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__5930 (
            .O(N__32187),
            .I(N__32181));
    InMux I__5929 (
            .O(N__32186),
            .I(N__32181));
    LocalMux I__5928 (
            .O(N__32181),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ));
    CEMux I__5927 (
            .O(N__32178),
            .I(N__32173));
    CEMux I__5926 (
            .O(N__32177),
            .I(N__32166));
    CEMux I__5925 (
            .O(N__32176),
            .I(N__32163));
    LocalMux I__5924 (
            .O(N__32173),
            .I(N__32160));
    InMux I__5923 (
            .O(N__32172),
            .I(N__32157));
    CEMux I__5922 (
            .O(N__32171),
            .I(N__32154));
    CEMux I__5921 (
            .O(N__32170),
            .I(N__32151));
    CEMux I__5920 (
            .O(N__32169),
            .I(N__32136));
    LocalMux I__5919 (
            .O(N__32166),
            .I(N__32122));
    LocalMux I__5918 (
            .O(N__32163),
            .I(N__32122));
    Span4Mux_v I__5917 (
            .O(N__32160),
            .I(N__32122));
    LocalMux I__5916 (
            .O(N__32157),
            .I(N__32122));
    LocalMux I__5915 (
            .O(N__32154),
            .I(N__32122));
    LocalMux I__5914 (
            .O(N__32151),
            .I(N__32119));
    InMux I__5913 (
            .O(N__32150),
            .I(N__32097));
    InMux I__5912 (
            .O(N__32149),
            .I(N__32097));
    InMux I__5911 (
            .O(N__32148),
            .I(N__32097));
    InMux I__5910 (
            .O(N__32147),
            .I(N__32088));
    InMux I__5909 (
            .O(N__32146),
            .I(N__32088));
    InMux I__5908 (
            .O(N__32145),
            .I(N__32088));
    InMux I__5907 (
            .O(N__32144),
            .I(N__32088));
    InMux I__5906 (
            .O(N__32143),
            .I(N__32075));
    InMux I__5905 (
            .O(N__32142),
            .I(N__32075));
    InMux I__5904 (
            .O(N__32141),
            .I(N__32075));
    InMux I__5903 (
            .O(N__32140),
            .I(N__32075));
    CEMux I__5902 (
            .O(N__32139),
            .I(N__32071));
    LocalMux I__5901 (
            .O(N__32136),
            .I(N__32068));
    CEMux I__5900 (
            .O(N__32135),
            .I(N__32065));
    CEMux I__5899 (
            .O(N__32134),
            .I(N__32062));
    CEMux I__5898 (
            .O(N__32133),
            .I(N__32059));
    Span4Mux_v I__5897 (
            .O(N__32122),
            .I(N__32056));
    Span4Mux_v I__5896 (
            .O(N__32119),
            .I(N__32053));
    InMux I__5895 (
            .O(N__32118),
            .I(N__32044));
    InMux I__5894 (
            .O(N__32117),
            .I(N__32044));
    InMux I__5893 (
            .O(N__32116),
            .I(N__32044));
    InMux I__5892 (
            .O(N__32115),
            .I(N__32044));
    InMux I__5891 (
            .O(N__32114),
            .I(N__32035));
    InMux I__5890 (
            .O(N__32113),
            .I(N__32035));
    InMux I__5889 (
            .O(N__32112),
            .I(N__32035));
    InMux I__5888 (
            .O(N__32111),
            .I(N__32035));
    InMux I__5887 (
            .O(N__32110),
            .I(N__32028));
    InMux I__5886 (
            .O(N__32109),
            .I(N__32028));
    InMux I__5885 (
            .O(N__32108),
            .I(N__32028));
    InMux I__5884 (
            .O(N__32107),
            .I(N__32019));
    InMux I__5883 (
            .O(N__32106),
            .I(N__32019));
    InMux I__5882 (
            .O(N__32105),
            .I(N__32019));
    InMux I__5881 (
            .O(N__32104),
            .I(N__32019));
    LocalMux I__5880 (
            .O(N__32097),
            .I(N__32016));
    LocalMux I__5879 (
            .O(N__32088),
            .I(N__32013));
    InMux I__5878 (
            .O(N__32087),
            .I(N__32004));
    InMux I__5877 (
            .O(N__32086),
            .I(N__32004));
    InMux I__5876 (
            .O(N__32085),
            .I(N__32004));
    InMux I__5875 (
            .O(N__32084),
            .I(N__32004));
    LocalMux I__5874 (
            .O(N__32075),
            .I(N__32001));
    CEMux I__5873 (
            .O(N__32074),
            .I(N__31998));
    LocalMux I__5872 (
            .O(N__32071),
            .I(N__31995));
    Span4Mux_h I__5871 (
            .O(N__32068),
            .I(N__31992));
    LocalMux I__5870 (
            .O(N__32065),
            .I(N__31981));
    LocalMux I__5869 (
            .O(N__32062),
            .I(N__31981));
    LocalMux I__5868 (
            .O(N__32059),
            .I(N__31981));
    Span4Mux_v I__5867 (
            .O(N__32056),
            .I(N__31981));
    Span4Mux_h I__5866 (
            .O(N__32053),
            .I(N__31981));
    LocalMux I__5865 (
            .O(N__32044),
            .I(N__31970));
    LocalMux I__5864 (
            .O(N__32035),
            .I(N__31970));
    LocalMux I__5863 (
            .O(N__32028),
            .I(N__31970));
    LocalMux I__5862 (
            .O(N__32019),
            .I(N__31970));
    Span4Mux_v I__5861 (
            .O(N__32016),
            .I(N__31970));
    Span4Mux_h I__5860 (
            .O(N__32013),
            .I(N__31963));
    LocalMux I__5859 (
            .O(N__32004),
            .I(N__31963));
    Span4Mux_v I__5858 (
            .O(N__32001),
            .I(N__31963));
    LocalMux I__5857 (
            .O(N__31998),
            .I(N__31960));
    Span4Mux_v I__5856 (
            .O(N__31995),
            .I(N__31957));
    Span4Mux_h I__5855 (
            .O(N__31992),
            .I(N__31954));
    Span4Mux_v I__5854 (
            .O(N__31981),
            .I(N__31951));
    Span4Mux_v I__5853 (
            .O(N__31970),
            .I(N__31946));
    Span4Mux_v I__5852 (
            .O(N__31963),
            .I(N__31946));
    Odrv12 I__5851 (
            .O(N__31960),
            .I(\phase_controller_inst1.m3 ));
    Odrv4 I__5850 (
            .O(N__31957),
            .I(\phase_controller_inst1.m3 ));
    Odrv4 I__5849 (
            .O(N__31954),
            .I(\phase_controller_inst1.m3 ));
    Odrv4 I__5848 (
            .O(N__31951),
            .I(\phase_controller_inst1.m3 ));
    Odrv4 I__5847 (
            .O(N__31946),
            .I(\phase_controller_inst1.m3 ));
    InMux I__5846 (
            .O(N__31935),
            .I(N__31932));
    LocalMux I__5845 (
            .O(N__31932),
            .I(N__31929));
    Span4Mux_v I__5844 (
            .O(N__31929),
            .I(N__31926));
    Span4Mux_v I__5843 (
            .O(N__31926),
            .I(N__31923));
    Span4Mux_h I__5842 (
            .O(N__31923),
            .I(N__31920));
    Odrv4 I__5841 (
            .O(N__31920),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    CascadeMux I__5840 (
            .O(N__31917),
            .I(N__31914));
    InMux I__5839 (
            .O(N__31914),
            .I(N__31911));
    LocalMux I__5838 (
            .O(N__31911),
            .I(N__31906));
    InMux I__5837 (
            .O(N__31910),
            .I(N__31903));
    InMux I__5836 (
            .O(N__31909),
            .I(N__31900));
    Span4Mux_v I__5835 (
            .O(N__31906),
            .I(N__31897));
    LocalMux I__5834 (
            .O(N__31903),
            .I(N__31894));
    LocalMux I__5833 (
            .O(N__31900),
            .I(N__31891));
    Odrv4 I__5832 (
            .O(N__31897),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv12 I__5831 (
            .O(N__31894),
            .I(\current_shift_inst.un4_control_input1_10 ));
    Odrv4 I__5830 (
            .O(N__31891),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__5829 (
            .O(N__31884),
            .I(N__31881));
    LocalMux I__5828 (
            .O(N__31881),
            .I(N__31878));
    Span4Mux_h I__5827 (
            .O(N__31878),
            .I(N__31875));
    Span4Mux_v I__5826 (
            .O(N__31875),
            .I(N__31872));
    Odrv4 I__5825 (
            .O(N__31872),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    InMux I__5824 (
            .O(N__31869),
            .I(N__31866));
    LocalMux I__5823 (
            .O(N__31866),
            .I(N__31862));
    CascadeMux I__5822 (
            .O(N__31865),
            .I(N__31858));
    Span12Mux_h I__5821 (
            .O(N__31862),
            .I(N__31855));
    InMux I__5820 (
            .O(N__31861),
            .I(N__31852));
    InMux I__5819 (
            .O(N__31858),
            .I(N__31849));
    Odrv12 I__5818 (
            .O(N__31855),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__5817 (
            .O(N__31852),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__5816 (
            .O(N__31849),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    CascadeMux I__5815 (
            .O(N__31842),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__5814 (
            .O(N__31839),
            .I(N__31835));
    CascadeMux I__5813 (
            .O(N__31838),
            .I(N__31832));
    LocalMux I__5812 (
            .O(N__31835),
            .I(N__31829));
    InMux I__5811 (
            .O(N__31832),
            .I(N__31826));
    Span4Mux_h I__5810 (
            .O(N__31829),
            .I(N__31821));
    LocalMux I__5809 (
            .O(N__31826),
            .I(N__31821));
    Span4Mux_v I__5808 (
            .O(N__31821),
            .I(N__31818));
    Odrv4 I__5807 (
            .O(N__31818),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__5806 (
            .O(N__31815),
            .I(N__31812));
    LocalMux I__5805 (
            .O(N__31812),
            .I(N__31807));
    InMux I__5804 (
            .O(N__31811),
            .I(N__31802));
    InMux I__5803 (
            .O(N__31810),
            .I(N__31802));
    Span4Mux_h I__5802 (
            .O(N__31807),
            .I(N__31796));
    LocalMux I__5801 (
            .O(N__31802),
            .I(N__31796));
    InMux I__5800 (
            .O(N__31801),
            .I(N__31793));
    Span4Mux_h I__5799 (
            .O(N__31796),
            .I(N__31790));
    LocalMux I__5798 (
            .O(N__31793),
            .I(N__31787));
    Odrv4 I__5797 (
            .O(N__31790),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    Odrv12 I__5796 (
            .O(N__31787),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__5795 (
            .O(N__31782),
            .I(N__31779));
    LocalMux I__5794 (
            .O(N__31779),
            .I(N__31775));
    InMux I__5793 (
            .O(N__31778),
            .I(N__31772));
    Odrv4 I__5792 (
            .O(N__31775),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    LocalMux I__5791 (
            .O(N__31772),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    InMux I__5790 (
            .O(N__31767),
            .I(N__31763));
    InMux I__5789 (
            .O(N__31766),
            .I(N__31759));
    LocalMux I__5788 (
            .O(N__31763),
            .I(N__31756));
    InMux I__5787 (
            .O(N__31762),
            .I(N__31753));
    LocalMux I__5786 (
            .O(N__31759),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    Odrv4 I__5785 (
            .O(N__31756),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    LocalMux I__5784 (
            .O(N__31753),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__5783 (
            .O(N__31746),
            .I(N__31742));
    CascadeMux I__5782 (
            .O(N__31745),
            .I(N__31737));
    LocalMux I__5781 (
            .O(N__31742),
            .I(N__31734));
    InMux I__5780 (
            .O(N__31741),
            .I(N__31731));
    InMux I__5779 (
            .O(N__31740),
            .I(N__31728));
    InMux I__5778 (
            .O(N__31737),
            .I(N__31725));
    Span4Mux_h I__5777 (
            .O(N__31734),
            .I(N__31720));
    LocalMux I__5776 (
            .O(N__31731),
            .I(N__31720));
    LocalMux I__5775 (
            .O(N__31728),
            .I(N__31715));
    LocalMux I__5774 (
            .O(N__31725),
            .I(N__31715));
    Span4Mux_h I__5773 (
            .O(N__31720),
            .I(N__31712));
    Span4Mux_h I__5772 (
            .O(N__31715),
            .I(N__31709));
    Odrv4 I__5771 (
            .O(N__31712),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    Odrv4 I__5770 (
            .O(N__31709),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    CEMux I__5769 (
            .O(N__31704),
            .I(N__31668));
    CEMux I__5768 (
            .O(N__31703),
            .I(N__31668));
    CEMux I__5767 (
            .O(N__31702),
            .I(N__31668));
    CEMux I__5766 (
            .O(N__31701),
            .I(N__31668));
    CEMux I__5765 (
            .O(N__31700),
            .I(N__31668));
    CEMux I__5764 (
            .O(N__31699),
            .I(N__31668));
    CEMux I__5763 (
            .O(N__31698),
            .I(N__31668));
    CEMux I__5762 (
            .O(N__31697),
            .I(N__31668));
    CEMux I__5761 (
            .O(N__31696),
            .I(N__31668));
    CEMux I__5760 (
            .O(N__31695),
            .I(N__31668));
    CEMux I__5759 (
            .O(N__31694),
            .I(N__31668));
    CEMux I__5758 (
            .O(N__31693),
            .I(N__31668));
    GlobalMux I__5757 (
            .O(N__31668),
            .I(N__31665));
    gio2CtrlBuf I__5756 (
            .O(N__31665),
            .I(\phase_controller_inst2.stoper_tr.un1_start_g ));
    InMux I__5755 (
            .O(N__31662),
            .I(N__31656));
    InMux I__5754 (
            .O(N__31661),
            .I(N__31656));
    LocalMux I__5753 (
            .O(N__31656),
            .I(N__31653));
    Odrv12 I__5752 (
            .O(N__31653),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ));
    CascadeMux I__5751 (
            .O(N__31650),
            .I(N__31647));
    InMux I__5750 (
            .O(N__31647),
            .I(N__31641));
    InMux I__5749 (
            .O(N__31646),
            .I(N__31641));
    LocalMux I__5748 (
            .O(N__31641),
            .I(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ));
    InMux I__5747 (
            .O(N__31638),
            .I(N__31635));
    LocalMux I__5746 (
            .O(N__31635),
            .I(N__31632));
    Span4Mux_h I__5745 (
            .O(N__31632),
            .I(N__31629));
    Odrv4 I__5744 (
            .O(N__31629),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt16 ));
    InMux I__5743 (
            .O(N__31626),
            .I(N__31620));
    InMux I__5742 (
            .O(N__31625),
            .I(N__31620));
    LocalMux I__5741 (
            .O(N__31620),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ));
    CascadeMux I__5740 (
            .O(N__31617),
            .I(N__31612));
    InMux I__5739 (
            .O(N__31616),
            .I(N__31609));
    InMux I__5738 (
            .O(N__31615),
            .I(N__31604));
    InMux I__5737 (
            .O(N__31612),
            .I(N__31604));
    LocalMux I__5736 (
            .O(N__31609),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    LocalMux I__5735 (
            .O(N__31604),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ));
    CascadeMux I__5734 (
            .O(N__31599),
            .I(N__31595));
    InMux I__5733 (
            .O(N__31598),
            .I(N__31591));
    InMux I__5732 (
            .O(N__31595),
            .I(N__31588));
    InMux I__5731 (
            .O(N__31594),
            .I(N__31585));
    LocalMux I__5730 (
            .O(N__31591),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__5729 (
            .O(N__31588),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    LocalMux I__5728 (
            .O(N__31585),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__5727 (
            .O(N__31578),
            .I(N__31574));
    InMux I__5726 (
            .O(N__31577),
            .I(N__31571));
    LocalMux I__5725 (
            .O(N__31574),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    LocalMux I__5724 (
            .O(N__31571),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ));
    CascadeMux I__5723 (
            .O(N__31566),
            .I(N__31563));
    InMux I__5722 (
            .O(N__31563),
            .I(N__31560));
    LocalMux I__5721 (
            .O(N__31560),
            .I(N__31557));
    Span4Mux_h I__5720 (
            .O(N__31557),
            .I(N__31554));
    Odrv4 I__5719 (
            .O(N__31554),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ));
    CascadeMux I__5718 (
            .O(N__31551),
            .I(N__31548));
    InMux I__5717 (
            .O(N__31548),
            .I(N__31545));
    LocalMux I__5716 (
            .O(N__31545),
            .I(N__31542));
    Span4Mux_h I__5715 (
            .O(N__31542),
            .I(N__31539));
    Odrv4 I__5714 (
            .O(N__31539),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt18 ));
    InMux I__5713 (
            .O(N__31536),
            .I(N__31530));
    InMux I__5712 (
            .O(N__31535),
            .I(N__31530));
    LocalMux I__5711 (
            .O(N__31530),
            .I(N__31526));
    InMux I__5710 (
            .O(N__31529),
            .I(N__31523));
    Span4Mux_h I__5709 (
            .O(N__31526),
            .I(N__31520));
    LocalMux I__5708 (
            .O(N__31523),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__5707 (
            .O(N__31520),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ));
    CascadeMux I__5706 (
            .O(N__31515),
            .I(N__31512));
    InMux I__5705 (
            .O(N__31512),
            .I(N__31506));
    InMux I__5704 (
            .O(N__31511),
            .I(N__31506));
    LocalMux I__5703 (
            .O(N__31506),
            .I(N__31502));
    InMux I__5702 (
            .O(N__31505),
            .I(N__31499));
    Span4Mux_h I__5701 (
            .O(N__31502),
            .I(N__31496));
    LocalMux I__5700 (
            .O(N__31499),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__5699 (
            .O(N__31496),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__5698 (
            .O(N__31491),
            .I(N__31488));
    LocalMux I__5697 (
            .O(N__31488),
            .I(N__31485));
    Odrv4 I__5696 (
            .O(N__31485),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ));
    InMux I__5695 (
            .O(N__31482),
            .I(N__31479));
    LocalMux I__5694 (
            .O(N__31479),
            .I(N__31476));
    Span4Mux_v I__5693 (
            .O(N__31476),
            .I(N__31473));
    Span4Mux_h I__5692 (
            .O(N__31473),
            .I(N__31466));
    InMux I__5691 (
            .O(N__31472),
            .I(N__31463));
    InMux I__5690 (
            .O(N__31471),
            .I(N__31460));
    InMux I__5689 (
            .O(N__31470),
            .I(N__31455));
    InMux I__5688 (
            .O(N__31469),
            .I(N__31455));
    Span4Mux_v I__5687 (
            .O(N__31466),
            .I(N__31448));
    LocalMux I__5686 (
            .O(N__31463),
            .I(N__31448));
    LocalMux I__5685 (
            .O(N__31460),
            .I(N__31448));
    LocalMux I__5684 (
            .O(N__31455),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    Odrv4 I__5683 (
            .O(N__31448),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__5682 (
            .O(N__31443),
            .I(N__31440));
    LocalMux I__5681 (
            .O(N__31440),
            .I(N__31436));
    InMux I__5680 (
            .O(N__31439),
            .I(N__31433));
    Odrv4 I__5679 (
            .O(N__31436),
            .I(\phase_controller_inst2.un4_running_cry_30_THRU_CO ));
    LocalMux I__5678 (
            .O(N__31433),
            .I(\phase_controller_inst2.un4_running_cry_30_THRU_CO ));
    InMux I__5677 (
            .O(N__31428),
            .I(N__31422));
    InMux I__5676 (
            .O(N__31427),
            .I(N__31422));
    LocalMux I__5675 (
            .O(N__31422),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ));
    CascadeMux I__5674 (
            .O(N__31419),
            .I(N__31415));
    InMux I__5673 (
            .O(N__31418),
            .I(N__31410));
    InMux I__5672 (
            .O(N__31415),
            .I(N__31410));
    LocalMux I__5671 (
            .O(N__31410),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ));
    InMux I__5670 (
            .O(N__31407),
            .I(N__31404));
    LocalMux I__5669 (
            .O(N__31404),
            .I(N__31398));
    InMux I__5668 (
            .O(N__31403),
            .I(N__31393));
    InMux I__5667 (
            .O(N__31402),
            .I(N__31393));
    InMux I__5666 (
            .O(N__31401),
            .I(N__31390));
    Span4Mux_h I__5665 (
            .O(N__31398),
            .I(N__31387));
    LocalMux I__5664 (
            .O(N__31393),
            .I(N__31384));
    LocalMux I__5663 (
            .O(N__31390),
            .I(N__31381));
    Span4Mux_h I__5662 (
            .O(N__31387),
            .I(N__31378));
    Span4Mux_h I__5661 (
            .O(N__31384),
            .I(N__31375));
    Span4Mux_v I__5660 (
            .O(N__31381),
            .I(N__31372));
    Odrv4 I__5659 (
            .O(N__31378),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__5658 (
            .O(N__31375),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    Odrv4 I__5657 (
            .O(N__31372),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__5656 (
            .O(N__31365),
            .I(N__31362));
    LocalMux I__5655 (
            .O(N__31362),
            .I(N__31359));
    Span4Mux_h I__5654 (
            .O(N__31359),
            .I(N__31355));
    InMux I__5653 (
            .O(N__31358),
            .I(N__31352));
    Odrv4 I__5652 (
            .O(N__31355),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    LocalMux I__5651 (
            .O(N__31352),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__5650 (
            .O(N__31347),
            .I(N__31341));
    InMux I__5649 (
            .O(N__31346),
            .I(N__31341));
    LocalMux I__5648 (
            .O(N__31341),
            .I(N__31338));
    Span4Mux_h I__5647 (
            .O(N__31338),
            .I(N__31335));
    Odrv4 I__5646 (
            .O(N__31335),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ));
    CascadeMux I__5645 (
            .O(N__31332),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ));
    InMux I__5644 (
            .O(N__31329),
            .I(N__31326));
    LocalMux I__5643 (
            .O(N__31326),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ));
    InMux I__5642 (
            .O(N__31323),
            .I(N__31320));
    LocalMux I__5641 (
            .O(N__31320),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ));
    InMux I__5640 (
            .O(N__31317),
            .I(N__31314));
    LocalMux I__5639 (
            .O(N__31314),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ));
    InMux I__5638 (
            .O(N__31311),
            .I(N__31307));
    InMux I__5637 (
            .O(N__31310),
            .I(N__31304));
    LocalMux I__5636 (
            .O(N__31307),
            .I(N__31299));
    LocalMux I__5635 (
            .O(N__31304),
            .I(N__31299));
    Span4Mux_h I__5634 (
            .O(N__31299),
            .I(N__31296));
    Span4Mux_h I__5633 (
            .O(N__31296),
            .I(N__31293));
    Span4Mux_v I__5632 (
            .O(N__31293),
            .I(N__31290));
    Span4Mux_v I__5631 (
            .O(N__31290),
            .I(N__31285));
    InMux I__5630 (
            .O(N__31289),
            .I(N__31282));
    InMux I__5629 (
            .O(N__31288),
            .I(N__31279));
    Span4Mux_v I__5628 (
            .O(N__31285),
            .I(N__31276));
    LocalMux I__5627 (
            .O(N__31282),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    LocalMux I__5626 (
            .O(N__31279),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__5625 (
            .O(N__31276),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__5624 (
            .O(N__31269),
            .I(N__31263));
    ClkMux I__5623 (
            .O(N__31268),
            .I(N__31263));
    GlobalMux I__5622 (
            .O(N__31263),
            .I(N__31260));
    gio2CtrlBuf I__5621 (
            .O(N__31260),
            .I(delay_tr_input_c_g));
    IoInMux I__5620 (
            .O(N__31257),
            .I(N__31254));
    LocalMux I__5619 (
            .O(N__31254),
            .I(N__31251));
    IoSpan4Mux I__5618 (
            .O(N__31251),
            .I(N__31248));
    Span4Mux_s1_v I__5617 (
            .O(N__31248),
            .I(N__31245));
    Odrv4 I__5616 (
            .O(N__31245),
            .I(s3_phy_c));
    IoInMux I__5615 (
            .O(N__31242),
            .I(N__31239));
    LocalMux I__5614 (
            .O(N__31239),
            .I(N__31236));
    Span4Mux_s0_v I__5613 (
            .O(N__31236),
            .I(N__31233));
    Odrv4 I__5612 (
            .O(N__31233),
            .I(GB_BUFFER_red_c_g_THRU_CO));
    InMux I__5611 (
            .O(N__31230),
            .I(N__31227));
    LocalMux I__5610 (
            .O(N__31227),
            .I(\phase_controller_inst1.stoper_hc.m34_1 ));
    InMux I__5609 (
            .O(N__31224),
            .I(N__31214));
    InMux I__5608 (
            .O(N__31223),
            .I(N__31214));
    InMux I__5607 (
            .O(N__31222),
            .I(N__31214));
    InMux I__5606 (
            .O(N__31221),
            .I(N__31210));
    LocalMux I__5605 (
            .O(N__31214),
            .I(N__31207));
    CascadeMux I__5604 (
            .O(N__31213),
            .I(N__31204));
    LocalMux I__5603 (
            .O(N__31210),
            .I(N__31199));
    Span4Mux_v I__5602 (
            .O(N__31207),
            .I(N__31199));
    InMux I__5601 (
            .O(N__31204),
            .I(N__31196));
    Span4Mux_h I__5600 (
            .O(N__31199),
            .I(N__31193));
    LocalMux I__5599 (
            .O(N__31196),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__5598 (
            .O(N__31193),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    InMux I__5597 (
            .O(N__31188),
            .I(N__31185));
    LocalMux I__5596 (
            .O(N__31185),
            .I(\phase_controller_inst2.stoper_hc.m10Z0Z_1 ));
    InMux I__5595 (
            .O(N__31182),
            .I(N__31179));
    LocalMux I__5594 (
            .O(N__31179),
            .I(N__31176));
    Span4Mux_v I__5593 (
            .O(N__31176),
            .I(N__31173));
    Odrv4 I__5592 (
            .O(N__31173),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__5591 (
            .O(N__31170),
            .I(N__31167));
    LocalMux I__5590 (
            .O(N__31167),
            .I(N__31164));
    Span4Mux_h I__5589 (
            .O(N__31164),
            .I(N__31161));
    Odrv4 I__5588 (
            .O(N__31161),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__5587 (
            .O(N__31158),
            .I(N__31155));
    LocalMux I__5586 (
            .O(N__31155),
            .I(N__31152));
    Span4Mux_h I__5585 (
            .O(N__31152),
            .I(N__31149));
    Odrv4 I__5584 (
            .O(N__31149),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__5583 (
            .O(N__31146),
            .I(N__31143));
    LocalMux I__5582 (
            .O(N__31143),
            .I(N__31140));
    Span4Mux_h I__5581 (
            .O(N__31140),
            .I(N__31137));
    Odrv4 I__5580 (
            .O(N__31137),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__5579 (
            .O(N__31134),
            .I(N__31131));
    LocalMux I__5578 (
            .O(N__31131),
            .I(N__31128));
    Span4Mux_h I__5577 (
            .O(N__31128),
            .I(N__31125));
    Odrv4 I__5576 (
            .O(N__31125),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    InMux I__5575 (
            .O(N__31122),
            .I(N__31119));
    LocalMux I__5574 (
            .O(N__31119),
            .I(N__31116));
    Odrv12 I__5573 (
            .O(N__31116),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__5572 (
            .O(N__31113),
            .I(N__31110));
    LocalMux I__5571 (
            .O(N__31110),
            .I(N__31105));
    InMux I__5570 (
            .O(N__31109),
            .I(N__31102));
    InMux I__5569 (
            .O(N__31108),
            .I(N__31099));
    Span4Mux_v I__5568 (
            .O(N__31105),
            .I(N__31096));
    LocalMux I__5567 (
            .O(N__31102),
            .I(N__31093));
    LocalMux I__5566 (
            .O(N__31099),
            .I(N__31090));
    Odrv4 I__5565 (
            .O(N__31096),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__5564 (
            .O(N__31093),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv12 I__5563 (
            .O(N__31090),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__5562 (
            .O(N__31083),
            .I(N__31080));
    LocalMux I__5561 (
            .O(N__31080),
            .I(N__31077));
    Span4Mux_h I__5560 (
            .O(N__31077),
            .I(N__31074));
    Odrv4 I__5559 (
            .O(N__31074),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__5558 (
            .O(N__31071),
            .I(N__31068));
    LocalMux I__5557 (
            .O(N__31068),
            .I(N__31065));
    Odrv4 I__5556 (
            .O(N__31065),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__5555 (
            .O(N__31062),
            .I(N__31059));
    LocalMux I__5554 (
            .O(N__31059),
            .I(N__31056));
    Span4Mux_v I__5553 (
            .O(N__31056),
            .I(N__31053));
    Odrv4 I__5552 (
            .O(N__31053),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    CascadeMux I__5551 (
            .O(N__31050),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ));
    InMux I__5550 (
            .O(N__31047),
            .I(N__31044));
    LocalMux I__5549 (
            .O(N__31044),
            .I(N__31041));
    Span4Mux_h I__5548 (
            .O(N__31041),
            .I(N__31038));
    Odrv4 I__5547 (
            .O(N__31038),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__5546 (
            .O(N__31035),
            .I(N__31032));
    LocalMux I__5545 (
            .O(N__31032),
            .I(N__31029));
    Span4Mux_h I__5544 (
            .O(N__31029),
            .I(N__31026));
    Odrv4 I__5543 (
            .O(N__31026),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__5542 (
            .O(N__31023),
            .I(N__31020));
    LocalMux I__5541 (
            .O(N__31020),
            .I(N__31017));
    Span4Mux_h I__5540 (
            .O(N__31017),
            .I(N__31014));
    Odrv4 I__5539 (
            .O(N__31014),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__5538 (
            .O(N__31011),
            .I(N__31008));
    LocalMux I__5537 (
            .O(N__31008),
            .I(N__31005));
    Span4Mux_v I__5536 (
            .O(N__31005),
            .I(N__31002));
    Odrv4 I__5535 (
            .O(N__31002),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    CascadeMux I__5534 (
            .O(N__30999),
            .I(N__30996));
    InMux I__5533 (
            .O(N__30996),
            .I(N__30993));
    LocalMux I__5532 (
            .O(N__30993),
            .I(N__30990));
    Span4Mux_v I__5531 (
            .O(N__30990),
            .I(N__30987));
    Odrv4 I__5530 (
            .O(N__30987),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__5529 (
            .O(N__30984),
            .I(N__30981));
    LocalMux I__5528 (
            .O(N__30981),
            .I(N__30978));
    Span4Mux_v I__5527 (
            .O(N__30978),
            .I(N__30975));
    Span4Mux_h I__5526 (
            .O(N__30975),
            .I(N__30972));
    Odrv4 I__5525 (
            .O(N__30972),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__5524 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__5523 (
            .O(N__30966),
            .I(N__30963));
    Odrv12 I__5522 (
            .O(N__30963),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__5521 (
            .O(N__30960),
            .I(N__30957));
    LocalMux I__5520 (
            .O(N__30957),
            .I(N__30954));
    Span4Mux_h I__5519 (
            .O(N__30954),
            .I(N__30951));
    Odrv4 I__5518 (
            .O(N__30951),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__5517 (
            .O(N__30948),
            .I(N__30945));
    LocalMux I__5516 (
            .O(N__30945),
            .I(N__30942));
    Span4Mux_h I__5515 (
            .O(N__30942),
            .I(N__30939));
    Odrv4 I__5514 (
            .O(N__30939),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__5513 (
            .O(N__30936),
            .I(N__30933));
    LocalMux I__5512 (
            .O(N__30933),
            .I(N__30930));
    Span4Mux_h I__5511 (
            .O(N__30930),
            .I(N__30927));
    Odrv4 I__5510 (
            .O(N__30927),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__5509 (
            .O(N__30924),
            .I(N__30921));
    LocalMux I__5508 (
            .O(N__30921),
            .I(N__30918));
    Span4Mux_v I__5507 (
            .O(N__30918),
            .I(N__30915));
    Odrv4 I__5506 (
            .O(N__30915),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__5505 (
            .O(N__30912),
            .I(N__30909));
    LocalMux I__5504 (
            .O(N__30909),
            .I(N__30906));
    Odrv4 I__5503 (
            .O(N__30906),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    CascadeMux I__5502 (
            .O(N__30903),
            .I(N__30900));
    InMux I__5501 (
            .O(N__30900),
            .I(N__30897));
    LocalMux I__5500 (
            .O(N__30897),
            .I(N__30893));
    InMux I__5499 (
            .O(N__30896),
            .I(N__30890));
    Span4Mux_v I__5498 (
            .O(N__30893),
            .I(N__30884));
    LocalMux I__5497 (
            .O(N__30890),
            .I(N__30884));
    InMux I__5496 (
            .O(N__30889),
            .I(N__30881));
    Span4Mux_v I__5495 (
            .O(N__30884),
            .I(N__30878));
    LocalMux I__5494 (
            .O(N__30881),
            .I(N__30875));
    Odrv4 I__5493 (
            .O(N__30878),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv12 I__5492 (
            .O(N__30875),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__5491 (
            .O(N__30870),
            .I(N__30867));
    LocalMux I__5490 (
            .O(N__30867),
            .I(N__30864));
    Odrv4 I__5489 (
            .O(N__30864),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    InMux I__5488 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__5487 (
            .O(N__30858),
            .I(N__30855));
    Span4Mux_v I__5486 (
            .O(N__30855),
            .I(N__30852));
    Odrv4 I__5485 (
            .O(N__30852),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__5484 (
            .O(N__30849),
            .I(N__30846));
    LocalMux I__5483 (
            .O(N__30846),
            .I(N__30843));
    Odrv4 I__5482 (
            .O(N__30843),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__5481 (
            .O(N__30840),
            .I(N__30837));
    LocalMux I__5480 (
            .O(N__30837),
            .I(N__30834));
    Span4Mux_v I__5479 (
            .O(N__30834),
            .I(N__30831));
    Odrv4 I__5478 (
            .O(N__30831),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__5477 (
            .O(N__30828),
            .I(N__30825));
    LocalMux I__5476 (
            .O(N__30825),
            .I(N__30822));
    Span4Mux_h I__5475 (
            .O(N__30822),
            .I(N__30819));
    Odrv4 I__5474 (
            .O(N__30819),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__5473 (
            .O(N__30816),
            .I(N__30813));
    LocalMux I__5472 (
            .O(N__30813),
            .I(N__30810));
    Span4Mux_h I__5471 (
            .O(N__30810),
            .I(N__30807));
    Odrv4 I__5470 (
            .O(N__30807),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__5469 (
            .O(N__30804),
            .I(N__30801));
    LocalMux I__5468 (
            .O(N__30801),
            .I(N__30798));
    Span4Mux_v I__5467 (
            .O(N__30798),
            .I(N__30795));
    Odrv4 I__5466 (
            .O(N__30795),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    CascadeMux I__5465 (
            .O(N__30792),
            .I(N__30789));
    InMux I__5464 (
            .O(N__30789),
            .I(N__30785));
    InMux I__5463 (
            .O(N__30788),
            .I(N__30782));
    LocalMux I__5462 (
            .O(N__30785),
            .I(N__30779));
    LocalMux I__5461 (
            .O(N__30782),
            .I(N__30776));
    Span4Mux_v I__5460 (
            .O(N__30779),
            .I(N__30773));
    Span4Mux_v I__5459 (
            .O(N__30776),
            .I(N__30770));
    Span4Mux_v I__5458 (
            .O(N__30773),
            .I(N__30766));
    Span4Mux_h I__5457 (
            .O(N__30770),
            .I(N__30763));
    InMux I__5456 (
            .O(N__30769),
            .I(N__30760));
    Odrv4 I__5455 (
            .O(N__30766),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__5454 (
            .O(N__30763),
            .I(\current_shift_inst.un4_control_input1_30 ));
    LocalMux I__5453 (
            .O(N__30760),
            .I(\current_shift_inst.un4_control_input1_30 ));
    CascadeMux I__5452 (
            .O(N__30753),
            .I(N__30750));
    InMux I__5451 (
            .O(N__30750),
            .I(N__30747));
    LocalMux I__5450 (
            .O(N__30747),
            .I(N__30744));
    Odrv4 I__5449 (
            .O(N__30744),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__5448 (
            .O(N__30741),
            .I(N__30738));
    LocalMux I__5447 (
            .O(N__30738),
            .I(N__30735));
    Odrv12 I__5446 (
            .O(N__30735),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__5445 (
            .O(N__30732),
            .I(N__30729));
    LocalMux I__5444 (
            .O(N__30729),
            .I(N__30726));
    Span4Mux_h I__5443 (
            .O(N__30726),
            .I(N__30723));
    Odrv4 I__5442 (
            .O(N__30723),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__5441 (
            .O(N__30720),
            .I(N__30717));
    LocalMux I__5440 (
            .O(N__30717),
            .I(N__30714));
    Odrv4 I__5439 (
            .O(N__30714),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__5438 (
            .O(N__30711),
            .I(N__30708));
    LocalMux I__5437 (
            .O(N__30708),
            .I(N__30705));
    Span4Mux_h I__5436 (
            .O(N__30705),
            .I(N__30702));
    Odrv4 I__5435 (
            .O(N__30702),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    CascadeMux I__5434 (
            .O(N__30699),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    InMux I__5433 (
            .O(N__30696),
            .I(N__30692));
    InMux I__5432 (
            .O(N__30695),
            .I(N__30689));
    LocalMux I__5431 (
            .O(N__30692),
            .I(N__30686));
    LocalMux I__5430 (
            .O(N__30689),
            .I(N__30683));
    Span4Mux_v I__5429 (
            .O(N__30686),
            .I(N__30680));
    Span4Mux_v I__5428 (
            .O(N__30683),
            .I(N__30677));
    Span4Mux_h I__5427 (
            .O(N__30680),
            .I(N__30674));
    Sp12to4 I__5426 (
            .O(N__30677),
            .I(N__30671));
    Span4Mux_h I__5425 (
            .O(N__30674),
            .I(N__30668));
    Span12Mux_h I__5424 (
            .O(N__30671),
            .I(N__30665));
    Odrv4 I__5423 (
            .O(N__30668),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv12 I__5422 (
            .O(N__30665),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    InMux I__5421 (
            .O(N__30660),
            .I(N__30657));
    LocalMux I__5420 (
            .O(N__30657),
            .I(N__30654));
    Span4Mux_h I__5419 (
            .O(N__30654),
            .I(N__30651));
    Odrv4 I__5418 (
            .O(N__30651),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__5417 (
            .O(N__30648),
            .I(N__30645));
    LocalMux I__5416 (
            .O(N__30645),
            .I(N__30642));
    Span4Mux_h I__5415 (
            .O(N__30642),
            .I(N__30639));
    Odrv4 I__5414 (
            .O(N__30639),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__5413 (
            .O(N__30636),
            .I(N__30633));
    LocalMux I__5412 (
            .O(N__30633),
            .I(N__30630));
    Odrv12 I__5411 (
            .O(N__30630),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__5410 (
            .O(N__30627),
            .I(N__30624));
    LocalMux I__5409 (
            .O(N__30624),
            .I(N__30621));
    Span4Mux_h I__5408 (
            .O(N__30621),
            .I(N__30618));
    Odrv4 I__5407 (
            .O(N__30618),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__5406 (
            .O(N__30615),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__5405 (
            .O(N__30612),
            .I(N__30609));
    LocalMux I__5404 (
            .O(N__30609),
            .I(N__30606));
    Span4Mux_v I__5403 (
            .O(N__30606),
            .I(N__30602));
    InMux I__5402 (
            .O(N__30605),
            .I(N__30599));
    Span4Mux_h I__5401 (
            .O(N__30602),
            .I(N__30593));
    LocalMux I__5400 (
            .O(N__30599),
            .I(N__30593));
    InMux I__5399 (
            .O(N__30598),
            .I(N__30590));
    Sp12to4 I__5398 (
            .O(N__30593),
            .I(N__30585));
    LocalMux I__5397 (
            .O(N__30590),
            .I(N__30585));
    Odrv12 I__5396 (
            .O(N__30585),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__5395 (
            .O(N__30582),
            .I(N__30578));
    InMux I__5394 (
            .O(N__30581),
            .I(N__30575));
    LocalMux I__5393 (
            .O(N__30578),
            .I(N__30572));
    LocalMux I__5392 (
            .O(N__30575),
            .I(N__30569));
    Span4Mux_v I__5391 (
            .O(N__30572),
            .I(N__30565));
    Span4Mux_h I__5390 (
            .O(N__30569),
            .I(N__30562));
    InMux I__5389 (
            .O(N__30568),
            .I(N__30559));
    Odrv4 I__5388 (
            .O(N__30565),
            .I(\current_shift_inst.un4_control_input1_26 ));
    Odrv4 I__5387 (
            .O(N__30562),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__5386 (
            .O(N__30559),
            .I(\current_shift_inst.un4_control_input1_26 ));
    CascadeMux I__5385 (
            .O(N__30552),
            .I(N__30549));
    InMux I__5384 (
            .O(N__30549),
            .I(N__30546));
    LocalMux I__5383 (
            .O(N__30546),
            .I(N__30543));
    Odrv4 I__5382 (
            .O(N__30543),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__5381 (
            .O(N__30540),
            .I(N__30537));
    InMux I__5380 (
            .O(N__30537),
            .I(N__30533));
    CascadeMux I__5379 (
            .O(N__30536),
            .I(N__30530));
    LocalMux I__5378 (
            .O(N__30533),
            .I(N__30527));
    InMux I__5377 (
            .O(N__30530),
            .I(N__30524));
    Span4Mux_v I__5376 (
            .O(N__30527),
            .I(N__30520));
    LocalMux I__5375 (
            .O(N__30524),
            .I(N__30517));
    InMux I__5374 (
            .O(N__30523),
            .I(N__30514));
    Odrv4 I__5373 (
            .O(N__30520),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv12 I__5372 (
            .O(N__30517),
            .I(\current_shift_inst.un4_control_input1_19 ));
    LocalMux I__5371 (
            .O(N__30514),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__5370 (
            .O(N__30507),
            .I(N__30504));
    LocalMux I__5369 (
            .O(N__30504),
            .I(N__30501));
    Odrv4 I__5368 (
            .O(N__30501),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    InMux I__5367 (
            .O(N__30498),
            .I(N__30495));
    LocalMux I__5366 (
            .O(N__30495),
            .I(N__30492));
    Span4Mux_h I__5365 (
            .O(N__30492),
            .I(N__30489));
    Odrv4 I__5364 (
            .O(N__30489),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__5363 (
            .O(N__30486),
            .I(N__30483));
    LocalMux I__5362 (
            .O(N__30483),
            .I(N__30480));
    Odrv12 I__5361 (
            .O(N__30480),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__5360 (
            .O(N__30477),
            .I(N__30474));
    LocalMux I__5359 (
            .O(N__30474),
            .I(N__30471));
    Odrv12 I__5358 (
            .O(N__30471),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__5357 (
            .O(N__30468),
            .I(N__30465));
    LocalMux I__5356 (
            .O(N__30465),
            .I(N__30462));
    Span12Mux_v I__5355 (
            .O(N__30462),
            .I(N__30459));
    Odrv12 I__5354 (
            .O(N__30459),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__5353 (
            .O(N__30456),
            .I(N__30453));
    LocalMux I__5352 (
            .O(N__30453),
            .I(N__30450));
    Span4Mux_h I__5351 (
            .O(N__30450),
            .I(N__30447));
    Odrv4 I__5350 (
            .O(N__30447),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__5349 (
            .O(N__30444),
            .I(N__30441));
    LocalMux I__5348 (
            .O(N__30441),
            .I(N__30438));
    Odrv12 I__5347 (
            .O(N__30438),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__5346 (
            .O(N__30435),
            .I(N__30432));
    LocalMux I__5345 (
            .O(N__30432),
            .I(N__30429));
    Span4Mux_h I__5344 (
            .O(N__30429),
            .I(N__30426));
    Odrv4 I__5343 (
            .O(N__30426),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__5342 (
            .O(N__30423),
            .I(N__30420));
    LocalMux I__5341 (
            .O(N__30420),
            .I(N__30417));
    Odrv12 I__5340 (
            .O(N__30417),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__5339 (
            .O(N__30414),
            .I(N__30411));
    LocalMux I__5338 (
            .O(N__30411),
            .I(N__30408));
    Span4Mux_h I__5337 (
            .O(N__30408),
            .I(N__30403));
    InMux I__5336 (
            .O(N__30407),
            .I(N__30400));
    InMux I__5335 (
            .O(N__30406),
            .I(N__30397));
    Span4Mux_v I__5334 (
            .O(N__30403),
            .I(N__30394));
    LocalMux I__5333 (
            .O(N__30400),
            .I(N__30391));
    LocalMux I__5332 (
            .O(N__30397),
            .I(N__30388));
    Odrv4 I__5331 (
            .O(N__30394),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv12 I__5330 (
            .O(N__30391),
            .I(\current_shift_inst.un4_control_input1_13 ));
    Odrv4 I__5329 (
            .O(N__30388),
            .I(\current_shift_inst.un4_control_input1_13 ));
    CascadeMux I__5328 (
            .O(N__30381),
            .I(N__30378));
    InMux I__5327 (
            .O(N__30378),
            .I(N__30375));
    LocalMux I__5326 (
            .O(N__30375),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__5325 (
            .O(N__30372),
            .I(N__30368));
    InMux I__5324 (
            .O(N__30371),
            .I(N__30365));
    LocalMux I__5323 (
            .O(N__30368),
            .I(N__30361));
    LocalMux I__5322 (
            .O(N__30365),
            .I(N__30358));
    InMux I__5321 (
            .O(N__30364),
            .I(N__30355));
    Span4Mux_h I__5320 (
            .O(N__30361),
            .I(N__30352));
    Span4Mux_h I__5319 (
            .O(N__30358),
            .I(N__30347));
    LocalMux I__5318 (
            .O(N__30355),
            .I(N__30347));
    Odrv4 I__5317 (
            .O(N__30352),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__5316 (
            .O(N__30347),
            .I(\current_shift_inst.un4_control_input1_24 ));
    CascadeMux I__5315 (
            .O(N__30342),
            .I(N__30339));
    InMux I__5314 (
            .O(N__30339),
            .I(N__30336));
    LocalMux I__5313 (
            .O(N__30336),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    InMux I__5312 (
            .O(N__30333),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__5311 (
            .O(N__30330),
            .I(N__30326));
    InMux I__5310 (
            .O(N__30329),
            .I(N__30323));
    LocalMux I__5309 (
            .O(N__30326),
            .I(N__30317));
    LocalMux I__5308 (
            .O(N__30323),
            .I(N__30317));
    InMux I__5307 (
            .O(N__30322),
            .I(N__30314));
    Span4Mux_v I__5306 (
            .O(N__30317),
            .I(N__30309));
    LocalMux I__5305 (
            .O(N__30314),
            .I(N__30309));
    Span4Mux_h I__5304 (
            .O(N__30309),
            .I(N__30306));
    Odrv4 I__5303 (
            .O(N__30306),
            .I(\current_shift_inst.un4_control_input1_23 ));
    InMux I__5302 (
            .O(N__30303),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__5301 (
            .O(N__30300),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__5300 (
            .O(N__30297),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__5299 (
            .O(N__30294),
            .I(bfn_12_16_0_));
    InMux I__5298 (
            .O(N__30291),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    CascadeMux I__5297 (
            .O(N__30288),
            .I(N__30284));
    InMux I__5296 (
            .O(N__30287),
            .I(N__30280));
    InMux I__5295 (
            .O(N__30284),
            .I(N__30275));
    InMux I__5294 (
            .O(N__30283),
            .I(N__30275));
    LocalMux I__5293 (
            .O(N__30280),
            .I(N__30272));
    LocalMux I__5292 (
            .O(N__30275),
            .I(N__30267));
    Span4Mux_v I__5291 (
            .O(N__30272),
            .I(N__30267));
    Span4Mux_h I__5290 (
            .O(N__30267),
            .I(N__30264));
    Odrv4 I__5289 (
            .O(N__30264),
            .I(\current_shift_inst.un4_control_input1_28 ));
    InMux I__5288 (
            .O(N__30261),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__5287 (
            .O(N__30258),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__5286 (
            .O(N__30255),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__5285 (
            .O(N__30252),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__5284 (
            .O(N__30249),
            .I(N__30244));
    InMux I__5283 (
            .O(N__30248),
            .I(N__30241));
    InMux I__5282 (
            .O(N__30247),
            .I(N__30238));
    LocalMux I__5281 (
            .O(N__30244),
            .I(N__30233));
    LocalMux I__5280 (
            .O(N__30241),
            .I(N__30233));
    LocalMux I__5279 (
            .O(N__30238),
            .I(N__30230));
    Span4Mux_h I__5278 (
            .O(N__30233),
            .I(N__30227));
    Odrv4 I__5277 (
            .O(N__30230),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__5276 (
            .O(N__30227),
            .I(\current_shift_inst.un4_control_input1_14 ));
    InMux I__5275 (
            .O(N__30222),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__5274 (
            .O(N__30219),
            .I(N__30214));
    InMux I__5273 (
            .O(N__30218),
            .I(N__30211));
    InMux I__5272 (
            .O(N__30217),
            .I(N__30208));
    LocalMux I__5271 (
            .O(N__30214),
            .I(N__30205));
    LocalMux I__5270 (
            .O(N__30211),
            .I(N__30200));
    LocalMux I__5269 (
            .O(N__30208),
            .I(N__30200));
    Span12Mux_h I__5268 (
            .O(N__30205),
            .I(N__30197));
    Span4Mux_h I__5267 (
            .O(N__30200),
            .I(N__30194));
    Odrv12 I__5266 (
            .O(N__30197),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__5265 (
            .O(N__30194),
            .I(\current_shift_inst.un4_control_input1_15 ));
    InMux I__5264 (
            .O(N__30189),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__5263 (
            .O(N__30186),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__5262 (
            .O(N__30183),
            .I(N__30178));
    InMux I__5261 (
            .O(N__30182),
            .I(N__30175));
    InMux I__5260 (
            .O(N__30181),
            .I(N__30172));
    LocalMux I__5259 (
            .O(N__30178),
            .I(N__30167));
    LocalMux I__5258 (
            .O(N__30175),
            .I(N__30167));
    LocalMux I__5257 (
            .O(N__30172),
            .I(N__30164));
    Span4Mux_h I__5256 (
            .O(N__30167),
            .I(N__30159));
    Span4Mux_v I__5255 (
            .O(N__30164),
            .I(N__30159));
    Odrv4 I__5254 (
            .O(N__30159),
            .I(\current_shift_inst.un4_control_input1_17 ));
    InMux I__5253 (
            .O(N__30156),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__5252 (
            .O(N__30153),
            .I(bfn_12_15_0_));
    InMux I__5251 (
            .O(N__30150),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__5250 (
            .O(N__30147),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__5249 (
            .O(N__30144),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__5248 (
            .O(N__30141),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    CascadeMux I__5247 (
            .O(N__30138),
            .I(N__30135));
    InMux I__5246 (
            .O(N__30135),
            .I(N__30130));
    InMux I__5245 (
            .O(N__30134),
            .I(N__30127));
    InMux I__5244 (
            .O(N__30133),
            .I(N__30124));
    LocalMux I__5243 (
            .O(N__30130),
            .I(N__30121));
    LocalMux I__5242 (
            .O(N__30127),
            .I(N__30116));
    LocalMux I__5241 (
            .O(N__30124),
            .I(N__30116));
    Span4Mux_v I__5240 (
            .O(N__30121),
            .I(N__30113));
    Span4Mux_h I__5239 (
            .O(N__30116),
            .I(N__30110));
    Odrv4 I__5238 (
            .O(N__30113),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv4 I__5237 (
            .O(N__30110),
            .I(\current_shift_inst.un4_control_input1_6 ));
    InMux I__5236 (
            .O(N__30105),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__5235 (
            .O(N__30102),
            .I(N__30097));
    InMux I__5234 (
            .O(N__30101),
            .I(N__30094));
    InMux I__5233 (
            .O(N__30100),
            .I(N__30091));
    LocalMux I__5232 (
            .O(N__30097),
            .I(N__30088));
    LocalMux I__5231 (
            .O(N__30094),
            .I(N__30083));
    LocalMux I__5230 (
            .O(N__30091),
            .I(N__30083));
    Span4Mux_h I__5229 (
            .O(N__30088),
            .I(N__30080));
    Span4Mux_v I__5228 (
            .O(N__30083),
            .I(N__30077));
    Odrv4 I__5227 (
            .O(N__30080),
            .I(\current_shift_inst.un4_control_input1_7 ));
    Odrv4 I__5226 (
            .O(N__30077),
            .I(\current_shift_inst.un4_control_input1_7 ));
    InMux I__5225 (
            .O(N__30072),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__5224 (
            .O(N__30069),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__5223 (
            .O(N__30066),
            .I(N__30061));
    InMux I__5222 (
            .O(N__30065),
            .I(N__30058));
    InMux I__5221 (
            .O(N__30064),
            .I(N__30055));
    LocalMux I__5220 (
            .O(N__30061),
            .I(N__30052));
    LocalMux I__5219 (
            .O(N__30058),
            .I(N__30049));
    LocalMux I__5218 (
            .O(N__30055),
            .I(N__30044));
    Span4Mux_v I__5217 (
            .O(N__30052),
            .I(N__30044));
    Span4Mux_h I__5216 (
            .O(N__30049),
            .I(N__30041));
    Span4Mux_v I__5215 (
            .O(N__30044),
            .I(N__30038));
    Odrv4 I__5214 (
            .O(N__30041),
            .I(\current_shift_inst.un4_control_input1_9 ));
    Odrv4 I__5213 (
            .O(N__30038),
            .I(\current_shift_inst.un4_control_input1_9 ));
    InMux I__5212 (
            .O(N__30033),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__5211 (
            .O(N__30030),
            .I(bfn_12_14_0_));
    InMux I__5210 (
            .O(N__30027),
            .I(N__30024));
    LocalMux I__5209 (
            .O(N__30024),
            .I(N__30020));
    CascadeMux I__5208 (
            .O(N__30023),
            .I(N__30017));
    Span4Mux_v I__5207 (
            .O(N__30020),
            .I(N__30013));
    InMux I__5206 (
            .O(N__30017),
            .I(N__30008));
    InMux I__5205 (
            .O(N__30016),
            .I(N__30008));
    Span4Mux_h I__5204 (
            .O(N__30013),
            .I(N__30005));
    LocalMux I__5203 (
            .O(N__30008),
            .I(N__30002));
    Odrv4 I__5202 (
            .O(N__30005),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__5201 (
            .O(N__30002),
            .I(\current_shift_inst.un4_control_input1_11 ));
    InMux I__5200 (
            .O(N__29997),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__5199 (
            .O(N__29994),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__5198 (
            .O(N__29991),
            .I(N__29971));
    InMux I__5197 (
            .O(N__29990),
            .I(N__29971));
    InMux I__5196 (
            .O(N__29989),
            .I(N__29971));
    InMux I__5195 (
            .O(N__29988),
            .I(N__29971));
    InMux I__5194 (
            .O(N__29987),
            .I(N__29962));
    InMux I__5193 (
            .O(N__29986),
            .I(N__29962));
    InMux I__5192 (
            .O(N__29985),
            .I(N__29962));
    InMux I__5191 (
            .O(N__29984),
            .I(N__29962));
    InMux I__5190 (
            .O(N__29983),
            .I(N__29934));
    InMux I__5189 (
            .O(N__29982),
            .I(N__29934));
    InMux I__5188 (
            .O(N__29981),
            .I(N__29934));
    InMux I__5187 (
            .O(N__29980),
            .I(N__29934));
    LocalMux I__5186 (
            .O(N__29971),
            .I(N__29929));
    LocalMux I__5185 (
            .O(N__29962),
            .I(N__29929));
    InMux I__5184 (
            .O(N__29961),
            .I(N__29922));
    InMux I__5183 (
            .O(N__29960),
            .I(N__29922));
    InMux I__5182 (
            .O(N__29959),
            .I(N__29922));
    InMux I__5181 (
            .O(N__29958),
            .I(N__29913));
    InMux I__5180 (
            .O(N__29957),
            .I(N__29913));
    InMux I__5179 (
            .O(N__29956),
            .I(N__29913));
    InMux I__5178 (
            .O(N__29955),
            .I(N__29913));
    InMux I__5177 (
            .O(N__29954),
            .I(N__29909));
    InMux I__5176 (
            .O(N__29953),
            .I(N__29900));
    InMux I__5175 (
            .O(N__29952),
            .I(N__29900));
    InMux I__5174 (
            .O(N__29951),
            .I(N__29900));
    InMux I__5173 (
            .O(N__29950),
            .I(N__29900));
    InMux I__5172 (
            .O(N__29949),
            .I(N__29893));
    InMux I__5171 (
            .O(N__29948),
            .I(N__29893));
    InMux I__5170 (
            .O(N__29947),
            .I(N__29893));
    InMux I__5169 (
            .O(N__29946),
            .I(N__29884));
    InMux I__5168 (
            .O(N__29945),
            .I(N__29884));
    InMux I__5167 (
            .O(N__29944),
            .I(N__29884));
    InMux I__5166 (
            .O(N__29943),
            .I(N__29884));
    LocalMux I__5165 (
            .O(N__29934),
            .I(N__29881));
    Sp12to4 I__5164 (
            .O(N__29929),
            .I(N__29874));
    LocalMux I__5163 (
            .O(N__29922),
            .I(N__29874));
    LocalMux I__5162 (
            .O(N__29913),
            .I(N__29874));
    IoInMux I__5161 (
            .O(N__29912),
            .I(N__29871));
    LocalMux I__5160 (
            .O(N__29909),
            .I(N__29858));
    LocalMux I__5159 (
            .O(N__29900),
            .I(N__29858));
    LocalMux I__5158 (
            .O(N__29893),
            .I(N__29858));
    LocalMux I__5157 (
            .O(N__29884),
            .I(N__29858));
    Span12Mux_h I__5156 (
            .O(N__29881),
            .I(N__29858));
    Span12Mux_v I__5155 (
            .O(N__29874),
            .I(N__29858));
    LocalMux I__5154 (
            .O(N__29871),
            .I(N__29855));
    Odrv12 I__5153 (
            .O(N__29858),
            .I(\phase_controller_inst2.m3_0 ));
    Odrv4 I__5152 (
            .O(N__29855),
            .I(\phase_controller_inst2.m3_0 ));
    InMux I__5151 (
            .O(N__29850),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ));
    CascadeMux I__5150 (
            .O(N__29847),
            .I(N__29843));
    InMux I__5149 (
            .O(N__29846),
            .I(N__29838));
    InMux I__5148 (
            .O(N__29843),
            .I(N__29838));
    LocalMux I__5147 (
            .O(N__29838),
            .I(N__29834));
    InMux I__5146 (
            .O(N__29837),
            .I(N__29831));
    Span4Mux_h I__5145 (
            .O(N__29834),
            .I(N__29828));
    LocalMux I__5144 (
            .O(N__29831),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__5143 (
            .O(N__29828),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__5142 (
            .O(N__29823),
            .I(N__29820));
    LocalMux I__5141 (
            .O(N__29820),
            .I(N__29817));
    Span4Mux_v I__5140 (
            .O(N__29817),
            .I(N__29813));
    InMux I__5139 (
            .O(N__29816),
            .I(N__29810));
    Span4Mux_h I__5138 (
            .O(N__29813),
            .I(N__29803));
    LocalMux I__5137 (
            .O(N__29810),
            .I(N__29803));
    InMux I__5136 (
            .O(N__29809),
            .I(N__29800));
    InMux I__5135 (
            .O(N__29808),
            .I(N__29797));
    Odrv4 I__5134 (
            .O(N__29803),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__5133 (
            .O(N__29800),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__5132 (
            .O(N__29797),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__5131 (
            .O(N__29790),
            .I(N__29787));
    InMux I__5130 (
            .O(N__29787),
            .I(N__29784));
    LocalMux I__5129 (
            .O(N__29784),
            .I(N__29781));
    Span4Mux_v I__5128 (
            .O(N__29781),
            .I(N__29778));
    Span4Mux_h I__5127 (
            .O(N__29778),
            .I(N__29775));
    Odrv4 I__5126 (
            .O(N__29775),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__5125 (
            .O(N__29772),
            .I(N__29769));
    LocalMux I__5124 (
            .O(N__29769),
            .I(N__29765));
    CascadeMux I__5123 (
            .O(N__29768),
            .I(N__29762));
    Span4Mux_v I__5122 (
            .O(N__29765),
            .I(N__29757));
    InMux I__5121 (
            .O(N__29762),
            .I(N__29750));
    InMux I__5120 (
            .O(N__29761),
            .I(N__29750));
    InMux I__5119 (
            .O(N__29760),
            .I(N__29750));
    Odrv4 I__5118 (
            .O(N__29757),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__5117 (
            .O(N__29750),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__5116 (
            .O(N__29745),
            .I(N__29742));
    InMux I__5115 (
            .O(N__29742),
            .I(N__29739));
    LocalMux I__5114 (
            .O(N__29739),
            .I(N__29736));
    Span4Mux_v I__5113 (
            .O(N__29736),
            .I(N__29733));
    Odrv4 I__5112 (
            .O(N__29733),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__5111 (
            .O(N__29730),
            .I(N__29727));
    LocalMux I__5110 (
            .O(N__29727),
            .I(N__29724));
    Span12Mux_v I__5109 (
            .O(N__29724),
            .I(N__29721));
    Odrv12 I__5108 (
            .O(N__29721),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__5107 (
            .O(N__29718),
            .I(N__29715));
    LocalMux I__5106 (
            .O(N__29715),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    CascadeMux I__5105 (
            .O(N__29712),
            .I(N__29709));
    InMux I__5104 (
            .O(N__29709),
            .I(N__29706));
    LocalMux I__5103 (
            .O(N__29706),
            .I(N__29703));
    Span4Mux_v I__5102 (
            .O(N__29703),
            .I(N__29698));
    InMux I__5101 (
            .O(N__29702),
            .I(N__29693));
    InMux I__5100 (
            .O(N__29701),
            .I(N__29693));
    Odrv4 I__5099 (
            .O(N__29698),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__5098 (
            .O(N__29693),
            .I(\current_shift_inst.un4_control_input1_2 ));
    CascadeMux I__5097 (
            .O(N__29688),
            .I(N__29685));
    InMux I__5096 (
            .O(N__29685),
            .I(N__29681));
    InMux I__5095 (
            .O(N__29684),
            .I(N__29677));
    LocalMux I__5094 (
            .O(N__29681),
            .I(N__29674));
    InMux I__5093 (
            .O(N__29680),
            .I(N__29671));
    LocalMux I__5092 (
            .O(N__29677),
            .I(N__29668));
    Span4Mux_v I__5091 (
            .O(N__29674),
            .I(N__29665));
    LocalMux I__5090 (
            .O(N__29671),
            .I(N__29662));
    Span4Mux_v I__5089 (
            .O(N__29668),
            .I(N__29657));
    Span4Mux_h I__5088 (
            .O(N__29665),
            .I(N__29657));
    Span4Mux_h I__5087 (
            .O(N__29662),
            .I(N__29654));
    Odrv4 I__5086 (
            .O(N__29657),
            .I(\current_shift_inst.un4_control_input1_3 ));
    Odrv4 I__5085 (
            .O(N__29654),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__5084 (
            .O(N__29649),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__5083 (
            .O(N__29646),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    CascadeMux I__5082 (
            .O(N__29643),
            .I(N__29639));
    InMux I__5081 (
            .O(N__29642),
            .I(N__29634));
    InMux I__5080 (
            .O(N__29639),
            .I(N__29634));
    LocalMux I__5079 (
            .O(N__29634),
            .I(N__29631));
    Span4Mux_h I__5078 (
            .O(N__29631),
            .I(N__29627));
    InMux I__5077 (
            .O(N__29630),
            .I(N__29624));
    Span4Mux_v I__5076 (
            .O(N__29627),
            .I(N__29621));
    LocalMux I__5075 (
            .O(N__29624),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__5074 (
            .O(N__29621),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__5073 (
            .O(N__29616),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ));
    CascadeMux I__5072 (
            .O(N__29613),
            .I(N__29609));
    InMux I__5071 (
            .O(N__29612),
            .I(N__29605));
    InMux I__5070 (
            .O(N__29609),
            .I(N__29602));
    InMux I__5069 (
            .O(N__29608),
            .I(N__29599));
    LocalMux I__5068 (
            .O(N__29605),
            .I(N__29594));
    LocalMux I__5067 (
            .O(N__29602),
            .I(N__29594));
    LocalMux I__5066 (
            .O(N__29599),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv12 I__5065 (
            .O(N__29594),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__5064 (
            .O(N__29589),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ));
    CascadeMux I__5063 (
            .O(N__29586),
            .I(N__29582));
    InMux I__5062 (
            .O(N__29585),
            .I(N__29578));
    InMux I__5061 (
            .O(N__29582),
            .I(N__29575));
    InMux I__5060 (
            .O(N__29581),
            .I(N__29572));
    LocalMux I__5059 (
            .O(N__29578),
            .I(N__29567));
    LocalMux I__5058 (
            .O(N__29575),
            .I(N__29567));
    LocalMux I__5057 (
            .O(N__29572),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv12 I__5056 (
            .O(N__29567),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__5055 (
            .O(N__29562),
            .I(bfn_12_11_0_));
    InMux I__5054 (
            .O(N__29559),
            .I(N__29552));
    InMux I__5053 (
            .O(N__29558),
            .I(N__29552));
    InMux I__5052 (
            .O(N__29557),
            .I(N__29549));
    LocalMux I__5051 (
            .O(N__29552),
            .I(N__29546));
    LocalMux I__5050 (
            .O(N__29549),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv12 I__5049 (
            .O(N__29546),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__5048 (
            .O(N__29541),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ));
    CascadeMux I__5047 (
            .O(N__29538),
            .I(N__29534));
    InMux I__5046 (
            .O(N__29537),
            .I(N__29529));
    InMux I__5045 (
            .O(N__29534),
            .I(N__29529));
    LocalMux I__5044 (
            .O(N__29529),
            .I(N__29525));
    InMux I__5043 (
            .O(N__29528),
            .I(N__29522));
    Span4Mux_h I__5042 (
            .O(N__29525),
            .I(N__29519));
    LocalMux I__5041 (
            .O(N__29522),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__5040 (
            .O(N__29519),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__5039 (
            .O(N__29514),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__5038 (
            .O(N__29511),
            .I(N__29504));
    InMux I__5037 (
            .O(N__29510),
            .I(N__29504));
    InMux I__5036 (
            .O(N__29509),
            .I(N__29501));
    LocalMux I__5035 (
            .O(N__29504),
            .I(N__29498));
    LocalMux I__5034 (
            .O(N__29501),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__5033 (
            .O(N__29498),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__5032 (
            .O(N__29493),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ));
    CascadeMux I__5031 (
            .O(N__29490),
            .I(N__29486));
    InMux I__5030 (
            .O(N__29489),
            .I(N__29480));
    InMux I__5029 (
            .O(N__29486),
            .I(N__29480));
    InMux I__5028 (
            .O(N__29485),
            .I(N__29477));
    LocalMux I__5027 (
            .O(N__29480),
            .I(N__29474));
    LocalMux I__5026 (
            .O(N__29477),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__5025 (
            .O(N__29474),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__5024 (
            .O(N__29469),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__5023 (
            .O(N__29466),
            .I(N__29459));
    InMux I__5022 (
            .O(N__29465),
            .I(N__29459));
    InMux I__5021 (
            .O(N__29464),
            .I(N__29456));
    LocalMux I__5020 (
            .O(N__29459),
            .I(N__29453));
    LocalMux I__5019 (
            .O(N__29456),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__5018 (
            .O(N__29453),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__5017 (
            .O(N__29448),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__5016 (
            .O(N__29445),
            .I(N__29441));
    InMux I__5015 (
            .O(N__29444),
            .I(N__29438));
    LocalMux I__5014 (
            .O(N__29441),
            .I(N__29435));
    LocalMux I__5013 (
            .O(N__29438),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__5012 (
            .O(N__29435),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__5011 (
            .O(N__29430),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__5010 (
            .O(N__29427),
            .I(N__29424));
    LocalMux I__5009 (
            .O(N__29424),
            .I(N__29420));
    InMux I__5008 (
            .O(N__29423),
            .I(N__29417));
    Span4Mux_h I__5007 (
            .O(N__29420),
            .I(N__29414));
    LocalMux I__5006 (
            .O(N__29417),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv4 I__5005 (
            .O(N__29414),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__5004 (
            .O(N__29409),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ));
    InMux I__5003 (
            .O(N__29406),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__5002 (
            .O(N__29403),
            .I(bfn_12_10_0_));
    CascadeMux I__5001 (
            .O(N__29400),
            .I(N__29396));
    InMux I__5000 (
            .O(N__29399),
            .I(N__29391));
    InMux I__4999 (
            .O(N__29396),
            .I(N__29391));
    LocalMux I__4998 (
            .O(N__29391),
            .I(N__29387));
    InMux I__4997 (
            .O(N__29390),
            .I(N__29384));
    Span4Mux_v I__4996 (
            .O(N__29387),
            .I(N__29381));
    LocalMux I__4995 (
            .O(N__29384),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    Odrv4 I__4994 (
            .O(N__29381),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ));
    InMux I__4993 (
            .O(N__29376),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__4992 (
            .O(N__29373),
            .I(N__29366));
    InMux I__4991 (
            .O(N__29372),
            .I(N__29366));
    InMux I__4990 (
            .O(N__29371),
            .I(N__29363));
    LocalMux I__4989 (
            .O(N__29366),
            .I(N__29360));
    LocalMux I__4988 (
            .O(N__29363),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    Odrv4 I__4987 (
            .O(N__29360),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ));
    InMux I__4986 (
            .O(N__29355),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ));
    InMux I__4985 (
            .O(N__29352),
            .I(N__29346));
    InMux I__4984 (
            .O(N__29351),
            .I(N__29346));
    LocalMux I__4983 (
            .O(N__29346),
            .I(N__29342));
    InMux I__4982 (
            .O(N__29345),
            .I(N__29339));
    Span4Mux_h I__4981 (
            .O(N__29342),
            .I(N__29336));
    LocalMux I__4980 (
            .O(N__29339),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__4979 (
            .O(N__29336),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__4978 (
            .O(N__29331),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ));
    CascadeMux I__4977 (
            .O(N__29328),
            .I(N__29324));
    InMux I__4976 (
            .O(N__29327),
            .I(N__29319));
    InMux I__4975 (
            .O(N__29324),
            .I(N__29319));
    LocalMux I__4974 (
            .O(N__29319),
            .I(N__29315));
    InMux I__4973 (
            .O(N__29318),
            .I(N__29312));
    Span4Mux_v I__4972 (
            .O(N__29315),
            .I(N__29309));
    LocalMux I__4971 (
            .O(N__29312),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__4970 (
            .O(N__29309),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__4969 (
            .O(N__29304),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ));
    InMux I__4968 (
            .O(N__29301),
            .I(N__29295));
    InMux I__4967 (
            .O(N__29300),
            .I(N__29295));
    LocalMux I__4966 (
            .O(N__29295),
            .I(N__29291));
    InMux I__4965 (
            .O(N__29294),
            .I(N__29288));
    Span4Mux_h I__4964 (
            .O(N__29291),
            .I(N__29285));
    LocalMux I__4963 (
            .O(N__29288),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__4962 (
            .O(N__29285),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__4961 (
            .O(N__29280),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__4960 (
            .O(N__29277),
            .I(N__29274));
    LocalMux I__4959 (
            .O(N__29274),
            .I(N__29270));
    InMux I__4958 (
            .O(N__29273),
            .I(N__29267));
    Span4Mux_v I__4957 (
            .O(N__29270),
            .I(N__29264));
    LocalMux I__4956 (
            .O(N__29267),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__4955 (
            .O(N__29264),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__4954 (
            .O(N__29259),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__4953 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__4952 (
            .O(N__29253),
            .I(N__29249));
    InMux I__4951 (
            .O(N__29252),
            .I(N__29246));
    Span4Mux_h I__4950 (
            .O(N__29249),
            .I(N__29243));
    LocalMux I__4949 (
            .O(N__29246),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv4 I__4948 (
            .O(N__29243),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__4947 (
            .O(N__29238),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__4946 (
            .O(N__29235),
            .I(N__29232));
    LocalMux I__4945 (
            .O(N__29232),
            .I(N__29228));
    InMux I__4944 (
            .O(N__29231),
            .I(N__29225));
    Span4Mux_h I__4943 (
            .O(N__29228),
            .I(N__29222));
    LocalMux I__4942 (
            .O(N__29225),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv4 I__4941 (
            .O(N__29222),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__4940 (
            .O(N__29217),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__4939 (
            .O(N__29214),
            .I(N__29210));
    InMux I__4938 (
            .O(N__29213),
            .I(N__29207));
    LocalMux I__4937 (
            .O(N__29210),
            .I(N__29204));
    LocalMux I__4936 (
            .O(N__29207),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__4935 (
            .O(N__29204),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__4934 (
            .O(N__29199),
            .I(bfn_12_9_0_));
    InMux I__4933 (
            .O(N__29196),
            .I(N__29192));
    InMux I__4932 (
            .O(N__29195),
            .I(N__29189));
    LocalMux I__4931 (
            .O(N__29192),
            .I(N__29186));
    LocalMux I__4930 (
            .O(N__29189),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__4929 (
            .O(N__29186),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__4928 (
            .O(N__29181),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__4927 (
            .O(N__29178),
            .I(N__29174));
    InMux I__4926 (
            .O(N__29177),
            .I(N__29171));
    LocalMux I__4925 (
            .O(N__29174),
            .I(N__29168));
    LocalMux I__4924 (
            .O(N__29171),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv4 I__4923 (
            .O(N__29168),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__4922 (
            .O(N__29163),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__4921 (
            .O(N__29160),
            .I(N__29156));
    InMux I__4920 (
            .O(N__29159),
            .I(N__29153));
    LocalMux I__4919 (
            .O(N__29156),
            .I(N__29150));
    LocalMux I__4918 (
            .O(N__29153),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__4917 (
            .O(N__29150),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__4916 (
            .O(N__29145),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__4915 (
            .O(N__29142),
            .I(N__29139));
    LocalMux I__4914 (
            .O(N__29139),
            .I(N__29135));
    InMux I__4913 (
            .O(N__29138),
            .I(N__29132));
    Span4Mux_v I__4912 (
            .O(N__29135),
            .I(N__29129));
    LocalMux I__4911 (
            .O(N__29132),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__4910 (
            .O(N__29129),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__4909 (
            .O(N__29124),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__4908 (
            .O(N__29121),
            .I(N__29117));
    InMux I__4907 (
            .O(N__29120),
            .I(N__29114));
    LocalMux I__4906 (
            .O(N__29117),
            .I(N__29109));
    LocalMux I__4905 (
            .O(N__29114),
            .I(N__29109));
    Span4Mux_v I__4904 (
            .O(N__29109),
            .I(N__29106));
    Odrv4 I__4903 (
            .O(N__29106),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ));
    InMux I__4902 (
            .O(N__29103),
            .I(N__29099));
    InMux I__4901 (
            .O(N__29102),
            .I(N__29096));
    LocalMux I__4900 (
            .O(N__29099),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    LocalMux I__4899 (
            .O(N__29096),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ));
    InMux I__4898 (
            .O(N__29091),
            .I(N__29088));
    LocalMux I__4897 (
            .O(N__29088),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt24 ));
    InMux I__4896 (
            .O(N__29085),
            .I(N__29081));
    InMux I__4895 (
            .O(N__29084),
            .I(N__29078));
    LocalMux I__4894 (
            .O(N__29081),
            .I(N__29075));
    LocalMux I__4893 (
            .O(N__29078),
            .I(N__29069));
    Span4Mux_v I__4892 (
            .O(N__29075),
            .I(N__29066));
    InMux I__4891 (
            .O(N__29074),
            .I(N__29059));
    InMux I__4890 (
            .O(N__29073),
            .I(N__29059));
    InMux I__4889 (
            .O(N__29072),
            .I(N__29059));
    Odrv12 I__4888 (
            .O(N__29069),
            .I(\phase_controller_inst1.start_latched ));
    Odrv4 I__4887 (
            .O(N__29066),
            .I(\phase_controller_inst1.start_latched ));
    LocalMux I__4886 (
            .O(N__29059),
            .I(\phase_controller_inst1.start_latched ));
    CascadeMux I__4885 (
            .O(N__29052),
            .I(N__29049));
    InMux I__4884 (
            .O(N__29049),
            .I(N__29043));
    InMux I__4883 (
            .O(N__29048),
            .I(N__29043));
    LocalMux I__4882 (
            .O(N__29043),
            .I(N__29040));
    Odrv4 I__4881 (
            .O(N__29040),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ));
    InMux I__4880 (
            .O(N__29037),
            .I(N__29031));
    InMux I__4879 (
            .O(N__29036),
            .I(N__29031));
    LocalMux I__4878 (
            .O(N__29031),
            .I(N__29028));
    Span4Mux_v I__4877 (
            .O(N__29028),
            .I(N__29025));
    Span4Mux_h I__4876 (
            .O(N__29025),
            .I(N__29022));
    Odrv4 I__4875 (
            .O(N__29022),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ));
    InMux I__4874 (
            .O(N__29019),
            .I(N__29016));
    LocalMux I__4873 (
            .O(N__29016),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt26 ));
    InMux I__4872 (
            .O(N__29013),
            .I(N__29009));
    InMux I__4871 (
            .O(N__29012),
            .I(N__29005));
    LocalMux I__4870 (
            .O(N__29009),
            .I(N__29002));
    InMux I__4869 (
            .O(N__29008),
            .I(N__28999));
    LocalMux I__4868 (
            .O(N__29005),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__4867 (
            .O(N__29002),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__4866 (
            .O(N__28999),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__4865 (
            .O(N__28992),
            .I(N__28989));
    LocalMux I__4864 (
            .O(N__28989),
            .I(N__28985));
    InMux I__4863 (
            .O(N__28988),
            .I(N__28982));
    Odrv4 I__4862 (
            .O(N__28985),
            .I(\phase_controller_inst2.N_38 ));
    LocalMux I__4861 (
            .O(N__28982),
            .I(\phase_controller_inst2.N_38 ));
    InMux I__4860 (
            .O(N__28977),
            .I(N__28974));
    LocalMux I__4859 (
            .O(N__28974),
            .I(N__28970));
    InMux I__4858 (
            .O(N__28973),
            .I(N__28967));
    Span4Mux_h I__4857 (
            .O(N__28970),
            .I(N__28964));
    LocalMux I__4856 (
            .O(N__28967),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv4 I__4855 (
            .O(N__28964),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__4854 (
            .O(N__28959),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__4853 (
            .O(N__28956),
            .I(N__28952));
    CascadeMux I__4852 (
            .O(N__28955),
            .I(N__28949));
    InMux I__4851 (
            .O(N__28952),
            .I(N__28944));
    InMux I__4850 (
            .O(N__28949),
            .I(N__28944));
    LocalMux I__4849 (
            .O(N__28944),
            .I(\phase_controller_inst2.stoper_tr.N_38_i ));
    InMux I__4848 (
            .O(N__28941),
            .I(N__28937));
    InMux I__4847 (
            .O(N__28940),
            .I(N__28934));
    LocalMux I__4846 (
            .O(N__28937),
            .I(N__28931));
    LocalMux I__4845 (
            .O(N__28934),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__4844 (
            .O(N__28931),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__4843 (
            .O(N__28926),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__4842 (
            .O(N__28923),
            .I(N__28919));
    InMux I__4841 (
            .O(N__28922),
            .I(N__28916));
    LocalMux I__4840 (
            .O(N__28919),
            .I(N__28913));
    LocalMux I__4839 (
            .O(N__28916),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__4838 (
            .O(N__28913),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__4837 (
            .O(N__28908),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__4836 (
            .O(N__28905),
            .I(N__28901));
    InMux I__4835 (
            .O(N__28904),
            .I(N__28898));
    LocalMux I__4834 (
            .O(N__28901),
            .I(N__28895));
    LocalMux I__4833 (
            .O(N__28898),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__4832 (
            .O(N__28895),
            .I(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__4831 (
            .O(N__28890),
            .I(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ));
    CascadeMux I__4830 (
            .O(N__28887),
            .I(N__28884));
    InMux I__4829 (
            .O(N__28884),
            .I(N__28881));
    LocalMux I__4828 (
            .O(N__28881),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ));
    InMux I__4827 (
            .O(N__28878),
            .I(N__28874));
    InMux I__4826 (
            .O(N__28877),
            .I(N__28870));
    LocalMux I__4825 (
            .O(N__28874),
            .I(N__28867));
    InMux I__4824 (
            .O(N__28873),
            .I(N__28864));
    LocalMux I__4823 (
            .O(N__28870),
            .I(N__28861));
    Span12Mux_v I__4822 (
            .O(N__28867),
            .I(N__28858));
    LocalMux I__4821 (
            .O(N__28864),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv12 I__4820 (
            .O(N__28861),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    Odrv12 I__4819 (
            .O(N__28858),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__4818 (
            .O(N__28851),
            .I(N__28848));
    LocalMux I__4817 (
            .O(N__28848),
            .I(N__28843));
    InMux I__4816 (
            .O(N__28847),
            .I(N__28840));
    InMux I__4815 (
            .O(N__28846),
            .I(N__28836));
    Span4Mux_v I__4814 (
            .O(N__28843),
            .I(N__28833));
    LocalMux I__4813 (
            .O(N__28840),
            .I(N__28830));
    InMux I__4812 (
            .O(N__28839),
            .I(N__28827));
    LocalMux I__4811 (
            .O(N__28836),
            .I(N__28824));
    Span4Mux_h I__4810 (
            .O(N__28833),
            .I(N__28817));
    Span4Mux_v I__4809 (
            .O(N__28830),
            .I(N__28817));
    LocalMux I__4808 (
            .O(N__28827),
            .I(N__28817));
    Span4Mux_h I__4807 (
            .O(N__28824),
            .I(N__28814));
    Span4Mux_v I__4806 (
            .O(N__28817),
            .I(N__28811));
    Odrv4 I__4805 (
            .O(N__28814),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    Odrv4 I__4804 (
            .O(N__28811),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__4803 (
            .O(N__28806),
            .I(N__28803));
    LocalMux I__4802 (
            .O(N__28803),
            .I(N__28798));
    InMux I__4801 (
            .O(N__28802),
            .I(N__28795));
    InMux I__4800 (
            .O(N__28801),
            .I(N__28792));
    Span4Mux_h I__4799 (
            .O(N__28798),
            .I(N__28789));
    LocalMux I__4798 (
            .O(N__28795),
            .I(N__28786));
    LocalMux I__4797 (
            .O(N__28792),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv4 I__4796 (
            .O(N__28789),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    Odrv12 I__4795 (
            .O(N__28786),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    InMux I__4794 (
            .O(N__28779),
            .I(N__28775));
    InMux I__4793 (
            .O(N__28778),
            .I(N__28771));
    LocalMux I__4792 (
            .O(N__28775),
            .I(N__28768));
    InMux I__4791 (
            .O(N__28774),
            .I(N__28765));
    LocalMux I__4790 (
            .O(N__28771),
            .I(N__28761));
    Span4Mux_h I__4789 (
            .O(N__28768),
            .I(N__28756));
    LocalMux I__4788 (
            .O(N__28765),
            .I(N__28756));
    InMux I__4787 (
            .O(N__28764),
            .I(N__28753));
    Span4Mux_h I__4786 (
            .O(N__28761),
            .I(N__28750));
    Span4Mux_h I__4785 (
            .O(N__28756),
            .I(N__28745));
    LocalMux I__4784 (
            .O(N__28753),
            .I(N__28745));
    Odrv4 I__4783 (
            .O(N__28750),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__4782 (
            .O(N__28745),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    CascadeMux I__4781 (
            .O(N__28740),
            .I(N__28737));
    InMux I__4780 (
            .O(N__28737),
            .I(N__28734));
    LocalMux I__4779 (
            .O(N__28734),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ));
    InMux I__4778 (
            .O(N__28731),
            .I(N__28728));
    LocalMux I__4777 (
            .O(N__28728),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ));
    CascadeMux I__4776 (
            .O(N__28725),
            .I(N__28722));
    InMux I__4775 (
            .O(N__28722),
            .I(N__28719));
    LocalMux I__4774 (
            .O(N__28719),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt18 ));
    CascadeMux I__4773 (
            .O(N__28716),
            .I(N__28713));
    InMux I__4772 (
            .O(N__28713),
            .I(N__28710));
    LocalMux I__4771 (
            .O(N__28710),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ));
    InMux I__4770 (
            .O(N__28707),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    CascadeMux I__4769 (
            .O(N__28704),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_ ));
    InMux I__4768 (
            .O(N__28701),
            .I(N__28698));
    LocalMux I__4767 (
            .O(N__28698),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    InMux I__4766 (
            .O(N__28695),
            .I(N__28691));
    CascadeMux I__4765 (
            .O(N__28694),
            .I(N__28688));
    LocalMux I__4764 (
            .O(N__28691),
            .I(N__28685));
    InMux I__4763 (
            .O(N__28688),
            .I(N__28682));
    Span4Mux_v I__4762 (
            .O(N__28685),
            .I(N__28678));
    LocalMux I__4761 (
            .O(N__28682),
            .I(N__28675));
    InMux I__4760 (
            .O(N__28681),
            .I(N__28669));
    Span4Mux_h I__4759 (
            .O(N__28678),
            .I(N__28664));
    Span4Mux_v I__4758 (
            .O(N__28675),
            .I(N__28664));
    InMux I__4757 (
            .O(N__28674),
            .I(N__28659));
    InMux I__4756 (
            .O(N__28673),
            .I(N__28659));
    InMux I__4755 (
            .O(N__28672),
            .I(N__28656));
    LocalMux I__4754 (
            .O(N__28669),
            .I(N__28653));
    Odrv4 I__4753 (
            .O(N__28664),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__4752 (
            .O(N__28659),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    LocalMux I__4751 (
            .O(N__28656),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv12 I__4750 (
            .O(N__28653),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    CascadeMux I__4749 (
            .O(N__28644),
            .I(N__28641));
    InMux I__4748 (
            .O(N__28641),
            .I(N__28638));
    LocalMux I__4747 (
            .O(N__28638),
            .I(N__28635));
    Span4Mux_h I__4746 (
            .O(N__28635),
            .I(N__28632));
    Odrv4 I__4745 (
            .O(N__28632),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    CascadeMux I__4744 (
            .O(N__28629),
            .I(N__28625));
    InMux I__4743 (
            .O(N__28628),
            .I(N__28621));
    InMux I__4742 (
            .O(N__28625),
            .I(N__28616));
    InMux I__4741 (
            .O(N__28624),
            .I(N__28616));
    LocalMux I__4740 (
            .O(N__28621),
            .I(N__28611));
    LocalMux I__4739 (
            .O(N__28616),
            .I(N__28611));
    Span4Mux_h I__4738 (
            .O(N__28611),
            .I(N__28608));
    Span4Mux_h I__4737 (
            .O(N__28608),
            .I(N__28605));
    Span4Mux_v I__4736 (
            .O(N__28605),
            .I(N__28602));
    Span4Mux_v I__4735 (
            .O(N__28602),
            .I(N__28599));
    Span4Mux_v I__4734 (
            .O(N__28599),
            .I(N__28596));
    Odrv4 I__4733 (
            .O(N__28596),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    IoInMux I__4732 (
            .O(N__28593),
            .I(N__28590));
    LocalMux I__4731 (
            .O(N__28590),
            .I(N__28587));
    Span4Mux_s1_v I__4730 (
            .O(N__28587),
            .I(N__28584));
    Span4Mux_h I__4729 (
            .O(N__28584),
            .I(N__28581));
    Odrv4 I__4728 (
            .O(N__28581),
            .I(s4_phy_c));
    InMux I__4727 (
            .O(N__28578),
            .I(N__28575));
    LocalMux I__4726 (
            .O(N__28575),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__4725 (
            .O(N__28572),
            .I(N__28569));
    LocalMux I__4724 (
            .O(N__28569),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    CascadeMux I__4723 (
            .O(N__28566),
            .I(N__28563));
    InMux I__4722 (
            .O(N__28563),
            .I(N__28560));
    LocalMux I__4721 (
            .O(N__28560),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__4720 (
            .O(N__28557),
            .I(N__28554));
    LocalMux I__4719 (
            .O(N__28554),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__4718 (
            .O(N__28551),
            .I(N__28548));
    InMux I__4717 (
            .O(N__28548),
            .I(N__28545));
    LocalMux I__4716 (
            .O(N__28545),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    InMux I__4715 (
            .O(N__28542),
            .I(N__28539));
    LocalMux I__4714 (
            .O(N__28539),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__4713 (
            .O(N__28536),
            .I(N__28533));
    InMux I__4712 (
            .O(N__28533),
            .I(N__28530));
    LocalMux I__4711 (
            .O(N__28530),
            .I(N__28527));
    Odrv4 I__4710 (
            .O(N__28527),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__4709 (
            .O(N__28524),
            .I(N__28521));
    LocalMux I__4708 (
            .O(N__28521),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__4707 (
            .O(N__28518),
            .I(N__28515));
    InMux I__4706 (
            .O(N__28515),
            .I(N__28512));
    LocalMux I__4705 (
            .O(N__28512),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    CascadeMux I__4704 (
            .O(N__28509),
            .I(N__28506));
    InMux I__4703 (
            .O(N__28506),
            .I(N__28503));
    LocalMux I__4702 (
            .O(N__28503),
            .I(N__28500));
    Odrv4 I__4701 (
            .O(N__28500),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__4700 (
            .O(N__28497),
            .I(N__28494));
    InMux I__4699 (
            .O(N__28494),
            .I(N__28488));
    InMux I__4698 (
            .O(N__28493),
            .I(N__28488));
    LocalMux I__4697 (
            .O(N__28488),
            .I(N__28484));
    InMux I__4696 (
            .O(N__28487),
            .I(N__28481));
    Span4Mux_h I__4695 (
            .O(N__28484),
            .I(N__28478));
    LocalMux I__4694 (
            .O(N__28481),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    Odrv4 I__4693 (
            .O(N__28478),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ));
    InMux I__4692 (
            .O(N__28473),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ));
    InMux I__4691 (
            .O(N__28470),
            .I(N__28464));
    InMux I__4690 (
            .O(N__28469),
            .I(N__28464));
    LocalMux I__4689 (
            .O(N__28464),
            .I(N__28460));
    InMux I__4688 (
            .O(N__28463),
            .I(N__28457));
    Span4Mux_h I__4687 (
            .O(N__28460),
            .I(N__28454));
    LocalMux I__4686 (
            .O(N__28457),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    Odrv4 I__4685 (
            .O(N__28454),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ));
    InMux I__4684 (
            .O(N__28449),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ));
    InMux I__4683 (
            .O(N__28446),
            .I(N__28440));
    InMux I__4682 (
            .O(N__28445),
            .I(N__28440));
    LocalMux I__4681 (
            .O(N__28440),
            .I(N__28436));
    InMux I__4680 (
            .O(N__28439),
            .I(N__28433));
    Span4Mux_h I__4679 (
            .O(N__28436),
            .I(N__28430));
    LocalMux I__4678 (
            .O(N__28433),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    Odrv4 I__4677 (
            .O(N__28430),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ));
    InMux I__4676 (
            .O(N__28425),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ));
    InMux I__4675 (
            .O(N__28422),
            .I(N__28419));
    LocalMux I__4674 (
            .O(N__28419),
            .I(N__28414));
    InMux I__4673 (
            .O(N__28418),
            .I(N__28411));
    InMux I__4672 (
            .O(N__28417),
            .I(N__28408));
    Span4Mux_h I__4671 (
            .O(N__28414),
            .I(N__28403));
    LocalMux I__4670 (
            .O(N__28411),
            .I(N__28403));
    LocalMux I__4669 (
            .O(N__28408),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    Odrv4 I__4668 (
            .O(N__28403),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ));
    InMux I__4667 (
            .O(N__28398),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ));
    InMux I__4666 (
            .O(N__28395),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ));
    InMux I__4665 (
            .O(N__28392),
            .I(N__28388));
    InMux I__4664 (
            .O(N__28391),
            .I(N__28385));
    LocalMux I__4663 (
            .O(N__28388),
            .I(N__28381));
    LocalMux I__4662 (
            .O(N__28385),
            .I(N__28378));
    InMux I__4661 (
            .O(N__28384),
            .I(N__28375));
    Span4Mux_h I__4660 (
            .O(N__28381),
            .I(N__28372));
    Span4Mux_v I__4659 (
            .O(N__28378),
            .I(N__28369));
    LocalMux I__4658 (
            .O(N__28375),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__4657 (
            .O(N__28372),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    Odrv4 I__4656 (
            .O(N__28369),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ));
    InMux I__4655 (
            .O(N__28362),
            .I(N__28359));
    LocalMux I__4654 (
            .O(N__28359),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__4653 (
            .O(N__28356),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ));
    InMux I__4652 (
            .O(N__28353),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ));
    CascadeMux I__4651 (
            .O(N__28350),
            .I(N__28346));
    InMux I__4650 (
            .O(N__28349),
            .I(N__28341));
    InMux I__4649 (
            .O(N__28346),
            .I(N__28341));
    LocalMux I__4648 (
            .O(N__28341),
            .I(N__28337));
    InMux I__4647 (
            .O(N__28340),
            .I(N__28334));
    Span4Mux_v I__4646 (
            .O(N__28337),
            .I(N__28331));
    LocalMux I__4645 (
            .O(N__28334),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    Odrv4 I__4644 (
            .O(N__28331),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ));
    InMux I__4643 (
            .O(N__28326),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ));
    InMux I__4642 (
            .O(N__28323),
            .I(N__28317));
    InMux I__4641 (
            .O(N__28322),
            .I(N__28317));
    LocalMux I__4640 (
            .O(N__28317),
            .I(N__28313));
    InMux I__4639 (
            .O(N__28316),
            .I(N__28310));
    Span4Mux_h I__4638 (
            .O(N__28313),
            .I(N__28307));
    LocalMux I__4637 (
            .O(N__28310),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    Odrv4 I__4636 (
            .O(N__28307),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ));
    InMux I__4635 (
            .O(N__28302),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ));
    CascadeMux I__4634 (
            .O(N__28299),
            .I(N__28296));
    InMux I__4633 (
            .O(N__28296),
            .I(N__28290));
    InMux I__4632 (
            .O(N__28295),
            .I(N__28290));
    LocalMux I__4631 (
            .O(N__28290),
            .I(N__28286));
    InMux I__4630 (
            .O(N__28289),
            .I(N__28283));
    Span4Mux_v I__4629 (
            .O(N__28286),
            .I(N__28280));
    LocalMux I__4628 (
            .O(N__28283),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    Odrv4 I__4627 (
            .O(N__28280),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ));
    InMux I__4626 (
            .O(N__28275),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ));
    InMux I__4625 (
            .O(N__28272),
            .I(N__28266));
    InMux I__4624 (
            .O(N__28271),
            .I(N__28266));
    LocalMux I__4623 (
            .O(N__28266),
            .I(N__28262));
    InMux I__4622 (
            .O(N__28265),
            .I(N__28259));
    Span4Mux_v I__4621 (
            .O(N__28262),
            .I(N__28256));
    LocalMux I__4620 (
            .O(N__28259),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    Odrv4 I__4619 (
            .O(N__28256),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ));
    InMux I__4618 (
            .O(N__28251),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ));
    CascadeMux I__4617 (
            .O(N__28248),
            .I(N__28244));
    CascadeMux I__4616 (
            .O(N__28247),
            .I(N__28241));
    InMux I__4615 (
            .O(N__28244),
            .I(N__28236));
    InMux I__4614 (
            .O(N__28241),
            .I(N__28236));
    LocalMux I__4613 (
            .O(N__28236),
            .I(N__28232));
    InMux I__4612 (
            .O(N__28235),
            .I(N__28229));
    Span4Mux_v I__4611 (
            .O(N__28232),
            .I(N__28226));
    LocalMux I__4610 (
            .O(N__28229),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    Odrv4 I__4609 (
            .O(N__28226),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ));
    InMux I__4608 (
            .O(N__28221),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ));
    InMux I__4607 (
            .O(N__28218),
            .I(N__28212));
    InMux I__4606 (
            .O(N__28217),
            .I(N__28212));
    LocalMux I__4605 (
            .O(N__28212),
            .I(N__28208));
    InMux I__4604 (
            .O(N__28211),
            .I(N__28205));
    Span4Mux_h I__4603 (
            .O(N__28208),
            .I(N__28202));
    LocalMux I__4602 (
            .O(N__28205),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    Odrv4 I__4601 (
            .O(N__28202),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ));
    InMux I__4600 (
            .O(N__28197),
            .I(bfn_11_15_0_));
    InMux I__4599 (
            .O(N__28194),
            .I(N__28187));
    InMux I__4598 (
            .O(N__28193),
            .I(N__28187));
    InMux I__4597 (
            .O(N__28192),
            .I(N__28184));
    LocalMux I__4596 (
            .O(N__28187),
            .I(N__28181));
    LocalMux I__4595 (
            .O(N__28184),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    Odrv4 I__4594 (
            .O(N__28181),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ));
    InMux I__4593 (
            .O(N__28176),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ));
    InMux I__4592 (
            .O(N__28173),
            .I(N__28169));
    InMux I__4591 (
            .O(N__28172),
            .I(N__28166));
    LocalMux I__4590 (
            .O(N__28169),
            .I(N__28163));
    LocalMux I__4589 (
            .O(N__28166),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    Odrv4 I__4588 (
            .O(N__28163),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ));
    InMux I__4587 (
            .O(N__28158),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ));
    InMux I__4586 (
            .O(N__28155),
            .I(N__28151));
    InMux I__4585 (
            .O(N__28154),
            .I(N__28148));
    LocalMux I__4584 (
            .O(N__28151),
            .I(N__28145));
    LocalMux I__4583 (
            .O(N__28148),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    Odrv12 I__4582 (
            .O(N__28145),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ));
    InMux I__4581 (
            .O(N__28140),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ));
    InMux I__4580 (
            .O(N__28137),
            .I(N__28133));
    InMux I__4579 (
            .O(N__28136),
            .I(N__28130));
    LocalMux I__4578 (
            .O(N__28133),
            .I(N__28127));
    LocalMux I__4577 (
            .O(N__28130),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    Odrv4 I__4576 (
            .O(N__28127),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ));
    InMux I__4575 (
            .O(N__28122),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ));
    InMux I__4574 (
            .O(N__28119),
            .I(N__28115));
    InMux I__4573 (
            .O(N__28118),
            .I(N__28112));
    LocalMux I__4572 (
            .O(N__28115),
            .I(N__28109));
    LocalMux I__4571 (
            .O(N__28112),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    Odrv4 I__4570 (
            .O(N__28109),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ));
    InMux I__4569 (
            .O(N__28104),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ));
    InMux I__4568 (
            .O(N__28101),
            .I(N__28097));
    InMux I__4567 (
            .O(N__28100),
            .I(N__28094));
    LocalMux I__4566 (
            .O(N__28097),
            .I(N__28091));
    LocalMux I__4565 (
            .O(N__28094),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    Odrv4 I__4564 (
            .O(N__28091),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ));
    InMux I__4563 (
            .O(N__28086),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ));
    InMux I__4562 (
            .O(N__28083),
            .I(N__28079));
    InMux I__4561 (
            .O(N__28082),
            .I(N__28076));
    LocalMux I__4560 (
            .O(N__28079),
            .I(N__28073));
    LocalMux I__4559 (
            .O(N__28076),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    Odrv12 I__4558 (
            .O(N__28073),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ));
    InMux I__4557 (
            .O(N__28068),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ));
    CascadeMux I__4556 (
            .O(N__28065),
            .I(N__28061));
    CascadeMux I__4555 (
            .O(N__28064),
            .I(N__28058));
    InMux I__4554 (
            .O(N__28061),
            .I(N__28053));
    InMux I__4553 (
            .O(N__28058),
            .I(N__28053));
    LocalMux I__4552 (
            .O(N__28053),
            .I(N__28049));
    InMux I__4551 (
            .O(N__28052),
            .I(N__28046));
    Sp12to4 I__4550 (
            .O(N__28049),
            .I(N__28043));
    LocalMux I__4549 (
            .O(N__28046),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    Odrv12 I__4548 (
            .O(N__28043),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ));
    InMux I__4547 (
            .O(N__28038),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ));
    InMux I__4546 (
            .O(N__28035),
            .I(N__28029));
    InMux I__4545 (
            .O(N__28034),
            .I(N__28029));
    LocalMux I__4544 (
            .O(N__28029),
            .I(N__28025));
    InMux I__4543 (
            .O(N__28028),
            .I(N__28022));
    Span4Mux_v I__4542 (
            .O(N__28025),
            .I(N__28019));
    LocalMux I__4541 (
            .O(N__28022),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    Odrv4 I__4540 (
            .O(N__28019),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ));
    InMux I__4539 (
            .O(N__28014),
            .I(bfn_11_14_0_));
    InMux I__4538 (
            .O(N__28011),
            .I(N__28007));
    InMux I__4537 (
            .O(N__28010),
            .I(N__28004));
    LocalMux I__4536 (
            .O(N__28007),
            .I(N__28001));
    LocalMux I__4535 (
            .O(N__28004),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    Odrv12 I__4534 (
            .O(N__28001),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ));
    InMux I__4533 (
            .O(N__27996),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ));
    CascadeMux I__4532 (
            .O(N__27993),
            .I(N__27989));
    CascadeMux I__4531 (
            .O(N__27992),
            .I(N__27986));
    InMux I__4530 (
            .O(N__27989),
            .I(N__27981));
    InMux I__4529 (
            .O(N__27986),
            .I(N__27981));
    LocalMux I__4528 (
            .O(N__27981),
            .I(\phase_controller_inst1.stoper_tr.N_42_i ));
    InMux I__4527 (
            .O(N__27978),
            .I(N__27974));
    InMux I__4526 (
            .O(N__27977),
            .I(N__27971));
    LocalMux I__4525 (
            .O(N__27974),
            .I(N__27968));
    LocalMux I__4524 (
            .O(N__27971),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    Odrv4 I__4523 (
            .O(N__27968),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ));
    InMux I__4522 (
            .O(N__27963),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ));
    InMux I__4521 (
            .O(N__27960),
            .I(N__27956));
    InMux I__4520 (
            .O(N__27959),
            .I(N__27953));
    LocalMux I__4519 (
            .O(N__27956),
            .I(N__27950));
    LocalMux I__4518 (
            .O(N__27953),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    Odrv4 I__4517 (
            .O(N__27950),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ));
    InMux I__4516 (
            .O(N__27945),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ));
    InMux I__4515 (
            .O(N__27942),
            .I(N__27938));
    InMux I__4514 (
            .O(N__27941),
            .I(N__27935));
    LocalMux I__4513 (
            .O(N__27938),
            .I(N__27932));
    LocalMux I__4512 (
            .O(N__27935),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    Odrv4 I__4511 (
            .O(N__27932),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ));
    InMux I__4510 (
            .O(N__27927),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ));
    InMux I__4509 (
            .O(N__27924),
            .I(N__27920));
    InMux I__4508 (
            .O(N__27923),
            .I(N__27917));
    LocalMux I__4507 (
            .O(N__27920),
            .I(N__27914));
    LocalMux I__4506 (
            .O(N__27917),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    Odrv4 I__4505 (
            .O(N__27914),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ));
    InMux I__4504 (
            .O(N__27909),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ));
    InMux I__4503 (
            .O(N__27906),
            .I(N__27902));
    InMux I__4502 (
            .O(N__27905),
            .I(N__27899));
    LocalMux I__4501 (
            .O(N__27902),
            .I(N__27896));
    LocalMux I__4500 (
            .O(N__27899),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    Odrv12 I__4499 (
            .O(N__27896),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ));
    InMux I__4498 (
            .O(N__27891),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ));
    InMux I__4497 (
            .O(N__27888),
            .I(N__27884));
    InMux I__4496 (
            .O(N__27887),
            .I(N__27881));
    LocalMux I__4495 (
            .O(N__27884),
            .I(N__27878));
    LocalMux I__4494 (
            .O(N__27881),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    Odrv12 I__4493 (
            .O(N__27878),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ));
    InMux I__4492 (
            .O(N__27873),
            .I(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ));
    InMux I__4491 (
            .O(N__27870),
            .I(N__27866));
    InMux I__4490 (
            .O(N__27869),
            .I(N__27863));
    LocalMux I__4489 (
            .O(N__27866),
            .I(N__27860));
    LocalMux I__4488 (
            .O(N__27863),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    Odrv4 I__4487 (
            .O(N__27860),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ));
    InMux I__4486 (
            .O(N__27855),
            .I(bfn_11_13_0_));
    InMux I__4485 (
            .O(N__27852),
            .I(N__27849));
    LocalMux I__4484 (
            .O(N__27849),
            .I(N__27846));
    Span4Mux_v I__4483 (
            .O(N__27846),
            .I(N__27843));
    Odrv4 I__4482 (
            .O(N__27843),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ));
    CascadeMux I__4481 (
            .O(N__27840),
            .I(N__27837));
    InMux I__4480 (
            .O(N__27837),
            .I(N__27834));
    LocalMux I__4479 (
            .O(N__27834),
            .I(N__27831));
    Span4Mux_v I__4478 (
            .O(N__27831),
            .I(N__27828));
    Odrv4 I__4477 (
            .O(N__27828),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt20 ));
    InMux I__4476 (
            .O(N__27825),
            .I(N__27822));
    LocalMux I__4475 (
            .O(N__27822),
            .I(N__27819));
    Span4Mux_v I__4474 (
            .O(N__27819),
            .I(N__27816));
    Odrv4 I__4473 (
            .O(N__27816),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ));
    CascadeMux I__4472 (
            .O(N__27813),
            .I(N__27810));
    InMux I__4471 (
            .O(N__27810),
            .I(N__27807));
    LocalMux I__4470 (
            .O(N__27807),
            .I(N__27804));
    Span4Mux_v I__4469 (
            .O(N__27804),
            .I(N__27801));
    Odrv4 I__4468 (
            .O(N__27801),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt22 ));
    InMux I__4467 (
            .O(N__27798),
            .I(N__27795));
    LocalMux I__4466 (
            .O(N__27795),
            .I(N__27792));
    Odrv12 I__4465 (
            .O(N__27792),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ));
    CascadeMux I__4464 (
            .O(N__27789),
            .I(N__27786));
    InMux I__4463 (
            .O(N__27786),
            .I(N__27783));
    LocalMux I__4462 (
            .O(N__27783),
            .I(N__27780));
    Odrv12 I__4461 (
            .O(N__27780),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt24 ));
    InMux I__4460 (
            .O(N__27777),
            .I(N__27774));
    LocalMux I__4459 (
            .O(N__27774),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ));
    CascadeMux I__4458 (
            .O(N__27771),
            .I(N__27768));
    InMux I__4457 (
            .O(N__27768),
            .I(N__27765));
    LocalMux I__4456 (
            .O(N__27765),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt26 ));
    InMux I__4455 (
            .O(N__27762),
            .I(N__27759));
    LocalMux I__4454 (
            .O(N__27759),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt28 ));
    CascadeMux I__4453 (
            .O(N__27756),
            .I(N__27753));
    InMux I__4452 (
            .O(N__27753),
            .I(N__27750));
    LocalMux I__4451 (
            .O(N__27750),
            .I(N__27747));
    Odrv4 I__4450 (
            .O(N__27747),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ));
    InMux I__4449 (
            .O(N__27744),
            .I(N__27741));
    LocalMux I__4448 (
            .O(N__27741),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt30 ));
    CascadeMux I__4447 (
            .O(N__27738),
            .I(N__27735));
    InMux I__4446 (
            .O(N__27735),
            .I(N__27732));
    LocalMux I__4445 (
            .O(N__27732),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ));
    InMux I__4444 (
            .O(N__27729),
            .I(\phase_controller_inst1.un4_running_cry_30 ));
    InMux I__4443 (
            .O(N__27726),
            .I(N__27720));
    InMux I__4442 (
            .O(N__27725),
            .I(N__27720));
    LocalMux I__4441 (
            .O(N__27720),
            .I(\phase_controller_inst1.un4_running_cry_30_THRU_CO ));
    InMux I__4440 (
            .O(N__27717),
            .I(N__27714));
    LocalMux I__4439 (
            .O(N__27714),
            .I(N__27711));
    Odrv4 I__4438 (
            .O(N__27711),
            .I(\phase_controller_inst1.N_42 ));
    InMux I__4437 (
            .O(N__27708),
            .I(N__27704));
    InMux I__4436 (
            .O(N__27707),
            .I(N__27700));
    LocalMux I__4435 (
            .O(N__27704),
            .I(N__27697));
    InMux I__4434 (
            .O(N__27703),
            .I(N__27694));
    LocalMux I__4433 (
            .O(N__27700),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    Odrv4 I__4432 (
            .O(N__27697),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    LocalMux I__4431 (
            .O(N__27694),
            .I(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ));
    InMux I__4430 (
            .O(N__27687),
            .I(N__27684));
    LocalMux I__4429 (
            .O(N__27684),
            .I(N__27681));
    Span4Mux_h I__4428 (
            .O(N__27681),
            .I(N__27678));
    Odrv4 I__4427 (
            .O(N__27678),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__4426 (
            .O(N__27675),
            .I(N__27672));
    InMux I__4425 (
            .O(N__27672),
            .I(N__27669));
    LocalMux I__4424 (
            .O(N__27669),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ));
    InMux I__4423 (
            .O(N__27666),
            .I(N__27663));
    LocalMux I__4422 (
            .O(N__27663),
            .I(N__27660));
    Span4Mux_h I__4421 (
            .O(N__27660),
            .I(N__27657));
    Odrv4 I__4420 (
            .O(N__27657),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__4419 (
            .O(N__27654),
            .I(N__27651));
    InMux I__4418 (
            .O(N__27651),
            .I(N__27648));
    LocalMux I__4417 (
            .O(N__27648),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ));
    InMux I__4416 (
            .O(N__27645),
            .I(N__27642));
    LocalMux I__4415 (
            .O(N__27642),
            .I(N__27639));
    Odrv12 I__4414 (
            .O(N__27639),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__4413 (
            .O(N__27636),
            .I(N__27633));
    InMux I__4412 (
            .O(N__27633),
            .I(N__27630));
    LocalMux I__4411 (
            .O(N__27630),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ));
    InMux I__4410 (
            .O(N__27627),
            .I(N__27624));
    LocalMux I__4409 (
            .O(N__27624),
            .I(N__27621));
    Span4Mux_v I__4408 (
            .O(N__27621),
            .I(N__27618));
    Odrv4 I__4407 (
            .O(N__27618),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__4406 (
            .O(N__27615),
            .I(N__27612));
    InMux I__4405 (
            .O(N__27612),
            .I(N__27609));
    LocalMux I__4404 (
            .O(N__27609),
            .I(N__27606));
    Odrv4 I__4403 (
            .O(N__27606),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__4402 (
            .O(N__27603),
            .I(N__27600));
    InMux I__4401 (
            .O(N__27600),
            .I(N__27597));
    LocalMux I__4400 (
            .O(N__27597),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ));
    CascadeMux I__4399 (
            .O(N__27594),
            .I(N__27591));
    InMux I__4398 (
            .O(N__27591),
            .I(N__27588));
    LocalMux I__4397 (
            .O(N__27588),
            .I(N__27585));
    Odrv12 I__4396 (
            .O(N__27585),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ));
    InMux I__4395 (
            .O(N__27582),
            .I(N__27579));
    LocalMux I__4394 (
            .O(N__27579),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ));
    InMux I__4393 (
            .O(N__27576),
            .I(N__27573));
    LocalMux I__4392 (
            .O(N__27573),
            .I(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__4391 (
            .O(N__27570),
            .I(N__27567));
    InMux I__4390 (
            .O(N__27567),
            .I(N__27564));
    LocalMux I__4389 (
            .O(N__27564),
            .I(\phase_controller_inst1.stoper_tr.un4_running_lt16 ));
    InMux I__4388 (
            .O(N__27561),
            .I(N__27558));
    LocalMux I__4387 (
            .O(N__27558),
            .I(N__27555));
    Span4Mux_h I__4386 (
            .O(N__27555),
            .I(N__27552));
    Odrv4 I__4385 (
            .O(N__27552),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__4384 (
            .O(N__27549),
            .I(N__27546));
    InMux I__4383 (
            .O(N__27546),
            .I(N__27543));
    LocalMux I__4382 (
            .O(N__27543),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ));
    InMux I__4381 (
            .O(N__27540),
            .I(N__27537));
    LocalMux I__4380 (
            .O(N__27537),
            .I(N__27534));
    Odrv4 I__4379 (
            .O(N__27534),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__4378 (
            .O(N__27531),
            .I(N__27528));
    InMux I__4377 (
            .O(N__27528),
            .I(N__27525));
    LocalMux I__4376 (
            .O(N__27525),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ));
    InMux I__4375 (
            .O(N__27522),
            .I(N__27519));
    LocalMux I__4374 (
            .O(N__27519),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__4373 (
            .O(N__27516),
            .I(N__27513));
    InMux I__4372 (
            .O(N__27513),
            .I(N__27510));
    LocalMux I__4371 (
            .O(N__27510),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ));
    InMux I__4370 (
            .O(N__27507),
            .I(N__27504));
    LocalMux I__4369 (
            .O(N__27504),
            .I(N__27501));
    Span4Mux_v I__4368 (
            .O(N__27501),
            .I(N__27498));
    Odrv4 I__4367 (
            .O(N__27498),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__4366 (
            .O(N__27495),
            .I(N__27492));
    InMux I__4365 (
            .O(N__27492),
            .I(N__27489));
    LocalMux I__4364 (
            .O(N__27489),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ));
    InMux I__4363 (
            .O(N__27486),
            .I(N__27483));
    LocalMux I__4362 (
            .O(N__27483),
            .I(N__27480));
    Odrv4 I__4361 (
            .O(N__27480),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__4360 (
            .O(N__27477),
            .I(N__27474));
    InMux I__4359 (
            .O(N__27474),
            .I(N__27471));
    LocalMux I__4358 (
            .O(N__27471),
            .I(N__27468));
    Odrv4 I__4357 (
            .O(N__27468),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ));
    InMux I__4356 (
            .O(N__27465),
            .I(N__27462));
    LocalMux I__4355 (
            .O(N__27462),
            .I(N__27459));
    Odrv12 I__4354 (
            .O(N__27459),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ));
    CascadeMux I__4353 (
            .O(N__27456),
            .I(N__27453));
    InMux I__4352 (
            .O(N__27453),
            .I(N__27450));
    LocalMux I__4351 (
            .O(N__27450),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ));
    InMux I__4350 (
            .O(N__27447),
            .I(N__27444));
    LocalMux I__4349 (
            .O(N__27444),
            .I(N__27441));
    Odrv4 I__4348 (
            .O(N__27441),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__4347 (
            .O(N__27438),
            .I(N__27435));
    InMux I__4346 (
            .O(N__27435),
            .I(N__27432));
    LocalMux I__4345 (
            .O(N__27432),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ));
    InMux I__4344 (
            .O(N__27429),
            .I(N__27426));
    LocalMux I__4343 (
            .O(N__27426),
            .I(N__27423));
    Odrv12 I__4342 (
            .O(N__27423),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__4341 (
            .O(N__27420),
            .I(N__27417));
    InMux I__4340 (
            .O(N__27417),
            .I(N__27414));
    LocalMux I__4339 (
            .O(N__27414),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ));
    InMux I__4338 (
            .O(N__27411),
            .I(\phase_controller_inst2.un4_running_cry_30 ));
    InMux I__4337 (
            .O(N__27408),
            .I(N__27405));
    LocalMux I__4336 (
            .O(N__27405),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt28 ));
    CascadeMux I__4335 (
            .O(N__27402),
            .I(N__27399));
    InMux I__4334 (
            .O(N__27399),
            .I(N__27393));
    InMux I__4333 (
            .O(N__27398),
            .I(N__27393));
    LocalMux I__4332 (
            .O(N__27393),
            .I(N__27390));
    Odrv12 I__4331 (
            .O(N__27390),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ));
    CascadeMux I__4330 (
            .O(N__27387),
            .I(N__27384));
    InMux I__4329 (
            .O(N__27384),
            .I(N__27381));
    LocalMux I__4328 (
            .O(N__27381),
            .I(N__27378));
    Odrv4 I__4327 (
            .O(N__27378),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ));
    InMux I__4326 (
            .O(N__27375),
            .I(N__27372));
    LocalMux I__4325 (
            .O(N__27372),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ));
    CascadeMux I__4324 (
            .O(N__27369),
            .I(N__27366));
    InMux I__4323 (
            .O(N__27366),
            .I(N__27360));
    InMux I__4322 (
            .O(N__27365),
            .I(N__27360));
    LocalMux I__4321 (
            .O(N__27360),
            .I(N__27357));
    Span4Mux_h I__4320 (
            .O(N__27357),
            .I(N__27354));
    Odrv4 I__4319 (
            .O(N__27354),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ));
    CascadeMux I__4318 (
            .O(N__27351),
            .I(N__27348));
    InMux I__4317 (
            .O(N__27348),
            .I(N__27345));
    LocalMux I__4316 (
            .O(N__27345),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt30 ));
    InMux I__4315 (
            .O(N__27342),
            .I(N__27337));
    InMux I__4314 (
            .O(N__27341),
            .I(N__27334));
    InMux I__4313 (
            .O(N__27340),
            .I(N__27331));
    LocalMux I__4312 (
            .O(N__27337),
            .I(N__27328));
    LocalMux I__4311 (
            .O(N__27334),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    LocalMux I__4310 (
            .O(N__27331),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    Odrv12 I__4309 (
            .O(N__27328),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    InMux I__4308 (
            .O(N__27321),
            .I(N__27318));
    LocalMux I__4307 (
            .O(N__27318),
            .I(N__27313));
    CascadeMux I__4306 (
            .O(N__27317),
            .I(N__27309));
    InMux I__4305 (
            .O(N__27316),
            .I(N__27306));
    Span4Mux_v I__4304 (
            .O(N__27313),
            .I(N__27303));
    InMux I__4303 (
            .O(N__27312),
            .I(N__27298));
    InMux I__4302 (
            .O(N__27309),
            .I(N__27298));
    LocalMux I__4301 (
            .O(N__27306),
            .I(N__27295));
    Span4Mux_h I__4300 (
            .O(N__27303),
            .I(N__27290));
    LocalMux I__4299 (
            .O(N__27298),
            .I(N__27290));
    Span4Mux_h I__4298 (
            .O(N__27295),
            .I(N__27287));
    Span4Mux_v I__4297 (
            .O(N__27290),
            .I(N__27284));
    Odrv4 I__4296 (
            .O(N__27287),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    Odrv4 I__4295 (
            .O(N__27284),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__4294 (
            .O(N__27279),
            .I(N__27273));
    InMux I__4293 (
            .O(N__27278),
            .I(N__27273));
    LocalMux I__4292 (
            .O(N__27273),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ));
    InMux I__4291 (
            .O(N__27270),
            .I(N__27267));
    LocalMux I__4290 (
            .O(N__27267),
            .I(N__27264));
    Odrv12 I__4289 (
            .O(N__27264),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__4288 (
            .O(N__27261),
            .I(N__27258));
    InMux I__4287 (
            .O(N__27258),
            .I(N__27255));
    LocalMux I__4286 (
            .O(N__27255),
            .I(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ));
    InMux I__4285 (
            .O(N__27252),
            .I(N__27249));
    LocalMux I__4284 (
            .O(N__27249),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ));
    CascadeMux I__4283 (
            .O(N__27246),
            .I(N__27243));
    InMux I__4282 (
            .O(N__27243),
            .I(N__27240));
    LocalMux I__4281 (
            .O(N__27240),
            .I(N__27237));
    Odrv4 I__4280 (
            .O(N__27237),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ));
    InMux I__4279 (
            .O(N__27234),
            .I(N__27231));
    LocalMux I__4278 (
            .O(N__27231),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ));
    CascadeMux I__4277 (
            .O(N__27228),
            .I(N__27225));
    InMux I__4276 (
            .O(N__27225),
            .I(N__27222));
    LocalMux I__4275 (
            .O(N__27222),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ));
    InMux I__4274 (
            .O(N__27219),
            .I(N__27216));
    LocalMux I__4273 (
            .O(N__27216),
            .I(N__27213));
    Odrv4 I__4272 (
            .O(N__27213),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ));
    CascadeMux I__4271 (
            .O(N__27210),
            .I(N__27207));
    InMux I__4270 (
            .O(N__27207),
            .I(N__27204));
    LocalMux I__4269 (
            .O(N__27204),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt20 ));
    InMux I__4268 (
            .O(N__27201),
            .I(N__27198));
    LocalMux I__4267 (
            .O(N__27198),
            .I(N__27195));
    Span12Mux_h I__4266 (
            .O(N__27195),
            .I(N__27192));
    Odrv12 I__4265 (
            .O(N__27192),
            .I(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ));
    CascadeMux I__4264 (
            .O(N__27189),
            .I(N__27186));
    InMux I__4263 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__4262 (
            .O(N__27183),
            .I(\phase_controller_inst2.stoper_tr.un4_running_lt22 ));
    InMux I__4261 (
            .O(N__27180),
            .I(N__27177));
    LocalMux I__4260 (
            .O(N__27177),
            .I(N__27174));
    Span4Mux_h I__4259 (
            .O(N__27174),
            .I(N__27171));
    Odrv4 I__4258 (
            .O(N__27171),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ));
    CascadeMux I__4257 (
            .O(N__27168),
            .I(N__27165));
    InMux I__4256 (
            .O(N__27165),
            .I(N__27162));
    LocalMux I__4255 (
            .O(N__27162),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ));
    InMux I__4254 (
            .O(N__27159),
            .I(N__27156));
    LocalMux I__4253 (
            .O(N__27156),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ));
    InMux I__4252 (
            .O(N__27153),
            .I(N__27150));
    LocalMux I__4251 (
            .O(N__27150),
            .I(N__27147));
    Odrv12 I__4250 (
            .O(N__27147),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ));
    CascadeMux I__4249 (
            .O(N__27144),
            .I(N__27141));
    InMux I__4248 (
            .O(N__27141),
            .I(N__27138));
    LocalMux I__4247 (
            .O(N__27138),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ));
    InMux I__4246 (
            .O(N__27135),
            .I(N__27132));
    LocalMux I__4245 (
            .O(N__27132),
            .I(N__27129));
    Span4Mux_h I__4244 (
            .O(N__27129),
            .I(N__27126));
    Odrv4 I__4243 (
            .O(N__27126),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ));
    CascadeMux I__4242 (
            .O(N__27123),
            .I(N__27120));
    InMux I__4241 (
            .O(N__27120),
            .I(N__27117));
    LocalMux I__4240 (
            .O(N__27117),
            .I(N__27114));
    Odrv4 I__4239 (
            .O(N__27114),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ));
    InMux I__4238 (
            .O(N__27111),
            .I(N__27108));
    LocalMux I__4237 (
            .O(N__27108),
            .I(N__27105));
    Span4Mux_h I__4236 (
            .O(N__27105),
            .I(N__27102));
    Odrv4 I__4235 (
            .O(N__27102),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ));
    CascadeMux I__4234 (
            .O(N__27099),
            .I(N__27096));
    InMux I__4233 (
            .O(N__27096),
            .I(N__27093));
    LocalMux I__4232 (
            .O(N__27093),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ));
    InMux I__4231 (
            .O(N__27090),
            .I(N__27087));
    LocalMux I__4230 (
            .O(N__27087),
            .I(N__27084));
    Span4Mux_h I__4229 (
            .O(N__27084),
            .I(N__27081));
    Odrv4 I__4228 (
            .O(N__27081),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ));
    CascadeMux I__4227 (
            .O(N__27078),
            .I(N__27075));
    InMux I__4226 (
            .O(N__27075),
            .I(N__27072));
    LocalMux I__4225 (
            .O(N__27072),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ));
    InMux I__4224 (
            .O(N__27069),
            .I(N__27066));
    LocalMux I__4223 (
            .O(N__27066),
            .I(N__27063));
    Odrv12 I__4222 (
            .O(N__27063),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ));
    CascadeMux I__4221 (
            .O(N__27060),
            .I(N__27057));
    InMux I__4220 (
            .O(N__27057),
            .I(N__27054));
    LocalMux I__4219 (
            .O(N__27054),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ));
    InMux I__4218 (
            .O(N__27051),
            .I(N__27048));
    LocalMux I__4217 (
            .O(N__27048),
            .I(N__27045));
    Odrv12 I__4216 (
            .O(N__27045),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ));
    CascadeMux I__4215 (
            .O(N__27042),
            .I(N__27039));
    InMux I__4214 (
            .O(N__27039),
            .I(N__27036));
    LocalMux I__4213 (
            .O(N__27036),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ));
    CascadeMux I__4212 (
            .O(N__27033),
            .I(N__27030));
    InMux I__4211 (
            .O(N__27030),
            .I(N__27027));
    LocalMux I__4210 (
            .O(N__27027),
            .I(N__27024));
    Odrv4 I__4209 (
            .O(N__27024),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__4208 (
            .O(N__27021),
            .I(N__27018));
    LocalMux I__4207 (
            .O(N__27018),
            .I(N__27015));
    Odrv4 I__4206 (
            .O(N__27015),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__4205 (
            .O(N__27012),
            .I(N__27009));
    LocalMux I__4204 (
            .O(N__27009),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    CascadeMux I__4203 (
            .O(N__27006),
            .I(N__27003));
    InMux I__4202 (
            .O(N__27003),
            .I(N__27000));
    LocalMux I__4201 (
            .O(N__27000),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__4200 (
            .O(N__26997),
            .I(N__26994));
    LocalMux I__4199 (
            .O(N__26994),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ));
    CascadeMux I__4198 (
            .O(N__26991),
            .I(N__26988));
    InMux I__4197 (
            .O(N__26988),
            .I(N__26985));
    LocalMux I__4196 (
            .O(N__26985),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ));
    InMux I__4195 (
            .O(N__26982),
            .I(N__26979));
    LocalMux I__4194 (
            .O(N__26979),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ));
    CascadeMux I__4193 (
            .O(N__26976),
            .I(N__26973));
    InMux I__4192 (
            .O(N__26973),
            .I(N__26970));
    LocalMux I__4191 (
            .O(N__26970),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ));
    InMux I__4190 (
            .O(N__26967),
            .I(N__26964));
    LocalMux I__4189 (
            .O(N__26964),
            .I(N__26961));
    Odrv12 I__4188 (
            .O(N__26961),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ));
    CascadeMux I__4187 (
            .O(N__26958),
            .I(N__26955));
    InMux I__4186 (
            .O(N__26955),
            .I(N__26952));
    LocalMux I__4185 (
            .O(N__26952),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ));
    InMux I__4184 (
            .O(N__26949),
            .I(N__26946));
    LocalMux I__4183 (
            .O(N__26946),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ));
    CascadeMux I__4182 (
            .O(N__26943),
            .I(N__26940));
    InMux I__4181 (
            .O(N__26940),
            .I(N__26937));
    LocalMux I__4180 (
            .O(N__26937),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ));
    InMux I__4179 (
            .O(N__26934),
            .I(N__26931));
    LocalMux I__4178 (
            .O(N__26931),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ));
    CascadeMux I__4177 (
            .O(N__26928),
            .I(N__26925));
    InMux I__4176 (
            .O(N__26925),
            .I(N__26922));
    LocalMux I__4175 (
            .O(N__26922),
            .I(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ));
    CascadeMux I__4174 (
            .O(N__26919),
            .I(N__26916));
    InMux I__4173 (
            .O(N__26916),
            .I(N__26913));
    LocalMux I__4172 (
            .O(N__26913),
            .I(N__26910));
    Span4Mux_h I__4171 (
            .O(N__26910),
            .I(N__26907));
    Odrv4 I__4170 (
            .O(N__26907),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    CascadeMux I__4169 (
            .O(N__26904),
            .I(N__26901));
    InMux I__4168 (
            .O(N__26901),
            .I(N__26898));
    LocalMux I__4167 (
            .O(N__26898),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    CascadeMux I__4166 (
            .O(N__26895),
            .I(N__26892));
    InMux I__4165 (
            .O(N__26892),
            .I(N__26889));
    LocalMux I__4164 (
            .O(N__26889),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    CascadeMux I__4163 (
            .O(N__26886),
            .I(N__26883));
    InMux I__4162 (
            .O(N__26883),
            .I(N__26880));
    LocalMux I__4161 (
            .O(N__26880),
            .I(N__26877));
    Odrv4 I__4160 (
            .O(N__26877),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    CascadeMux I__4159 (
            .O(N__26874),
            .I(N__26871));
    InMux I__4158 (
            .O(N__26871),
            .I(N__26868));
    LocalMux I__4157 (
            .O(N__26868),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__4156 (
            .O(N__26865),
            .I(N__26862));
    LocalMux I__4155 (
            .O(N__26862),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__4154 (
            .O(N__26859),
            .I(N__26856));
    LocalMux I__4153 (
            .O(N__26856),
            .I(N__26853));
    Odrv12 I__4152 (
            .O(N__26853),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__4151 (
            .O(N__26850),
            .I(N__26847));
    LocalMux I__4150 (
            .O(N__26847),
            .I(N__26844));
    Span4Mux_h I__4149 (
            .O(N__26844),
            .I(N__26841));
    Odrv4 I__4148 (
            .O(N__26841),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__4147 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__4146 (
            .O(N__26835),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__4145 (
            .O(N__26832),
            .I(N__26829));
    LocalMux I__4144 (
            .O(N__26829),
            .I(N__26826));
    Odrv12 I__4143 (
            .O(N__26826),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__4142 (
            .O(N__26823),
            .I(N__26820));
    LocalMux I__4141 (
            .O(N__26820),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__4140 (
            .O(N__26817),
            .I(N__26814));
    LocalMux I__4139 (
            .O(N__26814),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    CascadeMux I__4138 (
            .O(N__26811),
            .I(N__26808));
    InMux I__4137 (
            .O(N__26808),
            .I(N__26805));
    LocalMux I__4136 (
            .O(N__26805),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    CascadeMux I__4135 (
            .O(N__26802),
            .I(N__26799));
    InMux I__4134 (
            .O(N__26799),
            .I(N__26796));
    LocalMux I__4133 (
            .O(N__26796),
            .I(N__26793));
    Odrv4 I__4132 (
            .O(N__26793),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__4131 (
            .O(N__26790),
            .I(N__26787));
    LocalMux I__4130 (
            .O(N__26787),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__4129 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__4128 (
            .O(N__26781),
            .I(N__26778));
    Odrv4 I__4127 (
            .O(N__26778),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__4126 (
            .O(N__26775),
            .I(N__26772));
    LocalMux I__4125 (
            .O(N__26772),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__4124 (
            .O(N__26769),
            .I(N__26766));
    LocalMux I__4123 (
            .O(N__26766),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__4122 (
            .O(N__26763),
            .I(N__26760));
    LocalMux I__4121 (
            .O(N__26760),
            .I(N__26757));
    Odrv4 I__4120 (
            .O(N__26757),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__4119 (
            .O(N__26754),
            .I(N__26751));
    LocalMux I__4118 (
            .O(N__26751),
            .I(N__26748));
    Odrv4 I__4117 (
            .O(N__26748),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__4116 (
            .O(N__26745),
            .I(N__26742));
    LocalMux I__4115 (
            .O(N__26742),
            .I(N__26739));
    Odrv4 I__4114 (
            .O(N__26739),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    CascadeMux I__4113 (
            .O(N__26736),
            .I(N__26733));
    InMux I__4112 (
            .O(N__26733),
            .I(N__26730));
    LocalMux I__4111 (
            .O(N__26730),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    InMux I__4110 (
            .O(N__26727),
            .I(N__26724));
    LocalMux I__4109 (
            .O(N__26724),
            .I(N__26721));
    Span4Mux_h I__4108 (
            .O(N__26721),
            .I(N__26718));
    Odrv4 I__4107 (
            .O(N__26718),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__4106 (
            .O(N__26715),
            .I(N__26712));
    LocalMux I__4105 (
            .O(N__26712),
            .I(N__26709));
    Odrv4 I__4104 (
            .O(N__26709),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    CascadeMux I__4103 (
            .O(N__26706),
            .I(N__26703));
    InMux I__4102 (
            .O(N__26703),
            .I(N__26700));
    LocalMux I__4101 (
            .O(N__26700),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    InMux I__4100 (
            .O(N__26697),
            .I(N__26694));
    LocalMux I__4099 (
            .O(N__26694),
            .I(N__26691));
    Span4Mux_v I__4098 (
            .O(N__26691),
            .I(N__26688));
    Odrv4 I__4097 (
            .O(N__26688),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__4096 (
            .O(N__26685),
            .I(N__26682));
    LocalMux I__4095 (
            .O(N__26682),
            .I(N__26679));
    Span4Mux_v I__4094 (
            .O(N__26679),
            .I(N__26676));
    Odrv4 I__4093 (
            .O(N__26676),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__4092 (
            .O(N__26673),
            .I(N__26670));
    LocalMux I__4091 (
            .O(N__26670),
            .I(N__26667));
    Odrv4 I__4090 (
            .O(N__26667),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    InMux I__4089 (
            .O(N__26664),
            .I(N__26661));
    LocalMux I__4088 (
            .O(N__26661),
            .I(N__26658));
    Sp12to4 I__4087 (
            .O(N__26658),
            .I(N__26655));
    Odrv12 I__4086 (
            .O(N__26655),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    CascadeMux I__4085 (
            .O(N__26652),
            .I(N__26649));
    InMux I__4084 (
            .O(N__26649),
            .I(N__26646));
    LocalMux I__4083 (
            .O(N__26646),
            .I(N__26643));
    Span4Mux_h I__4082 (
            .O(N__26643),
            .I(N__26640));
    Span4Mux_v I__4081 (
            .O(N__26640),
            .I(N__26637));
    Odrv4 I__4080 (
            .O(N__26637),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    CascadeMux I__4079 (
            .O(N__26634),
            .I(N__26631));
    InMux I__4078 (
            .O(N__26631),
            .I(N__26628));
    LocalMux I__4077 (
            .O(N__26628),
            .I(N__26625));
    Odrv4 I__4076 (
            .O(N__26625),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__4075 (
            .O(N__26622),
            .I(N__26619));
    LocalMux I__4074 (
            .O(N__26619),
            .I(N__26616));
    Span12Mux_v I__4073 (
            .O(N__26616),
            .I(N__26613));
    Odrv12 I__4072 (
            .O(N__26613),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__4071 (
            .O(N__26610),
            .I(N__26606));
    InMux I__4070 (
            .O(N__26609),
            .I(N__26601));
    LocalMux I__4069 (
            .O(N__26606),
            .I(N__26598));
    InMux I__4068 (
            .O(N__26605),
            .I(N__26593));
    InMux I__4067 (
            .O(N__26604),
            .I(N__26593));
    LocalMux I__4066 (
            .O(N__26601),
            .I(N__26590));
    Span4Mux_h I__4065 (
            .O(N__26598),
            .I(N__26587));
    LocalMux I__4064 (
            .O(N__26593),
            .I(N__26584));
    Span4Mux_v I__4063 (
            .O(N__26590),
            .I(N__26581));
    Odrv4 I__4062 (
            .O(N__26587),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv12 I__4061 (
            .O(N__26584),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    Odrv4 I__4060 (
            .O(N__26581),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    CascadeMux I__4059 (
            .O(N__26574),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_));
    InMux I__4058 (
            .O(N__26571),
            .I(N__26565));
    InMux I__4057 (
            .O(N__26570),
            .I(N__26565));
    LocalMux I__4056 (
            .O(N__26565),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ));
    InMux I__4055 (
            .O(N__26562),
            .I(N__26558));
    InMux I__4054 (
            .O(N__26561),
            .I(N__26555));
    LocalMux I__4053 (
            .O(N__26558),
            .I(N__26550));
    LocalMux I__4052 (
            .O(N__26555),
            .I(N__26550));
    Odrv4 I__4051 (
            .O(N__26550),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ));
    CascadeMux I__4050 (
            .O(N__26547),
            .I(N__26543));
    CascadeMux I__4049 (
            .O(N__26546),
            .I(N__26540));
    InMux I__4048 (
            .O(N__26543),
            .I(N__26537));
    InMux I__4047 (
            .O(N__26540),
            .I(N__26534));
    LocalMux I__4046 (
            .O(N__26537),
            .I(N__26531));
    LocalMux I__4045 (
            .O(N__26534),
            .I(N__26528));
    Span4Mux_h I__4044 (
            .O(N__26531),
            .I(N__26525));
    Span4Mux_v I__4043 (
            .O(N__26528),
            .I(N__26522));
    Span4Mux_v I__4042 (
            .O(N__26525),
            .I(N__26519));
    Odrv4 I__4041 (
            .O(N__26522),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    Odrv4 I__4040 (
            .O(N__26519),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ));
    CascadeMux I__4039 (
            .O(N__26514),
            .I(N__26511));
    InMux I__4038 (
            .O(N__26511),
            .I(N__26508));
    LocalMux I__4037 (
            .O(N__26508),
            .I(N__26505));
    Span4Mux_h I__4036 (
            .O(N__26505),
            .I(N__26502));
    Span4Mux_v I__4035 (
            .O(N__26502),
            .I(N__26499));
    Odrv4 I__4034 (
            .O(N__26499),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    CascadeMux I__4033 (
            .O(N__26496),
            .I(N__26493));
    InMux I__4032 (
            .O(N__26493),
            .I(N__26490));
    LocalMux I__4031 (
            .O(N__26490),
            .I(N__26487));
    Span4Mux_v I__4030 (
            .O(N__26487),
            .I(N__26484));
    Odrv4 I__4029 (
            .O(N__26484),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    CascadeMux I__4028 (
            .O(N__26481),
            .I(N__26478));
    InMux I__4027 (
            .O(N__26478),
            .I(N__26475));
    LocalMux I__4026 (
            .O(N__26475),
            .I(N__26472));
    Span4Mux_v I__4025 (
            .O(N__26472),
            .I(N__26469));
    Odrv4 I__4024 (
            .O(N__26469),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    CascadeMux I__4023 (
            .O(N__26466),
            .I(N__26463));
    InMux I__4022 (
            .O(N__26463),
            .I(N__26460));
    LocalMux I__4021 (
            .O(N__26460),
            .I(N__26457));
    Span4Mux_v I__4020 (
            .O(N__26457),
            .I(N__26454));
    Odrv4 I__4019 (
            .O(N__26454),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    CascadeMux I__4018 (
            .O(N__26451),
            .I(N__26448));
    InMux I__4017 (
            .O(N__26448),
            .I(N__26445));
    LocalMux I__4016 (
            .O(N__26445),
            .I(N__26442));
    Span4Mux_v I__4015 (
            .O(N__26442),
            .I(N__26439));
    Odrv4 I__4014 (
            .O(N__26439),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__4013 (
            .O(N__26436),
            .I(N__26433));
    LocalMux I__4012 (
            .O(N__26433),
            .I(N__26430));
    Span4Mux_v I__4011 (
            .O(N__26430),
            .I(N__26427));
    Odrv4 I__4010 (
            .O(N__26427),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    CascadeMux I__4009 (
            .O(N__26424),
            .I(\phase_controller_inst1.N_42_cascade_ ));
    CascadeMux I__4008 (
            .O(N__26421),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_));
    InMux I__4007 (
            .O(N__26418),
            .I(N__26412));
    InMux I__4006 (
            .O(N__26417),
            .I(N__26412));
    LocalMux I__4005 (
            .O(N__26412),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ));
    CascadeMux I__4004 (
            .O(N__26409),
            .I(N__26405));
    CascadeMux I__4003 (
            .O(N__26408),
            .I(N__26402));
    InMux I__4002 (
            .O(N__26405),
            .I(N__26397));
    InMux I__4001 (
            .O(N__26402),
            .I(N__26397));
    LocalMux I__4000 (
            .O(N__26397),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ));
    InMux I__3999 (
            .O(N__26394),
            .I(N__26390));
    InMux I__3998 (
            .O(N__26393),
            .I(N__26386));
    LocalMux I__3997 (
            .O(N__26390),
            .I(N__26383));
    InMux I__3996 (
            .O(N__26389),
            .I(N__26380));
    LocalMux I__3995 (
            .O(N__26386),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    Odrv12 I__3994 (
            .O(N__26383),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    LocalMux I__3993 (
            .O(N__26380),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    InMux I__3992 (
            .O(N__26373),
            .I(N__26370));
    LocalMux I__3991 (
            .O(N__26370),
            .I(N__26364));
    InMux I__3990 (
            .O(N__26369),
            .I(N__26361));
    InMux I__3989 (
            .O(N__26368),
            .I(N__26358));
    InMux I__3988 (
            .O(N__26367),
            .I(N__26355));
    Span4Mux_v I__3987 (
            .O(N__26364),
            .I(N__26350));
    LocalMux I__3986 (
            .O(N__26361),
            .I(N__26350));
    LocalMux I__3985 (
            .O(N__26358),
            .I(N__26347));
    LocalMux I__3984 (
            .O(N__26355),
            .I(N__26344));
    Span4Mux_v I__3983 (
            .O(N__26350),
            .I(N__26341));
    Span4Mux_h I__3982 (
            .O(N__26347),
            .I(N__26336));
    Span4Mux_v I__3981 (
            .O(N__26344),
            .I(N__26336));
    Odrv4 I__3980 (
            .O(N__26341),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    Odrv4 I__3979 (
            .O(N__26336),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    CascadeMux I__3978 (
            .O(N__26331),
            .I(N__26328));
    InMux I__3977 (
            .O(N__26328),
            .I(N__26322));
    InMux I__3976 (
            .O(N__26327),
            .I(N__26322));
    LocalMux I__3975 (
            .O(N__26322),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ));
    InMux I__3974 (
            .O(N__26319),
            .I(N__26315));
    InMux I__3973 (
            .O(N__26318),
            .I(N__26312));
    LocalMux I__3972 (
            .O(N__26315),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    LocalMux I__3971 (
            .O(N__26312),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__3970 (
            .O(N__26307),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_));
    InMux I__3969 (
            .O(N__26304),
            .I(N__26298));
    InMux I__3968 (
            .O(N__26303),
            .I(N__26298));
    LocalMux I__3967 (
            .O(N__26298),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ));
    InMux I__3966 (
            .O(N__26295),
            .I(N__26289));
    InMux I__3965 (
            .O(N__26294),
            .I(N__26289));
    LocalMux I__3964 (
            .O(N__26289),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ));
    InMux I__3963 (
            .O(N__26286),
            .I(N__26283));
    LocalMux I__3962 (
            .O(N__26283),
            .I(\phase_controller_inst1.N_43 ));
    CascadeMux I__3961 (
            .O(N__26280),
            .I(\phase_controller_inst1.N_43_cascade_ ));
    CEMux I__3960 (
            .O(N__26277),
            .I(N__26274));
    LocalMux I__3959 (
            .O(N__26274),
            .I(N__26271));
    Odrv12 I__3958 (
            .O(N__26271),
            .I(\phase_controller_inst1.stoper_tr.N_43_0 ));
    CascadeMux I__3957 (
            .O(N__26268),
            .I(N__26263));
    CascadeMux I__3956 (
            .O(N__26267),
            .I(N__26260));
    InMux I__3955 (
            .O(N__26266),
            .I(N__26253));
    InMux I__3954 (
            .O(N__26263),
            .I(N__26253));
    InMux I__3953 (
            .O(N__26260),
            .I(N__26253));
    LocalMux I__3952 (
            .O(N__26253),
            .I(\phase_controller_inst1.running ));
    InMux I__3951 (
            .O(N__26250),
            .I(N__26247));
    LocalMux I__3950 (
            .O(N__26247),
            .I(N__26242));
    InMux I__3949 (
            .O(N__26246),
            .I(N__26239));
    InMux I__3948 (
            .O(N__26245),
            .I(N__26236));
    Span4Mux_v I__3947 (
            .O(N__26242),
            .I(N__26233));
    LocalMux I__3946 (
            .O(N__26239),
            .I(N__26230));
    LocalMux I__3945 (
            .O(N__26236),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv4 I__3944 (
            .O(N__26233),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    Odrv12 I__3943 (
            .O(N__26230),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__3942 (
            .O(N__26223),
            .I(N__26219));
    InMux I__3941 (
            .O(N__26222),
            .I(N__26216));
    LocalMux I__3940 (
            .O(N__26219),
            .I(N__26211));
    LocalMux I__3939 (
            .O(N__26216),
            .I(N__26208));
    InMux I__3938 (
            .O(N__26215),
            .I(N__26203));
    InMux I__3937 (
            .O(N__26214),
            .I(N__26203));
    Span4Mux_h I__3936 (
            .O(N__26211),
            .I(N__26200));
    Span4Mux_h I__3935 (
            .O(N__26208),
            .I(N__26197));
    LocalMux I__3934 (
            .O(N__26203),
            .I(N__26194));
    Odrv4 I__3933 (
            .O(N__26200),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv4 I__3932 (
            .O(N__26197),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    Odrv12 I__3931 (
            .O(N__26194),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    InMux I__3930 (
            .O(N__26187),
            .I(N__26184));
    LocalMux I__3929 (
            .O(N__26184),
            .I(N__26180));
    InMux I__3928 (
            .O(N__26183),
            .I(N__26177));
    Odrv4 I__3927 (
            .O(N__26180),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__3926 (
            .O(N__26177),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__3925 (
            .O(N__26172),
            .I(N__26169));
    LocalMux I__3924 (
            .O(N__26169),
            .I(N__26164));
    InMux I__3923 (
            .O(N__26168),
            .I(N__26159));
    InMux I__3922 (
            .O(N__26167),
            .I(N__26159));
    Span4Mux_v I__3921 (
            .O(N__26164),
            .I(N__26153));
    LocalMux I__3920 (
            .O(N__26159),
            .I(N__26153));
    InMux I__3919 (
            .O(N__26158),
            .I(N__26150));
    Span4Mux_h I__3918 (
            .O(N__26153),
            .I(N__26147));
    LocalMux I__3917 (
            .O(N__26150),
            .I(N__26144));
    Odrv4 I__3916 (
            .O(N__26147),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    Odrv12 I__3915 (
            .O(N__26144),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    CascadeMux I__3914 (
            .O(N__26139),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_));
    CascadeMux I__3913 (
            .O(N__26136),
            .I(N__26133));
    InMux I__3912 (
            .O(N__26133),
            .I(N__26127));
    InMux I__3911 (
            .O(N__26132),
            .I(N__26127));
    LocalMux I__3910 (
            .O(N__26127),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ));
    InMux I__3909 (
            .O(N__26124),
            .I(N__26121));
    LocalMux I__3908 (
            .O(N__26121),
            .I(N__26117));
    InMux I__3907 (
            .O(N__26120),
            .I(N__26114));
    Odrv4 I__3906 (
            .O(N__26117),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__3905 (
            .O(N__26114),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__3904 (
            .O(N__26109),
            .I(N__26104));
    InMux I__3903 (
            .O(N__26108),
            .I(N__26099));
    InMux I__3902 (
            .O(N__26107),
            .I(N__26099));
    LocalMux I__3901 (
            .O(N__26104),
            .I(N__26096));
    LocalMux I__3900 (
            .O(N__26099),
            .I(N__26092));
    Span4Mux_h I__3899 (
            .O(N__26096),
            .I(N__26089));
    InMux I__3898 (
            .O(N__26095),
            .I(N__26086));
    Span4Mux_h I__3897 (
            .O(N__26092),
            .I(N__26083));
    Sp12to4 I__3896 (
            .O(N__26089),
            .I(N__26078));
    LocalMux I__3895 (
            .O(N__26086),
            .I(N__26078));
    Odrv4 I__3894 (
            .O(N__26083),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    Odrv12 I__3893 (
            .O(N__26078),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    CascadeMux I__3892 (
            .O(N__26073),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_));
    InMux I__3891 (
            .O(N__26070),
            .I(N__26064));
    InMux I__3890 (
            .O(N__26069),
            .I(N__26064));
    LocalMux I__3889 (
            .O(N__26064),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ));
    InMux I__3888 (
            .O(N__26061),
            .I(N__26058));
    LocalMux I__3887 (
            .O(N__26058),
            .I(N__26054));
    InMux I__3886 (
            .O(N__26057),
            .I(N__26051));
    Span4Mux_v I__3885 (
            .O(N__26054),
            .I(N__26047));
    LocalMux I__3884 (
            .O(N__26051),
            .I(N__26044));
    InMux I__3883 (
            .O(N__26050),
            .I(N__26041));
    Span4Mux_h I__3882 (
            .O(N__26047),
            .I(N__26036));
    Span4Mux_h I__3881 (
            .O(N__26044),
            .I(N__26036));
    LocalMux I__3880 (
            .O(N__26041),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    Odrv4 I__3879 (
            .O(N__26036),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__3878 (
            .O(N__26031),
            .I(N__26028));
    LocalMux I__3877 (
            .O(N__26028),
            .I(N__26024));
    InMux I__3876 (
            .O(N__26027),
            .I(N__26021));
    Span4Mux_v I__3875 (
            .O(N__26024),
            .I(N__26015));
    LocalMux I__3874 (
            .O(N__26021),
            .I(N__26015));
    InMux I__3873 (
            .O(N__26020),
            .I(N__26012));
    Span4Mux_h I__3872 (
            .O(N__26015),
            .I(N__26008));
    LocalMux I__3871 (
            .O(N__26012),
            .I(N__26005));
    InMux I__3870 (
            .O(N__26011),
            .I(N__26002));
    Odrv4 I__3869 (
            .O(N__26008),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    Odrv12 I__3868 (
            .O(N__26005),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__3867 (
            .O(N__26002),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__3866 (
            .O(N__25995),
            .I(N__25992));
    LocalMux I__3865 (
            .O(N__25992),
            .I(N__25988));
    InMux I__3864 (
            .O(N__25991),
            .I(N__25984));
    Span4Mux_v I__3863 (
            .O(N__25988),
            .I(N__25981));
    InMux I__3862 (
            .O(N__25987),
            .I(N__25978));
    LocalMux I__3861 (
            .O(N__25984),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    Odrv4 I__3860 (
            .O(N__25981),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    LocalMux I__3859 (
            .O(N__25978),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__3858 (
            .O(N__25971),
            .I(N__25967));
    InMux I__3857 (
            .O(N__25970),
            .I(N__25963));
    LocalMux I__3856 (
            .O(N__25967),
            .I(N__25960));
    InMux I__3855 (
            .O(N__25966),
            .I(N__25957));
    LocalMux I__3854 (
            .O(N__25963),
            .I(N__25953));
    Span4Mux_h I__3853 (
            .O(N__25960),
            .I(N__25950));
    LocalMux I__3852 (
            .O(N__25957),
            .I(N__25947));
    CascadeMux I__3851 (
            .O(N__25956),
            .I(N__25944));
    Span4Mux_v I__3850 (
            .O(N__25953),
            .I(N__25937));
    Span4Mux_v I__3849 (
            .O(N__25950),
            .I(N__25937));
    Span4Mux_v I__3848 (
            .O(N__25947),
            .I(N__25937));
    InMux I__3847 (
            .O(N__25944),
            .I(N__25934));
    Odrv4 I__3846 (
            .O(N__25937),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    LocalMux I__3845 (
            .O(N__25934),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__3844 (
            .O(N__25929),
            .I(N__25923));
    InMux I__3843 (
            .O(N__25928),
            .I(N__25923));
    LocalMux I__3842 (
            .O(N__25923),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ));
    CascadeMux I__3841 (
            .O(N__25920),
            .I(N__25917));
    InMux I__3840 (
            .O(N__25917),
            .I(N__25911));
    InMux I__3839 (
            .O(N__25916),
            .I(N__25911));
    LocalMux I__3838 (
            .O(N__25911),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ));
    InMux I__3837 (
            .O(N__25908),
            .I(N__25903));
    InMux I__3836 (
            .O(N__25907),
            .I(N__25900));
    InMux I__3835 (
            .O(N__25906),
            .I(N__25897));
    LocalMux I__3834 (
            .O(N__25903),
            .I(N__25891));
    LocalMux I__3833 (
            .O(N__25900),
            .I(N__25891));
    LocalMux I__3832 (
            .O(N__25897),
            .I(N__25888));
    InMux I__3831 (
            .O(N__25896),
            .I(N__25885));
    Span4Mux_h I__3830 (
            .O(N__25891),
            .I(N__25882));
    Span4Mux_v I__3829 (
            .O(N__25888),
            .I(N__25877));
    LocalMux I__3828 (
            .O(N__25885),
            .I(N__25877));
    Odrv4 I__3827 (
            .O(N__25882),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    Odrv4 I__3826 (
            .O(N__25877),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__3825 (
            .O(N__25872),
            .I(N__25868));
    InMux I__3824 (
            .O(N__25871),
            .I(N__25864));
    LocalMux I__3823 (
            .O(N__25868),
            .I(N__25861));
    InMux I__3822 (
            .O(N__25867),
            .I(N__25858));
    LocalMux I__3821 (
            .O(N__25864),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    Odrv12 I__3820 (
            .O(N__25861),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    LocalMux I__3819 (
            .O(N__25858),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    InMux I__3818 (
            .O(N__25851),
            .I(N__25845));
    InMux I__3817 (
            .O(N__25850),
            .I(N__25845));
    LocalMux I__3816 (
            .O(N__25845),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__3815 (
            .O(N__25842),
            .I(N__25839));
    InMux I__3814 (
            .O(N__25839),
            .I(N__25833));
    InMux I__3813 (
            .O(N__25838),
            .I(N__25833));
    LocalMux I__3812 (
            .O(N__25833),
            .I(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ));
    InMux I__3811 (
            .O(N__25830),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    InMux I__3810 (
            .O(N__25827),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__3809 (
            .O(N__25824),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    InMux I__3808 (
            .O(N__25821),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    InMux I__3807 (
            .O(N__25818),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__3806 (
            .O(N__25815),
            .I(N__25812));
    LocalMux I__3805 (
            .O(N__25812),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__3804 (
            .O(N__25809),
            .I(N__25806));
    LocalMux I__3803 (
            .O(N__25806),
            .I(N__25803));
    Glb2LocalMux I__3802 (
            .O(N__25803),
            .I(N__25800));
    GlobalMux I__3801 (
            .O(N__25800),
            .I(clk_12mhz));
    IoInMux I__3800 (
            .O(N__25797),
            .I(N__25794));
    LocalMux I__3799 (
            .O(N__25794),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__3798 (
            .O(N__25791),
            .I(N__25788));
    LocalMux I__3797 (
            .O(N__25788),
            .I(N__25783));
    InMux I__3796 (
            .O(N__25787),
            .I(N__25780));
    InMux I__3795 (
            .O(N__25786),
            .I(N__25777));
    Span4Mux_v I__3794 (
            .O(N__25783),
            .I(N__25774));
    LocalMux I__3793 (
            .O(N__25780),
            .I(N__25771));
    LocalMux I__3792 (
            .O(N__25777),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__3791 (
            .O(N__25774),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__3790 (
            .O(N__25771),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__3789 (
            .O(N__25764),
            .I(N__25759));
    InMux I__3788 (
            .O(N__25763),
            .I(N__25756));
    InMux I__3787 (
            .O(N__25762),
            .I(N__25753));
    LocalMux I__3786 (
            .O(N__25759),
            .I(N__25748));
    LocalMux I__3785 (
            .O(N__25756),
            .I(N__25748));
    LocalMux I__3784 (
            .O(N__25753),
            .I(N__25744));
    Span4Mux_h I__3783 (
            .O(N__25748),
            .I(N__25741));
    InMux I__3782 (
            .O(N__25747),
            .I(N__25738));
    Span4Mux_h I__3781 (
            .O(N__25744),
            .I(N__25731));
    Span4Mux_v I__3780 (
            .O(N__25741),
            .I(N__25731));
    LocalMux I__3779 (
            .O(N__25738),
            .I(N__25731));
    Odrv4 I__3778 (
            .O(N__25731),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    CascadeMux I__3777 (
            .O(N__25728),
            .I(N__25725));
    InMux I__3776 (
            .O(N__25725),
            .I(N__25721));
    InMux I__3775 (
            .O(N__25724),
            .I(N__25718));
    LocalMux I__3774 (
            .O(N__25721),
            .I(N__25715));
    LocalMux I__3773 (
            .O(N__25718),
            .I(N__25709));
    Span4Mux_v I__3772 (
            .O(N__25715),
            .I(N__25709));
    InMux I__3771 (
            .O(N__25714),
            .I(N__25706));
    Span4Mux_v I__3770 (
            .O(N__25709),
            .I(N__25703));
    LocalMux I__3769 (
            .O(N__25706),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    Odrv4 I__3768 (
            .O(N__25703),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__3767 (
            .O(N__25698),
            .I(N__25692));
    CascadeMux I__3766 (
            .O(N__25697),
            .I(N__25689));
    InMux I__3765 (
            .O(N__25696),
            .I(N__25686));
    InMux I__3764 (
            .O(N__25695),
            .I(N__25683));
    LocalMux I__3763 (
            .O(N__25692),
            .I(N__25680));
    InMux I__3762 (
            .O(N__25689),
            .I(N__25677));
    LocalMux I__3761 (
            .O(N__25686),
            .I(N__25674));
    LocalMux I__3760 (
            .O(N__25683),
            .I(N__25671));
    Span4Mux_v I__3759 (
            .O(N__25680),
            .I(N__25666));
    LocalMux I__3758 (
            .O(N__25677),
            .I(N__25666));
    Span4Mux_h I__3757 (
            .O(N__25674),
            .I(N__25663));
    Span12Mux_h I__3756 (
            .O(N__25671),
            .I(N__25660));
    Span4Mux_v I__3755 (
            .O(N__25666),
            .I(N__25657));
    Odrv4 I__3754 (
            .O(N__25663),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv12 I__3753 (
            .O(N__25660),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    Odrv4 I__3752 (
            .O(N__25657),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__3751 (
            .O(N__25650),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    InMux I__3750 (
            .O(N__25647),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    InMux I__3749 (
            .O(N__25644),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    InMux I__3748 (
            .O(N__25641),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    CascadeMux I__3747 (
            .O(N__25638),
            .I(N__25635));
    InMux I__3746 (
            .O(N__25635),
            .I(N__25632));
    LocalMux I__3745 (
            .O(N__25632),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__3744 (
            .O(N__25629),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    InMux I__3743 (
            .O(N__25626),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    InMux I__3742 (
            .O(N__25623),
            .I(bfn_9_21_0_));
    InMux I__3741 (
            .O(N__25620),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    InMux I__3740 (
            .O(N__25617),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__3739 (
            .O(N__25614),
            .I(N__25611));
    LocalMux I__3738 (
            .O(N__25611),
            .I(N__25608));
    Odrv12 I__3737 (
            .O(N__25608),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__3736 (
            .O(N__25605),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    InMux I__3735 (
            .O(N__25602),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__3734 (
            .O(N__25599),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    InMux I__3733 (
            .O(N__25596),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__3732 (
            .O(N__25593),
            .I(N__25590));
    LocalMux I__3731 (
            .O(N__25590),
            .I(N__25587));
    Odrv4 I__3730 (
            .O(N__25587),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__3729 (
            .O(N__25584),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    InMux I__3728 (
            .O(N__25581),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__3727 (
            .O(N__25578),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__3726 (
            .O(N__25575),
            .I(bfn_9_20_0_));
    InMux I__3725 (
            .O(N__25572),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    CascadeMux I__3724 (
            .O(N__25569),
            .I(N__25566));
    InMux I__3723 (
            .O(N__25566),
            .I(N__25562));
    InMux I__3722 (
            .O(N__25565),
            .I(N__25559));
    LocalMux I__3721 (
            .O(N__25562),
            .I(N__25556));
    LocalMux I__3720 (
            .O(N__25559),
            .I(N__25553));
    Odrv4 I__3719 (
            .O(N__25556),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    Odrv4 I__3718 (
            .O(N__25553),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__3717 (
            .O(N__25548),
            .I(N__25545));
    InMux I__3716 (
            .O(N__25545),
            .I(N__25541));
    InMux I__3715 (
            .O(N__25544),
            .I(N__25538));
    LocalMux I__3714 (
            .O(N__25541),
            .I(N__25535));
    LocalMux I__3713 (
            .O(N__25538),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__3712 (
            .O(N__25535),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    InMux I__3711 (
            .O(N__25530),
            .I(N__25527));
    LocalMux I__3710 (
            .O(N__25527),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    InMux I__3709 (
            .O(N__25524),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__3708 (
            .O(N__25521),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__3707 (
            .O(N__25518),
            .I(N__25515));
    LocalMux I__3706 (
            .O(N__25515),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    InMux I__3705 (
            .O(N__25512),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    CascadeMux I__3704 (
            .O(N__25509),
            .I(N__25506));
    InMux I__3703 (
            .O(N__25506),
            .I(N__25503));
    LocalMux I__3702 (
            .O(N__25503),
            .I(N__25500));
    Odrv12 I__3701 (
            .O(N__25500),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__3700 (
            .O(N__25497),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    InMux I__3699 (
            .O(N__25494),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    InMux I__3698 (
            .O(N__25491),
            .I(bfn_9_19_0_));
    CascadeMux I__3697 (
            .O(N__25488),
            .I(N__25485));
    InMux I__3696 (
            .O(N__25485),
            .I(N__25482));
    LocalMux I__3695 (
            .O(N__25482),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    CascadeMux I__3694 (
            .O(N__25479),
            .I(N__25476));
    InMux I__3693 (
            .O(N__25476),
            .I(N__25473));
    LocalMux I__3692 (
            .O(N__25473),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__3691 (
            .O(N__25470),
            .I(N__25467));
    LocalMux I__3690 (
            .O(N__25467),
            .I(N__25464));
    Odrv4 I__3689 (
            .O(N__25464),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__3688 (
            .O(N__25461),
            .I(N__25458));
    LocalMux I__3687 (
            .O(N__25458),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__3686 (
            .O(N__25455),
            .I(N__25452));
    LocalMux I__3685 (
            .O(N__25452),
            .I(N__25449));
    Odrv4 I__3684 (
            .O(N__25449),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__3683 (
            .O(N__25446),
            .I(N__25443));
    LocalMux I__3682 (
            .O(N__25443),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    CascadeMux I__3681 (
            .O(N__25440),
            .I(N__25437));
    InMux I__3680 (
            .O(N__25437),
            .I(N__25434));
    LocalMux I__3679 (
            .O(N__25434),
            .I(N__25431));
    Span4Mux_v I__3678 (
            .O(N__25431),
            .I(N__25428));
    Odrv4 I__3677 (
            .O(N__25428),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    CascadeMux I__3676 (
            .O(N__25425),
            .I(N__25422));
    InMux I__3675 (
            .O(N__25422),
            .I(N__25419));
    LocalMux I__3674 (
            .O(N__25419),
            .I(N__25416));
    Span4Mux_v I__3673 (
            .O(N__25416),
            .I(N__25413));
    Odrv4 I__3672 (
            .O(N__25413),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    CascadeMux I__3671 (
            .O(N__25410),
            .I(N__25407));
    InMux I__3670 (
            .O(N__25407),
            .I(N__25404));
    LocalMux I__3669 (
            .O(N__25404),
            .I(N__25401));
    Odrv4 I__3668 (
            .O(N__25401),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    CascadeMux I__3667 (
            .O(N__25398),
            .I(N__25395));
    InMux I__3666 (
            .O(N__25395),
            .I(N__25392));
    LocalMux I__3665 (
            .O(N__25392),
            .I(N__25389));
    Odrv4 I__3664 (
            .O(N__25389),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    InMux I__3663 (
            .O(N__25386),
            .I(N__25383));
    LocalMux I__3662 (
            .O(N__25383),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    InMux I__3661 (
            .O(N__25380),
            .I(N__25374));
    InMux I__3660 (
            .O(N__25379),
            .I(N__25374));
    LocalMux I__3659 (
            .O(N__25374),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ));
    InMux I__3658 (
            .O(N__25371),
            .I(N__25365));
    InMux I__3657 (
            .O(N__25370),
            .I(N__25365));
    LocalMux I__3656 (
            .O(N__25365),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ));
    InMux I__3655 (
            .O(N__25362),
            .I(N__25358));
    InMux I__3654 (
            .O(N__25361),
            .I(N__25354));
    LocalMux I__3653 (
            .O(N__25358),
            .I(N__25351));
    InMux I__3652 (
            .O(N__25357),
            .I(N__25347));
    LocalMux I__3651 (
            .O(N__25354),
            .I(N__25342));
    Span4Mux_v I__3650 (
            .O(N__25351),
            .I(N__25342));
    InMux I__3649 (
            .O(N__25350),
            .I(N__25339));
    LocalMux I__3648 (
            .O(N__25347),
            .I(N__25336));
    Span4Mux_v I__3647 (
            .O(N__25342),
            .I(N__25333));
    LocalMux I__3646 (
            .O(N__25339),
            .I(N__25330));
    Span4Mux_h I__3645 (
            .O(N__25336),
            .I(N__25327));
    Odrv4 I__3644 (
            .O(N__25333),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv12 I__3643 (
            .O(N__25330),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    Odrv4 I__3642 (
            .O(N__25327),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__3641 (
            .O(N__25320),
            .I(N__25317));
    LocalMux I__3640 (
            .O(N__25317),
            .I(N__25313));
    InMux I__3639 (
            .O(N__25316),
            .I(N__25309));
    Span4Mux_v I__3638 (
            .O(N__25313),
            .I(N__25306));
    InMux I__3637 (
            .O(N__25312),
            .I(N__25303));
    LocalMux I__3636 (
            .O(N__25309),
            .I(N__25296));
    Span4Mux_v I__3635 (
            .O(N__25306),
            .I(N__25296));
    LocalMux I__3634 (
            .O(N__25303),
            .I(N__25296));
    Odrv4 I__3633 (
            .O(N__25296),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__3632 (
            .O(N__25293),
            .I(N__25287));
    InMux I__3631 (
            .O(N__25292),
            .I(N__25287));
    LocalMux I__3630 (
            .O(N__25287),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ));
    CascadeMux I__3629 (
            .O(N__25284),
            .I(N__25280));
    InMux I__3628 (
            .O(N__25283),
            .I(N__25275));
    InMux I__3627 (
            .O(N__25280),
            .I(N__25275));
    LocalMux I__3626 (
            .O(N__25275),
            .I(N__25272));
    Odrv4 I__3625 (
            .O(N__25272),
            .I(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ));
    InMux I__3624 (
            .O(N__25269),
            .I(N__25266));
    LocalMux I__3623 (
            .O(N__25266),
            .I(N__25261));
    InMux I__3622 (
            .O(N__25265),
            .I(N__25258));
    InMux I__3621 (
            .O(N__25264),
            .I(N__25255));
    Span4Mux_v I__3620 (
            .O(N__25261),
            .I(N__25250));
    LocalMux I__3619 (
            .O(N__25258),
            .I(N__25250));
    LocalMux I__3618 (
            .O(N__25255),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    Odrv4 I__3617 (
            .O(N__25250),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    InMux I__3616 (
            .O(N__25245),
            .I(N__25241));
    InMux I__3615 (
            .O(N__25244),
            .I(N__25237));
    LocalMux I__3614 (
            .O(N__25241),
            .I(N__25234));
    InMux I__3613 (
            .O(N__25240),
            .I(N__25231));
    LocalMux I__3612 (
            .O(N__25237),
            .I(N__25227));
    Span4Mux_h I__3611 (
            .O(N__25234),
            .I(N__25224));
    LocalMux I__3610 (
            .O(N__25231),
            .I(N__25221));
    InMux I__3609 (
            .O(N__25230),
            .I(N__25218));
    Span4Mux_h I__3608 (
            .O(N__25227),
            .I(N__25213));
    Span4Mux_v I__3607 (
            .O(N__25224),
            .I(N__25213));
    Span4Mux_v I__3606 (
            .O(N__25221),
            .I(N__25208));
    LocalMux I__3605 (
            .O(N__25218),
            .I(N__25208));
    Odrv4 I__3604 (
            .O(N__25213),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    Odrv4 I__3603 (
            .O(N__25208),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__3602 (
            .O(N__25203),
            .I(N__25200));
    LocalMux I__3601 (
            .O(N__25200),
            .I(N__25196));
    InMux I__3600 (
            .O(N__25199),
            .I(N__25192));
    Span4Mux_v I__3599 (
            .O(N__25196),
            .I(N__25189));
    InMux I__3598 (
            .O(N__25195),
            .I(N__25186));
    LocalMux I__3597 (
            .O(N__25192),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    Odrv4 I__3596 (
            .O(N__25189),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    LocalMux I__3595 (
            .O(N__25186),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__3594 (
            .O(N__25179),
            .I(N__25175));
    InMux I__3593 (
            .O(N__25178),
            .I(N__25170));
    LocalMux I__3592 (
            .O(N__25175),
            .I(N__25167));
    InMux I__3591 (
            .O(N__25174),
            .I(N__25164));
    CascadeMux I__3590 (
            .O(N__25173),
            .I(N__25161));
    LocalMux I__3589 (
            .O(N__25170),
            .I(N__25156));
    Span4Mux_v I__3588 (
            .O(N__25167),
            .I(N__25156));
    LocalMux I__3587 (
            .O(N__25164),
            .I(N__25153));
    InMux I__3586 (
            .O(N__25161),
            .I(N__25150));
    Span4Mux_v I__3585 (
            .O(N__25156),
            .I(N__25147));
    Span4Mux_v I__3584 (
            .O(N__25153),
            .I(N__25144));
    LocalMux I__3583 (
            .O(N__25150),
            .I(N__25141));
    Odrv4 I__3582 (
            .O(N__25147),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__3581 (
            .O(N__25144),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    Odrv4 I__3580 (
            .O(N__25141),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__3579 (
            .O(N__25134),
            .I(N__25131));
    LocalMux I__3578 (
            .O(N__25131),
            .I(N__25126));
    InMux I__3577 (
            .O(N__25130),
            .I(N__25123));
    InMux I__3576 (
            .O(N__25129),
            .I(N__25120));
    Span4Mux_v I__3575 (
            .O(N__25126),
            .I(N__25114));
    LocalMux I__3574 (
            .O(N__25123),
            .I(N__25114));
    LocalMux I__3573 (
            .O(N__25120),
            .I(N__25111));
    InMux I__3572 (
            .O(N__25119),
            .I(N__25108));
    Span4Mux_v I__3571 (
            .O(N__25114),
            .I(N__25105));
    Span4Mux_h I__3570 (
            .O(N__25111),
            .I(N__25102));
    LocalMux I__3569 (
            .O(N__25108),
            .I(N__25099));
    Odrv4 I__3568 (
            .O(N__25105),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv4 I__3567 (
            .O(N__25102),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    Odrv12 I__3566 (
            .O(N__25099),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__3565 (
            .O(N__25092),
            .I(N__25088));
    InMux I__3564 (
            .O(N__25091),
            .I(N__25084));
    LocalMux I__3563 (
            .O(N__25088),
            .I(N__25081));
    InMux I__3562 (
            .O(N__25087),
            .I(N__25078));
    LocalMux I__3561 (
            .O(N__25084),
            .I(N__25073));
    Span4Mux_h I__3560 (
            .O(N__25081),
            .I(N__25073));
    LocalMux I__3559 (
            .O(N__25078),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv4 I__3558 (
            .O(N__25073),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__3557 (
            .O(N__25068),
            .I(N__25065));
    LocalMux I__3556 (
            .O(N__25065),
            .I(N__25060));
    InMux I__3555 (
            .O(N__25064),
            .I(N__25057));
    InMux I__3554 (
            .O(N__25063),
            .I(N__25054));
    Span12Mux_h I__3553 (
            .O(N__25060),
            .I(N__25051));
    LocalMux I__3552 (
            .O(N__25057),
            .I(N__25048));
    LocalMux I__3551 (
            .O(N__25054),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv12 I__3550 (
            .O(N__25051),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    Odrv4 I__3549 (
            .O(N__25048),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    InMux I__3548 (
            .O(N__25041),
            .I(N__25037));
    InMux I__3547 (
            .O(N__25040),
            .I(N__25034));
    LocalMux I__3546 (
            .O(N__25037),
            .I(N__25029));
    LocalMux I__3545 (
            .O(N__25034),
            .I(N__25026));
    InMux I__3544 (
            .O(N__25033),
            .I(N__25023));
    InMux I__3543 (
            .O(N__25032),
            .I(N__25020));
    Span4Mux_h I__3542 (
            .O(N__25029),
            .I(N__25017));
    Span4Mux_h I__3541 (
            .O(N__25026),
            .I(N__25012));
    LocalMux I__3540 (
            .O(N__25023),
            .I(N__25012));
    LocalMux I__3539 (
            .O(N__25020),
            .I(N__25009));
    Span4Mux_v I__3538 (
            .O(N__25017),
            .I(N__25006));
    Span4Mux_v I__3537 (
            .O(N__25012),
            .I(N__25001));
    Span4Mux_v I__3536 (
            .O(N__25009),
            .I(N__25001));
    Odrv4 I__3535 (
            .O(N__25006),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    Odrv4 I__3534 (
            .O(N__25001),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    InMux I__3533 (
            .O(N__24996),
            .I(N__24992));
    CascadeMux I__3532 (
            .O(N__24995),
            .I(N__24988));
    LocalMux I__3531 (
            .O(N__24992),
            .I(N__24985));
    InMux I__3530 (
            .O(N__24991),
            .I(N__24982));
    InMux I__3529 (
            .O(N__24988),
            .I(N__24979));
    Span4Mux_h I__3528 (
            .O(N__24985),
            .I(N__24974));
    LocalMux I__3527 (
            .O(N__24982),
            .I(N__24974));
    LocalMux I__3526 (
            .O(N__24979),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    Odrv4 I__3525 (
            .O(N__24974),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    InMux I__3524 (
            .O(N__24969),
            .I(N__24966));
    LocalMux I__3523 (
            .O(N__24966),
            .I(N__24960));
    InMux I__3522 (
            .O(N__24965),
            .I(N__24957));
    InMux I__3521 (
            .O(N__24964),
            .I(N__24954));
    InMux I__3520 (
            .O(N__24963),
            .I(N__24951));
    Span4Mux_v I__3519 (
            .O(N__24960),
            .I(N__24946));
    LocalMux I__3518 (
            .O(N__24957),
            .I(N__24946));
    LocalMux I__3517 (
            .O(N__24954),
            .I(N__24943));
    LocalMux I__3516 (
            .O(N__24951),
            .I(N__24940));
    Odrv4 I__3515 (
            .O(N__24946),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv4 I__3514 (
            .O(N__24943),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    Odrv4 I__3513 (
            .O(N__24940),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__3512 (
            .O(N__24933),
            .I(N__24929));
    InMux I__3511 (
            .O(N__24932),
            .I(N__24925));
    LocalMux I__3510 (
            .O(N__24929),
            .I(N__24922));
    InMux I__3509 (
            .O(N__24928),
            .I(N__24919));
    LocalMux I__3508 (
            .O(N__24925),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    Odrv12 I__3507 (
            .O(N__24922),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    LocalMux I__3506 (
            .O(N__24919),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    InMux I__3505 (
            .O(N__24912),
            .I(N__24907));
    InMux I__3504 (
            .O(N__24911),
            .I(N__24904));
    InMux I__3503 (
            .O(N__24910),
            .I(N__24901));
    LocalMux I__3502 (
            .O(N__24907),
            .I(N__24893));
    LocalMux I__3501 (
            .O(N__24904),
            .I(N__24893));
    LocalMux I__3500 (
            .O(N__24901),
            .I(N__24893));
    InMux I__3499 (
            .O(N__24900),
            .I(N__24890));
    Span4Mux_h I__3498 (
            .O(N__24893),
            .I(N__24885));
    LocalMux I__3497 (
            .O(N__24890),
            .I(N__24885));
    Odrv4 I__3496 (
            .O(N__24885),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__3495 (
            .O(N__24882),
            .I(N__24877));
    InMux I__3494 (
            .O(N__24881),
            .I(N__24874));
    InMux I__3493 (
            .O(N__24880),
            .I(N__24871));
    LocalMux I__3492 (
            .O(N__24877),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__3491 (
            .O(N__24874),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__3490 (
            .O(N__24871),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__3489 (
            .O(N__24864),
            .I(N__24859));
    InMux I__3488 (
            .O(N__24863),
            .I(N__24855));
    InMux I__3487 (
            .O(N__24862),
            .I(N__24852));
    LocalMux I__3486 (
            .O(N__24859),
            .I(N__24849));
    InMux I__3485 (
            .O(N__24858),
            .I(N__24846));
    LocalMux I__3484 (
            .O(N__24855),
            .I(N__24843));
    LocalMux I__3483 (
            .O(N__24852),
            .I(N__24840));
    Span4Mux_h I__3482 (
            .O(N__24849),
            .I(N__24835));
    LocalMux I__3481 (
            .O(N__24846),
            .I(N__24835));
    Span4Mux_h I__3480 (
            .O(N__24843),
            .I(N__24830));
    Span4Mux_h I__3479 (
            .O(N__24840),
            .I(N__24830));
    Odrv4 I__3478 (
            .O(N__24835),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    Odrv4 I__3477 (
            .O(N__24830),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__3476 (
            .O(N__24825),
            .I(N__24821));
    InMux I__3475 (
            .O(N__24824),
            .I(N__24817));
    LocalMux I__3474 (
            .O(N__24821),
            .I(N__24814));
    InMux I__3473 (
            .O(N__24820),
            .I(N__24811));
    LocalMux I__3472 (
            .O(N__24817),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    Odrv4 I__3471 (
            .O(N__24814),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    LocalMux I__3470 (
            .O(N__24811),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    InMux I__3469 (
            .O(N__24804),
            .I(N__24801));
    LocalMux I__3468 (
            .O(N__24801),
            .I(N__24796));
    InMux I__3467 (
            .O(N__24800),
            .I(N__24793));
    InMux I__3466 (
            .O(N__24799),
            .I(N__24790));
    Span4Mux_h I__3465 (
            .O(N__24796),
            .I(N__24786));
    LocalMux I__3464 (
            .O(N__24793),
            .I(N__24783));
    LocalMux I__3463 (
            .O(N__24790),
            .I(N__24780));
    InMux I__3462 (
            .O(N__24789),
            .I(N__24777));
    Span4Mux_v I__3461 (
            .O(N__24786),
            .I(N__24774));
    Span4Mux_h I__3460 (
            .O(N__24783),
            .I(N__24769));
    Span4Mux_v I__3459 (
            .O(N__24780),
            .I(N__24769));
    LocalMux I__3458 (
            .O(N__24777),
            .I(N__24766));
    Odrv4 I__3457 (
            .O(N__24774),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv4 I__3456 (
            .O(N__24769),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    Odrv12 I__3455 (
            .O(N__24766),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__3454 (
            .O(N__24759),
            .I(N__24755));
    InMux I__3453 (
            .O(N__24758),
            .I(N__24752));
    LocalMux I__3452 (
            .O(N__24755),
            .I(N__24748));
    LocalMux I__3451 (
            .O(N__24752),
            .I(N__24745));
    InMux I__3450 (
            .O(N__24751),
            .I(N__24742));
    Span4Mux_v I__3449 (
            .O(N__24748),
            .I(N__24737));
    Span4Mux_v I__3448 (
            .O(N__24745),
            .I(N__24737));
    LocalMux I__3447 (
            .O(N__24742),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    Odrv4 I__3446 (
            .O(N__24737),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__3445 (
            .O(N__24732),
            .I(N__24728));
    InMux I__3444 (
            .O(N__24731),
            .I(N__24725));
    LocalMux I__3443 (
            .O(N__24728),
            .I(N__24722));
    LocalMux I__3442 (
            .O(N__24725),
            .I(N__24716));
    Span4Mux_v I__3441 (
            .O(N__24722),
            .I(N__24716));
    InMux I__3440 (
            .O(N__24721),
            .I(N__24713));
    Span4Mux_v I__3439 (
            .O(N__24716),
            .I(N__24709));
    LocalMux I__3438 (
            .O(N__24713),
            .I(N__24706));
    InMux I__3437 (
            .O(N__24712),
            .I(N__24703));
    Odrv4 I__3436 (
            .O(N__24709),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    Odrv4 I__3435 (
            .O(N__24706),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__3434 (
            .O(N__24703),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    CascadeMux I__3433 (
            .O(N__24696),
            .I(N__24693));
    InMux I__3432 (
            .O(N__24693),
            .I(N__24689));
    InMux I__3431 (
            .O(N__24692),
            .I(N__24686));
    LocalMux I__3430 (
            .O(N__24689),
            .I(N__24681));
    LocalMux I__3429 (
            .O(N__24686),
            .I(N__24678));
    InMux I__3428 (
            .O(N__24685),
            .I(N__24675));
    InMux I__3427 (
            .O(N__24684),
            .I(N__24672));
    Span4Mux_h I__3426 (
            .O(N__24681),
            .I(N__24669));
    Span4Mux_h I__3425 (
            .O(N__24678),
            .I(N__24664));
    LocalMux I__3424 (
            .O(N__24675),
            .I(N__24664));
    LocalMux I__3423 (
            .O(N__24672),
            .I(N__24661));
    Odrv4 I__3422 (
            .O(N__24669),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__3421 (
            .O(N__24664),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    Odrv4 I__3420 (
            .O(N__24661),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__3419 (
            .O(N__24654),
            .I(N__24649));
    InMux I__3418 (
            .O(N__24653),
            .I(N__24646));
    InMux I__3417 (
            .O(N__24652),
            .I(N__24643));
    LocalMux I__3416 (
            .O(N__24649),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__3415 (
            .O(N__24646),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    LocalMux I__3414 (
            .O(N__24643),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    InMux I__3413 (
            .O(N__24636),
            .I(N__24631));
    InMux I__3412 (
            .O(N__24635),
            .I(N__24628));
    InMux I__3411 (
            .O(N__24634),
            .I(N__24625));
    LocalMux I__3410 (
            .O(N__24631),
            .I(N__24622));
    LocalMux I__3409 (
            .O(N__24628),
            .I(N__24617));
    LocalMux I__3408 (
            .O(N__24625),
            .I(N__24617));
    Odrv4 I__3407 (
            .O(N__24622),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__3406 (
            .O(N__24617),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__3405 (
            .O(N__24612),
            .I(N__24607));
    InMux I__3404 (
            .O(N__24611),
            .I(N__24604));
    InMux I__3403 (
            .O(N__24610),
            .I(N__24601));
    LocalMux I__3402 (
            .O(N__24607),
            .I(N__24597));
    LocalMux I__3401 (
            .O(N__24604),
            .I(N__24594));
    LocalMux I__3400 (
            .O(N__24601),
            .I(N__24591));
    InMux I__3399 (
            .O(N__24600),
            .I(N__24588));
    Span4Mux_v I__3398 (
            .O(N__24597),
            .I(N__24585));
    Span12Mux_h I__3397 (
            .O(N__24594),
            .I(N__24578));
    Span12Mux_s4_v I__3396 (
            .O(N__24591),
            .I(N__24578));
    LocalMux I__3395 (
            .O(N__24588),
            .I(N__24578));
    Odrv4 I__3394 (
            .O(N__24585),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv12 I__3393 (
            .O(N__24578),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__3392 (
            .O(N__24573),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__3391 (
            .O(N__24570),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    InMux I__3390 (
            .O(N__24567),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__3389 (
            .O(N__24564),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    InMux I__3388 (
            .O(N__24561),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__3387 (
            .O(N__24558),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__3386 (
            .O(N__24555),
            .I(N__24552));
    LocalMux I__3385 (
            .O(N__24552),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    CascadeMux I__3384 (
            .O(N__24549),
            .I(N__24546));
    InMux I__3383 (
            .O(N__24546),
            .I(N__24543));
    LocalMux I__3382 (
            .O(N__24543),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__3381 (
            .O(N__24540),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    InMux I__3380 (
            .O(N__24537),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__3379 (
            .O(N__24534),
            .I(N__24531));
    LocalMux I__3378 (
            .O(N__24531),
            .I(N__24528));
    Span4Mux_v I__3377 (
            .O(N__24528),
            .I(N__24525));
    Odrv4 I__3376 (
            .O(N__24525),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__3375 (
            .O(N__24522),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    CascadeMux I__3374 (
            .O(N__24519),
            .I(N__24516));
    InMux I__3373 (
            .O(N__24516),
            .I(N__24513));
    LocalMux I__3372 (
            .O(N__24513),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__3371 (
            .O(N__24510),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__3370 (
            .O(N__24507),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    CascadeMux I__3369 (
            .O(N__24504),
            .I(N__24501));
    InMux I__3368 (
            .O(N__24501),
            .I(N__24498));
    LocalMux I__3367 (
            .O(N__24498),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__3366 (
            .O(N__24495),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__3365 (
            .O(N__24492),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    InMux I__3364 (
            .O(N__24489),
            .I(bfn_8_20_0_));
    InMux I__3363 (
            .O(N__24486),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    InMux I__3362 (
            .O(N__24483),
            .I(N__24480));
    LocalMux I__3361 (
            .O(N__24480),
            .I(N__24477));
    Odrv4 I__3360 (
            .O(N__24477),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__3359 (
            .O(N__24474),
            .I(bfn_8_18_0_));
    InMux I__3358 (
            .O(N__24471),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    InMux I__3357 (
            .O(N__24468),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__3356 (
            .O(N__24465),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    InMux I__3355 (
            .O(N__24462),
            .I(N__24459));
    LocalMux I__3354 (
            .O(N__24459),
            .I(N__24456));
    Odrv12 I__3353 (
            .O(N__24456),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    InMux I__3352 (
            .O(N__24453),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__3351 (
            .O(N__24450),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    InMux I__3350 (
            .O(N__24447),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    CascadeMux I__3349 (
            .O(N__24444),
            .I(N__24441));
    InMux I__3348 (
            .O(N__24441),
            .I(N__24438));
    LocalMux I__3347 (
            .O(N__24438),
            .I(N__24435));
    Odrv12 I__3346 (
            .O(N__24435),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__3345 (
            .O(N__24432),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    InMux I__3344 (
            .O(N__24429),
            .I(bfn_8_19_0_));
    CascadeMux I__3343 (
            .O(N__24426),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__3342 (
            .O(N__24423),
            .I(N__24420));
    LocalMux I__3341 (
            .O(N__24420),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    InMux I__3340 (
            .O(N__24417),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    InMux I__3339 (
            .O(N__24414),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__3338 (
            .O(N__24411),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    CascadeMux I__3337 (
            .O(N__24408),
            .I(N__24405));
    InMux I__3336 (
            .O(N__24405),
            .I(N__24402));
    LocalMux I__3335 (
            .O(N__24402),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__3334 (
            .O(N__24399),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    CascadeMux I__3333 (
            .O(N__24396),
            .I(N__24393));
    InMux I__3332 (
            .O(N__24393),
            .I(N__24390));
    LocalMux I__3331 (
            .O(N__24390),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__3330 (
            .O(N__24387),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    InMux I__3329 (
            .O(N__24384),
            .I(N__24381));
    LocalMux I__3328 (
            .O(N__24381),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__3327 (
            .O(N__24378),
            .I(N__24375));
    LocalMux I__3326 (
            .O(N__24375),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__3325 (
            .O(N__24372),
            .I(N__24369));
    InMux I__3324 (
            .O(N__24369),
            .I(N__24364));
    InMux I__3323 (
            .O(N__24368),
            .I(N__24361));
    InMux I__3322 (
            .O(N__24367),
            .I(N__24358));
    LocalMux I__3321 (
            .O(N__24364),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3320 (
            .O(N__24361),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3319 (
            .O(N__24358),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__3318 (
            .O(N__24351),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    CascadeMux I__3317 (
            .O(N__24348),
            .I(N__24345));
    InMux I__3316 (
            .O(N__24345),
            .I(N__24340));
    InMux I__3315 (
            .O(N__24344),
            .I(N__24337));
    InMux I__3314 (
            .O(N__24343),
            .I(N__24334));
    LocalMux I__3313 (
            .O(N__24340),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3312 (
            .O(N__24337),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3311 (
            .O(N__24334),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__3310 (
            .O(N__24327),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    CascadeMux I__3309 (
            .O(N__24324),
            .I(N__24321));
    InMux I__3308 (
            .O(N__24321),
            .I(N__24316));
    InMux I__3307 (
            .O(N__24320),
            .I(N__24313));
    InMux I__3306 (
            .O(N__24319),
            .I(N__24310));
    LocalMux I__3305 (
            .O(N__24316),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3304 (
            .O(N__24313),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3303 (
            .O(N__24310),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__3302 (
            .O(N__24303),
            .I(bfn_8_12_0_));
    InMux I__3301 (
            .O(N__24300),
            .I(N__24295));
    InMux I__3300 (
            .O(N__24299),
            .I(N__24292));
    InMux I__3299 (
            .O(N__24298),
            .I(N__24289));
    LocalMux I__3298 (
            .O(N__24295),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3297 (
            .O(N__24292),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3296 (
            .O(N__24289),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__3295 (
            .O(N__24282),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    CascadeMux I__3294 (
            .O(N__24279),
            .I(N__24276));
    InMux I__3293 (
            .O(N__24276),
            .I(N__24271));
    InMux I__3292 (
            .O(N__24275),
            .I(N__24268));
    InMux I__3291 (
            .O(N__24274),
            .I(N__24265));
    LocalMux I__3290 (
            .O(N__24271),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3289 (
            .O(N__24268),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3288 (
            .O(N__24265),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__3287 (
            .O(N__24258),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    CascadeMux I__3286 (
            .O(N__24255),
            .I(N__24250));
    CascadeMux I__3285 (
            .O(N__24254),
            .I(N__24247));
    InMux I__3284 (
            .O(N__24253),
            .I(N__24244));
    InMux I__3283 (
            .O(N__24250),
            .I(N__24239));
    InMux I__3282 (
            .O(N__24247),
            .I(N__24239));
    LocalMux I__3281 (
            .O(N__24244),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__3280 (
            .O(N__24239),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__3279 (
            .O(N__24234),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__3278 (
            .O(N__24231),
            .I(N__24227));
    InMux I__3277 (
            .O(N__24230),
            .I(N__24224));
    LocalMux I__3276 (
            .O(N__24227),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__3275 (
            .O(N__24224),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    InMux I__3274 (
            .O(N__24219),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__3273 (
            .O(N__24216),
            .I(N__24194));
    InMux I__3272 (
            .O(N__24215),
            .I(N__24194));
    InMux I__3271 (
            .O(N__24214),
            .I(N__24194));
    InMux I__3270 (
            .O(N__24213),
            .I(N__24194));
    InMux I__3269 (
            .O(N__24212),
            .I(N__24185));
    InMux I__3268 (
            .O(N__24211),
            .I(N__24185));
    InMux I__3267 (
            .O(N__24210),
            .I(N__24185));
    InMux I__3266 (
            .O(N__24209),
            .I(N__24185));
    InMux I__3265 (
            .O(N__24208),
            .I(N__24180));
    InMux I__3264 (
            .O(N__24207),
            .I(N__24180));
    InMux I__3263 (
            .O(N__24206),
            .I(N__24155));
    InMux I__3262 (
            .O(N__24205),
            .I(N__24155));
    InMux I__3261 (
            .O(N__24204),
            .I(N__24155));
    InMux I__3260 (
            .O(N__24203),
            .I(N__24155));
    LocalMux I__3259 (
            .O(N__24194),
            .I(N__24152));
    LocalMux I__3258 (
            .O(N__24185),
            .I(N__24149));
    LocalMux I__3257 (
            .O(N__24180),
            .I(N__24146));
    InMux I__3256 (
            .O(N__24179),
            .I(N__24137));
    InMux I__3255 (
            .O(N__24178),
            .I(N__24137));
    InMux I__3254 (
            .O(N__24177),
            .I(N__24137));
    InMux I__3253 (
            .O(N__24176),
            .I(N__24137));
    InMux I__3252 (
            .O(N__24175),
            .I(N__24128));
    InMux I__3251 (
            .O(N__24174),
            .I(N__24128));
    InMux I__3250 (
            .O(N__24173),
            .I(N__24128));
    InMux I__3249 (
            .O(N__24172),
            .I(N__24128));
    InMux I__3248 (
            .O(N__24171),
            .I(N__24119));
    InMux I__3247 (
            .O(N__24170),
            .I(N__24119));
    InMux I__3246 (
            .O(N__24169),
            .I(N__24119));
    InMux I__3245 (
            .O(N__24168),
            .I(N__24119));
    InMux I__3244 (
            .O(N__24167),
            .I(N__24110));
    InMux I__3243 (
            .O(N__24166),
            .I(N__24110));
    InMux I__3242 (
            .O(N__24165),
            .I(N__24110));
    InMux I__3241 (
            .O(N__24164),
            .I(N__24110));
    LocalMux I__3240 (
            .O(N__24155),
            .I(N__24107));
    Span4Mux_v I__3239 (
            .O(N__24152),
            .I(N__24096));
    Span4Mux_v I__3238 (
            .O(N__24149),
            .I(N__24096));
    Span4Mux_v I__3237 (
            .O(N__24146),
            .I(N__24096));
    LocalMux I__3236 (
            .O(N__24137),
            .I(N__24096));
    LocalMux I__3235 (
            .O(N__24128),
            .I(N__24096));
    LocalMux I__3234 (
            .O(N__24119),
            .I(N__24091));
    LocalMux I__3233 (
            .O(N__24110),
            .I(N__24091));
    Span4Mux_h I__3232 (
            .O(N__24107),
            .I(N__24088));
    Span4Mux_h I__3231 (
            .O(N__24096),
            .I(N__24085));
    Odrv4 I__3230 (
            .O(N__24091),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__3229 (
            .O(N__24088),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__3228 (
            .O(N__24085),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__3227 (
            .O(N__24078),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__3226 (
            .O(N__24075),
            .I(N__24071));
    InMux I__3225 (
            .O(N__24074),
            .I(N__24068));
    LocalMux I__3224 (
            .O(N__24071),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__3223 (
            .O(N__24068),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CEMux I__3222 (
            .O(N__24063),
            .I(N__24057));
    CEMux I__3221 (
            .O(N__24062),
            .I(N__24054));
    CEMux I__3220 (
            .O(N__24061),
            .I(N__24051));
    CEMux I__3219 (
            .O(N__24060),
            .I(N__24048));
    LocalMux I__3218 (
            .O(N__24057),
            .I(N__24045));
    LocalMux I__3217 (
            .O(N__24054),
            .I(N__24042));
    LocalMux I__3216 (
            .O(N__24051),
            .I(N__24039));
    LocalMux I__3215 (
            .O(N__24048),
            .I(N__24036));
    Span4Mux_h I__3214 (
            .O(N__24045),
            .I(N__24033));
    Span4Mux_v I__3213 (
            .O(N__24042),
            .I(N__24026));
    Span4Mux_v I__3212 (
            .O(N__24039),
            .I(N__24026));
    Span4Mux_h I__3211 (
            .O(N__24036),
            .I(N__24026));
    Odrv4 I__3210 (
            .O(N__24033),
            .I(\delay_measurement_inst.delay_tr_timer.N_344_i ));
    Odrv4 I__3209 (
            .O(N__24026),
            .I(\delay_measurement_inst.delay_tr_timer.N_344_i ));
    CascadeMux I__3208 (
            .O(N__24021),
            .I(N__24018));
    InMux I__3207 (
            .O(N__24018),
            .I(N__24013));
    InMux I__3206 (
            .O(N__24017),
            .I(N__24010));
    InMux I__3205 (
            .O(N__24016),
            .I(N__24007));
    LocalMux I__3204 (
            .O(N__24013),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__3203 (
            .O(N__24010),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__3202 (
            .O(N__24007),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__3201 (
            .O(N__24000),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    CascadeMux I__3200 (
            .O(N__23997),
            .I(N__23994));
    InMux I__3199 (
            .O(N__23994),
            .I(N__23989));
    InMux I__3198 (
            .O(N__23993),
            .I(N__23986));
    InMux I__3197 (
            .O(N__23992),
            .I(N__23983));
    LocalMux I__3196 (
            .O(N__23989),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__3195 (
            .O(N__23986),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__3194 (
            .O(N__23983),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__3193 (
            .O(N__23976),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    CascadeMux I__3192 (
            .O(N__23973),
            .I(N__23970));
    InMux I__3191 (
            .O(N__23970),
            .I(N__23965));
    InMux I__3190 (
            .O(N__23969),
            .I(N__23962));
    InMux I__3189 (
            .O(N__23968),
            .I(N__23959));
    LocalMux I__3188 (
            .O(N__23965),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__3187 (
            .O(N__23962),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__3186 (
            .O(N__23959),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__3185 (
            .O(N__23952),
            .I(bfn_8_11_0_));
    CascadeMux I__3184 (
            .O(N__23949),
            .I(N__23946));
    InMux I__3183 (
            .O(N__23946),
            .I(N__23941));
    InMux I__3182 (
            .O(N__23945),
            .I(N__23938));
    InMux I__3181 (
            .O(N__23944),
            .I(N__23935));
    LocalMux I__3180 (
            .O(N__23941),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__3179 (
            .O(N__23938),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__3178 (
            .O(N__23935),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__3177 (
            .O(N__23928),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    CascadeMux I__3176 (
            .O(N__23925),
            .I(N__23922));
    InMux I__3175 (
            .O(N__23922),
            .I(N__23917));
    InMux I__3174 (
            .O(N__23921),
            .I(N__23914));
    InMux I__3173 (
            .O(N__23920),
            .I(N__23911));
    LocalMux I__3172 (
            .O(N__23917),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__3171 (
            .O(N__23914),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__3170 (
            .O(N__23911),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__3169 (
            .O(N__23904),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    CascadeMux I__3168 (
            .O(N__23901),
            .I(N__23898));
    InMux I__3167 (
            .O(N__23898),
            .I(N__23893));
    InMux I__3166 (
            .O(N__23897),
            .I(N__23890));
    InMux I__3165 (
            .O(N__23896),
            .I(N__23887));
    LocalMux I__3164 (
            .O(N__23893),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__3163 (
            .O(N__23890),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__3162 (
            .O(N__23887),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__3161 (
            .O(N__23880),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    CascadeMux I__3160 (
            .O(N__23877),
            .I(N__23874));
    InMux I__3159 (
            .O(N__23874),
            .I(N__23869));
    InMux I__3158 (
            .O(N__23873),
            .I(N__23866));
    InMux I__3157 (
            .O(N__23872),
            .I(N__23863));
    LocalMux I__3156 (
            .O(N__23869),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3155 (
            .O(N__23866),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3154 (
            .O(N__23863),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__3153 (
            .O(N__23856),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    CascadeMux I__3152 (
            .O(N__23853),
            .I(N__23850));
    InMux I__3151 (
            .O(N__23850),
            .I(N__23845));
    InMux I__3150 (
            .O(N__23849),
            .I(N__23842));
    InMux I__3149 (
            .O(N__23848),
            .I(N__23839));
    LocalMux I__3148 (
            .O(N__23845),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3147 (
            .O(N__23842),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3146 (
            .O(N__23839),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__3145 (
            .O(N__23832),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    CascadeMux I__3144 (
            .O(N__23829),
            .I(N__23826));
    InMux I__3143 (
            .O(N__23826),
            .I(N__23821));
    InMux I__3142 (
            .O(N__23825),
            .I(N__23818));
    InMux I__3141 (
            .O(N__23824),
            .I(N__23815));
    LocalMux I__3140 (
            .O(N__23821),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__3139 (
            .O(N__23818),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__3138 (
            .O(N__23815),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__3137 (
            .O(N__23808),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    CascadeMux I__3136 (
            .O(N__23805),
            .I(N__23802));
    InMux I__3135 (
            .O(N__23802),
            .I(N__23797));
    InMux I__3134 (
            .O(N__23801),
            .I(N__23794));
    InMux I__3133 (
            .O(N__23800),
            .I(N__23791));
    LocalMux I__3132 (
            .O(N__23797),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__3131 (
            .O(N__23794),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__3130 (
            .O(N__23791),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__3129 (
            .O(N__23784),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    CascadeMux I__3128 (
            .O(N__23781),
            .I(N__23778));
    InMux I__3127 (
            .O(N__23778),
            .I(N__23773));
    InMux I__3126 (
            .O(N__23777),
            .I(N__23770));
    InMux I__3125 (
            .O(N__23776),
            .I(N__23767));
    LocalMux I__3124 (
            .O(N__23773),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__3123 (
            .O(N__23770),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__3122 (
            .O(N__23767),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__3121 (
            .O(N__23760),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    CascadeMux I__3120 (
            .O(N__23757),
            .I(N__23754));
    InMux I__3119 (
            .O(N__23754),
            .I(N__23749));
    InMux I__3118 (
            .O(N__23753),
            .I(N__23746));
    InMux I__3117 (
            .O(N__23752),
            .I(N__23743));
    LocalMux I__3116 (
            .O(N__23749),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__3115 (
            .O(N__23746),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__3114 (
            .O(N__23743),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__3113 (
            .O(N__23736),
            .I(bfn_8_10_0_));
    CascadeMux I__3112 (
            .O(N__23733),
            .I(N__23730));
    InMux I__3111 (
            .O(N__23730),
            .I(N__23725));
    InMux I__3110 (
            .O(N__23729),
            .I(N__23722));
    InMux I__3109 (
            .O(N__23728),
            .I(N__23719));
    LocalMux I__3108 (
            .O(N__23725),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__3107 (
            .O(N__23722),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__3106 (
            .O(N__23719),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__3105 (
            .O(N__23712),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    CascadeMux I__3104 (
            .O(N__23709),
            .I(N__23706));
    InMux I__3103 (
            .O(N__23706),
            .I(N__23701));
    InMux I__3102 (
            .O(N__23705),
            .I(N__23698));
    InMux I__3101 (
            .O(N__23704),
            .I(N__23695));
    LocalMux I__3100 (
            .O(N__23701),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__3099 (
            .O(N__23698),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__3098 (
            .O(N__23695),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__3097 (
            .O(N__23688),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    CascadeMux I__3096 (
            .O(N__23685),
            .I(N__23682));
    InMux I__3095 (
            .O(N__23682),
            .I(N__23677));
    InMux I__3094 (
            .O(N__23681),
            .I(N__23674));
    InMux I__3093 (
            .O(N__23680),
            .I(N__23671));
    LocalMux I__3092 (
            .O(N__23677),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__3091 (
            .O(N__23674),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__3090 (
            .O(N__23671),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__3089 (
            .O(N__23664),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    CascadeMux I__3088 (
            .O(N__23661),
            .I(N__23658));
    InMux I__3087 (
            .O(N__23658),
            .I(N__23653));
    InMux I__3086 (
            .O(N__23657),
            .I(N__23650));
    InMux I__3085 (
            .O(N__23656),
            .I(N__23647));
    LocalMux I__3084 (
            .O(N__23653),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3083 (
            .O(N__23650),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3082 (
            .O(N__23647),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__3081 (
            .O(N__23640),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    CascadeMux I__3080 (
            .O(N__23637),
            .I(N__23634));
    InMux I__3079 (
            .O(N__23634),
            .I(N__23629));
    InMux I__3078 (
            .O(N__23633),
            .I(N__23626));
    InMux I__3077 (
            .O(N__23632),
            .I(N__23623));
    LocalMux I__3076 (
            .O(N__23629),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3075 (
            .O(N__23626),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3074 (
            .O(N__23623),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__3073 (
            .O(N__23616),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__3072 (
            .O(N__23613),
            .I(N__23610));
    LocalMux I__3071 (
            .O(N__23610),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__3070 (
            .O(N__23607),
            .I(N__23604));
    LocalMux I__3069 (
            .O(N__23604),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ));
    InMux I__3068 (
            .O(N__23601),
            .I(N__23597));
    CascadeMux I__3067 (
            .O(N__23600),
            .I(N__23594));
    LocalMux I__3066 (
            .O(N__23597),
            .I(N__23590));
    InMux I__3065 (
            .O(N__23594),
            .I(N__23587));
    InMux I__3064 (
            .O(N__23593),
            .I(N__23584));
    Odrv12 I__3063 (
            .O(N__23590),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__3062 (
            .O(N__23587),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__3061 (
            .O(N__23584),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    InMux I__3060 (
            .O(N__23577),
            .I(bfn_8_9_0_));
    InMux I__3059 (
            .O(N__23574),
            .I(N__23569));
    InMux I__3058 (
            .O(N__23573),
            .I(N__23566));
    InMux I__3057 (
            .O(N__23572),
            .I(N__23563));
    LocalMux I__3056 (
            .O(N__23569),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3055 (
            .O(N__23566),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__3054 (
            .O(N__23563),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__3053 (
            .O(N__23556),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    CascadeMux I__3052 (
            .O(N__23553),
            .I(N__23550));
    InMux I__3051 (
            .O(N__23550),
            .I(N__23545));
    InMux I__3050 (
            .O(N__23549),
            .I(N__23542));
    InMux I__3049 (
            .O(N__23548),
            .I(N__23539));
    LocalMux I__3048 (
            .O(N__23545),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__3047 (
            .O(N__23542),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__3046 (
            .O(N__23539),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__3045 (
            .O(N__23532),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    CascadeMux I__3044 (
            .O(N__23529),
            .I(N__23524));
    CascadeMux I__3043 (
            .O(N__23528),
            .I(N__23521));
    InMux I__3042 (
            .O(N__23527),
            .I(N__23518));
    InMux I__3041 (
            .O(N__23524),
            .I(N__23513));
    InMux I__3040 (
            .O(N__23521),
            .I(N__23513));
    LocalMux I__3039 (
            .O(N__23518),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__3038 (
            .O(N__23513),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__3037 (
            .O(N__23508),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    CascadeMux I__3036 (
            .O(N__23505),
            .I(N__23502));
    InMux I__3035 (
            .O(N__23502),
            .I(N__23497));
    InMux I__3034 (
            .O(N__23501),
            .I(N__23494));
    InMux I__3033 (
            .O(N__23500),
            .I(N__23491));
    LocalMux I__3032 (
            .O(N__23497),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__3031 (
            .O(N__23494),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__3030 (
            .O(N__23491),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__3029 (
            .O(N__23484),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    CascadeMux I__3028 (
            .O(N__23481),
            .I(N__23478));
    InMux I__3027 (
            .O(N__23478),
            .I(N__23475));
    LocalMux I__3026 (
            .O(N__23475),
            .I(N__23472));
    Span4Mux_h I__3025 (
            .O(N__23472),
            .I(N__23469));
    Odrv4 I__3024 (
            .O(N__23469),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    InMux I__3023 (
            .O(N__23466),
            .I(N__23463));
    LocalMux I__3022 (
            .O(N__23463),
            .I(N__23460));
    Odrv12 I__3021 (
            .O(N__23460),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__3020 (
            .O(N__23457),
            .I(N__23454));
    LocalMux I__3019 (
            .O(N__23454),
            .I(N__23451));
    Span4Mux_h I__3018 (
            .O(N__23451),
            .I(N__23448));
    Odrv4 I__3017 (
            .O(N__23448),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    InMux I__3016 (
            .O(N__23445),
            .I(N__23442));
    LocalMux I__3015 (
            .O(N__23442),
            .I(N__23439));
    Span12Mux_v I__3014 (
            .O(N__23439),
            .I(N__23436));
    Odrv12 I__3013 (
            .O(N__23436),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    InMux I__3012 (
            .O(N__23433),
            .I(N__23430));
    LocalMux I__3011 (
            .O(N__23430),
            .I(N__23427));
    Span4Mux_h I__3010 (
            .O(N__23427),
            .I(N__23424));
    Odrv4 I__3009 (
            .O(N__23424),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    InMux I__3008 (
            .O(N__23421),
            .I(N__23418));
    LocalMux I__3007 (
            .O(N__23418),
            .I(N__23415));
    Odrv12 I__3006 (
            .O(N__23415),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    InMux I__3005 (
            .O(N__23412),
            .I(N__23409));
    LocalMux I__3004 (
            .O(N__23409),
            .I(N__23406));
    Span4Mux_h I__3003 (
            .O(N__23406),
            .I(N__23403));
    Odrv4 I__3002 (
            .O(N__23403),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    CascadeMux I__3001 (
            .O(N__23400),
            .I(N__23397));
    InMux I__3000 (
            .O(N__23397),
            .I(N__23394));
    LocalMux I__2999 (
            .O(N__23394),
            .I(N__23391));
    Span12Mux_s7_h I__2998 (
            .O(N__23391),
            .I(N__23388));
    Odrv12 I__2997 (
            .O(N__23388),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__2996 (
            .O(N__23385),
            .I(N__23382));
    InMux I__2995 (
            .O(N__23382),
            .I(N__23379));
    LocalMux I__2994 (
            .O(N__23379),
            .I(N__23376));
    Odrv12 I__2993 (
            .O(N__23376),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__2992 (
            .O(N__23373),
            .I(N__23370));
    LocalMux I__2991 (
            .O(N__23370),
            .I(N__23367));
    Span4Mux_h I__2990 (
            .O(N__23367),
            .I(N__23364));
    Odrv4 I__2989 (
            .O(N__23364),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    InMux I__2988 (
            .O(N__23361),
            .I(N__23358));
    LocalMux I__2987 (
            .O(N__23358),
            .I(N__23355));
    Odrv4 I__2986 (
            .O(N__23355),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__2985 (
            .O(N__23352),
            .I(N__23349));
    LocalMux I__2984 (
            .O(N__23349),
            .I(N__23346));
    Span4Mux_h I__2983 (
            .O(N__23346),
            .I(N__23343));
    Odrv4 I__2982 (
            .O(N__23343),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    InMux I__2981 (
            .O(N__23340),
            .I(N__23337));
    LocalMux I__2980 (
            .O(N__23337),
            .I(N__23334));
    Odrv4 I__2979 (
            .O(N__23334),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    CascadeMux I__2978 (
            .O(N__23331),
            .I(N__23328));
    InMux I__2977 (
            .O(N__23328),
            .I(N__23325));
    LocalMux I__2976 (
            .O(N__23325),
            .I(N__23322));
    Span4Mux_h I__2975 (
            .O(N__23322),
            .I(N__23319));
    Odrv4 I__2974 (
            .O(N__23319),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    InMux I__2973 (
            .O(N__23316),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__2972 (
            .O(N__23313),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__2971 (
            .O(N__23310),
            .I(bfn_7_13_0_));
    InMux I__2970 (
            .O(N__23307),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__2969 (
            .O(N__23304),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__2968 (
            .O(N__23301),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__2967 (
            .O(N__23298),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__2966 (
            .O(N__23295),
            .I(N__23290));
    CEMux I__2965 (
            .O(N__23294),
            .I(N__23287));
    CEMux I__2964 (
            .O(N__23293),
            .I(N__23284));
    LocalMux I__2963 (
            .O(N__23290),
            .I(N__23276));
    LocalMux I__2962 (
            .O(N__23287),
            .I(N__23276));
    LocalMux I__2961 (
            .O(N__23284),
            .I(N__23273));
    CEMux I__2960 (
            .O(N__23283),
            .I(N__23270));
    CEMux I__2959 (
            .O(N__23282),
            .I(N__23267));
    CEMux I__2958 (
            .O(N__23281),
            .I(N__23264));
    Span4Mux_v I__2957 (
            .O(N__23276),
            .I(N__23261));
    Span4Mux_v I__2956 (
            .O(N__23273),
            .I(N__23256));
    LocalMux I__2955 (
            .O(N__23270),
            .I(N__23256));
    LocalMux I__2954 (
            .O(N__23267),
            .I(N__23251));
    LocalMux I__2953 (
            .O(N__23264),
            .I(N__23251));
    Span4Mux_h I__2952 (
            .O(N__23261),
            .I(N__23246));
    Span4Mux_h I__2951 (
            .O(N__23256),
            .I(N__23246));
    Span4Mux_h I__2950 (
            .O(N__23251),
            .I(N__23243));
    Odrv4 I__2949 (
            .O(N__23246),
            .I(\delay_measurement_inst.delay_tr_timer.N_343_i ));
    Odrv4 I__2948 (
            .O(N__23243),
            .I(\delay_measurement_inst.delay_tr_timer.N_343_i ));
    InMux I__2947 (
            .O(N__23238),
            .I(N__23235));
    LocalMux I__2946 (
            .O(N__23235),
            .I(N__23232));
    Span4Mux_h I__2945 (
            .O(N__23232),
            .I(N__23229));
    Odrv4 I__2944 (
            .O(N__23229),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__2943 (
            .O(N__23226),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__2942 (
            .O(N__23223),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__2941 (
            .O(N__23220),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__2940 (
            .O(N__23217),
            .I(bfn_7_12_0_));
    InMux I__2939 (
            .O(N__23214),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__2938 (
            .O(N__23211),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__2937 (
            .O(N__23208),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__2936 (
            .O(N__23205),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__2935 (
            .O(N__23202),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__2934 (
            .O(N__23199),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__2933 (
            .O(N__23196),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    InMux I__2932 (
            .O(N__23193),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__2931 (
            .O(N__23190),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__2930 (
            .O(N__23187),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__2929 (
            .O(N__23184),
            .I(bfn_7_11_0_));
    InMux I__2928 (
            .O(N__23181),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__2927 (
            .O(N__23178),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__2926 (
            .O(N__23175),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__2925 (
            .O(N__23172),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__2924 (
            .O(N__23169),
            .I(N__23166));
    LocalMux I__2923 (
            .O(N__23166),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    CascadeMux I__2922 (
            .O(N__23163),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ));
    CascadeMux I__2921 (
            .O(N__23160),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    CascadeMux I__2920 (
            .O(N__23157),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ));
    InMux I__2919 (
            .O(N__23154),
            .I(N__23151));
    LocalMux I__2918 (
            .O(N__23151),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    InMux I__2917 (
            .O(N__23148),
            .I(N__23145));
    LocalMux I__2916 (
            .O(N__23145),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ));
    InMux I__2915 (
            .O(N__23142),
            .I(N__23139));
    LocalMux I__2914 (
            .O(N__23139),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ));
    InMux I__2913 (
            .O(N__23136),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__2912 (
            .O(N__23133),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__2911 (
            .O(N__23130),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ));
    InMux I__2910 (
            .O(N__23127),
            .I(N__23124));
    LocalMux I__2909 (
            .O(N__23124),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__2908 (
            .O(N__23121),
            .I(N__23118));
    LocalMux I__2907 (
            .O(N__23118),
            .I(N__23115));
    Odrv4 I__2906 (
            .O(N__23115),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    InMux I__2905 (
            .O(N__23112),
            .I(N__23109));
    LocalMux I__2904 (
            .O(N__23109),
            .I(N__23106));
    Odrv4 I__2903 (
            .O(N__23106),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__2902 (
            .O(N__23103),
            .I(N__23100));
    LocalMux I__2901 (
            .O(N__23100),
            .I(N__23097));
    Odrv4 I__2900 (
            .O(N__23097),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    InMux I__2899 (
            .O(N__23094),
            .I(N__23091));
    LocalMux I__2898 (
            .O(N__23091),
            .I(N__23087));
    InMux I__2897 (
            .O(N__23090),
            .I(N__23084));
    Span4Mux_v I__2896 (
            .O(N__23087),
            .I(N__23081));
    LocalMux I__2895 (
            .O(N__23084),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv4 I__2894 (
            .O(N__23081),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    InMux I__2893 (
            .O(N__23076),
            .I(N__23073));
    LocalMux I__2892 (
            .O(N__23073),
            .I(N__23069));
    InMux I__2891 (
            .O(N__23072),
            .I(N__23066));
    Odrv4 I__2890 (
            .O(N__23069),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    LocalMux I__2889 (
            .O(N__23066),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__2888 (
            .O(N__23061),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__2887 (
            .O(N__23058),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    InMux I__2886 (
            .O(N__23055),
            .I(N__23050));
    CascadeMux I__2885 (
            .O(N__23054),
            .I(N__23047));
    InMux I__2884 (
            .O(N__23053),
            .I(N__23044));
    LocalMux I__2883 (
            .O(N__23050),
            .I(N__23041));
    InMux I__2882 (
            .O(N__23047),
            .I(N__23038));
    LocalMux I__2881 (
            .O(N__23044),
            .I(N__23028));
    Span4Mux_h I__2880 (
            .O(N__23041),
            .I(N__23023));
    LocalMux I__2879 (
            .O(N__23038),
            .I(N__23023));
    InMux I__2878 (
            .O(N__23037),
            .I(N__23020));
    InMux I__2877 (
            .O(N__23036),
            .I(N__23011));
    InMux I__2876 (
            .O(N__23035),
            .I(N__23011));
    InMux I__2875 (
            .O(N__23034),
            .I(N__23011));
    InMux I__2874 (
            .O(N__23033),
            .I(N__23011));
    InMux I__2873 (
            .O(N__23032),
            .I(N__23006));
    InMux I__2872 (
            .O(N__23031),
            .I(N__23006));
    Span4Mux_v I__2871 (
            .O(N__23028),
            .I(N__22999));
    Span4Mux_v I__2870 (
            .O(N__23023),
            .I(N__22999));
    LocalMux I__2869 (
            .O(N__23020),
            .I(N__22999));
    LocalMux I__2868 (
            .O(N__23011),
            .I(N__22996));
    LocalMux I__2867 (
            .O(N__23006),
            .I(N__22993));
    Span4Mux_h I__2866 (
            .O(N__22999),
            .I(N__22990));
    Span12Mux_s3_h I__2865 (
            .O(N__22996),
            .I(N__22985));
    Sp12to4 I__2864 (
            .O(N__22993),
            .I(N__22985));
    Span4Mux_v I__2863 (
            .O(N__22990),
            .I(N__22982));
    Span12Mux_v I__2862 (
            .O(N__22985),
            .I(N__22979));
    Span4Mux_v I__2861 (
            .O(N__22982),
            .I(N__22976));
    Odrv12 I__2860 (
            .O(N__22979),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    Odrv4 I__2859 (
            .O(N__22976),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__2858 (
            .O(N__22971),
            .I(N__22968));
    LocalMux I__2857 (
            .O(N__22968),
            .I(N__22965));
    Odrv4 I__2856 (
            .O(N__22965),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__2855 (
            .O(N__22962),
            .I(N__22959));
    LocalMux I__2854 (
            .O(N__22959),
            .I(N__22956));
    Odrv4 I__2853 (
            .O(N__22956),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    InMux I__2852 (
            .O(N__22953),
            .I(N__22950));
    LocalMux I__2851 (
            .O(N__22950),
            .I(N__22947));
    Odrv4 I__2850 (
            .O(N__22947),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    InMux I__2849 (
            .O(N__22944),
            .I(N__22941));
    LocalMux I__2848 (
            .O(N__22941),
            .I(N__22938));
    Odrv12 I__2847 (
            .O(N__22938),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    InMux I__2846 (
            .O(N__22935),
            .I(N__22932));
    LocalMux I__2845 (
            .O(N__22932),
            .I(N__22929));
    Odrv4 I__2844 (
            .O(N__22929),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__2843 (
            .O(N__22926),
            .I(N__22923));
    LocalMux I__2842 (
            .O(N__22923),
            .I(N__22920));
    Odrv4 I__2841 (
            .O(N__22920),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__2840 (
            .O(N__22917),
            .I(N__22914));
    LocalMux I__2839 (
            .O(N__22914),
            .I(N__22911));
    Odrv4 I__2838 (
            .O(N__22911),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__2837 (
            .O(N__22908),
            .I(N__22904));
    InMux I__2836 (
            .O(N__22907),
            .I(N__22901));
    LocalMux I__2835 (
            .O(N__22904),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    LocalMux I__2834 (
            .O(N__22901),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__2833 (
            .O(N__22896),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    InMux I__2832 (
            .O(N__22893),
            .I(N__22889));
    InMux I__2831 (
            .O(N__22892),
            .I(N__22886));
    LocalMux I__2830 (
            .O(N__22889),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    LocalMux I__2829 (
            .O(N__22886),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__2828 (
            .O(N__22881),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    InMux I__2827 (
            .O(N__22878),
            .I(N__22875));
    LocalMux I__2826 (
            .O(N__22875),
            .I(N__22872));
    Odrv4 I__2825 (
            .O(N__22872),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__2824 (
            .O(N__22869),
            .I(N__22865));
    InMux I__2823 (
            .O(N__22868),
            .I(N__22862));
    LocalMux I__2822 (
            .O(N__22865),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    LocalMux I__2821 (
            .O(N__22862),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__2820 (
            .O(N__22857),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    InMux I__2819 (
            .O(N__22854),
            .I(N__22848));
    InMux I__2818 (
            .O(N__22853),
            .I(N__22848));
    LocalMux I__2817 (
            .O(N__22848),
            .I(N__22845));
    Odrv4 I__2816 (
            .O(N__22845),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    InMux I__2815 (
            .O(N__22842),
            .I(bfn_5_18_0_));
    InMux I__2814 (
            .O(N__22839),
            .I(N__22833));
    InMux I__2813 (
            .O(N__22838),
            .I(N__22833));
    LocalMux I__2812 (
            .O(N__22833),
            .I(N__22830));
    Odrv4 I__2811 (
            .O(N__22830),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    InMux I__2810 (
            .O(N__22827),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    InMux I__2809 (
            .O(N__22824),
            .I(N__22821));
    LocalMux I__2808 (
            .O(N__22821),
            .I(N__22818));
    Odrv12 I__2807 (
            .O(N__22818),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    InMux I__2806 (
            .O(N__22815),
            .I(N__22812));
    LocalMux I__2805 (
            .O(N__22812),
            .I(N__22808));
    InMux I__2804 (
            .O(N__22811),
            .I(N__22805));
    Span4Mux_h I__2803 (
            .O(N__22808),
            .I(N__22802));
    LocalMux I__2802 (
            .O(N__22805),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    Odrv4 I__2801 (
            .O(N__22802),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__2800 (
            .O(N__22797),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    InMux I__2799 (
            .O(N__22794),
            .I(N__22791));
    LocalMux I__2798 (
            .O(N__22791),
            .I(N__22787));
    InMux I__2797 (
            .O(N__22790),
            .I(N__22784));
    Odrv4 I__2796 (
            .O(N__22787),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    LocalMux I__2795 (
            .O(N__22784),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__2794 (
            .O(N__22779),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__2793 (
            .O(N__22776),
            .I(N__22772));
    CascadeMux I__2792 (
            .O(N__22775),
            .I(N__22769));
    LocalMux I__2791 (
            .O(N__22772),
            .I(N__22766));
    InMux I__2790 (
            .O(N__22769),
            .I(N__22763));
    Odrv4 I__2789 (
            .O(N__22766),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    LocalMux I__2788 (
            .O(N__22763),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    InMux I__2787 (
            .O(N__22758),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    InMux I__2786 (
            .O(N__22755),
            .I(N__22752));
    LocalMux I__2785 (
            .O(N__22752),
            .I(N__22748));
    InMux I__2784 (
            .O(N__22751),
            .I(N__22745));
    Odrv4 I__2783 (
            .O(N__22748),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    LocalMux I__2782 (
            .O(N__22745),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    InMux I__2781 (
            .O(N__22740),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    CascadeMux I__2780 (
            .O(N__22737),
            .I(N__22734));
    InMux I__2779 (
            .O(N__22734),
            .I(N__22730));
    CascadeMux I__2778 (
            .O(N__22733),
            .I(N__22727));
    LocalMux I__2777 (
            .O(N__22730),
            .I(N__22724));
    InMux I__2776 (
            .O(N__22727),
            .I(N__22721));
    Odrv4 I__2775 (
            .O(N__22724),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    LocalMux I__2774 (
            .O(N__22721),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    InMux I__2773 (
            .O(N__22716),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    CascadeMux I__2772 (
            .O(N__22713),
            .I(N__22710));
    InMux I__2771 (
            .O(N__22710),
            .I(N__22704));
    InMux I__2770 (
            .O(N__22709),
            .I(N__22704));
    LocalMux I__2769 (
            .O(N__22704),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__2768 (
            .O(N__22701),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__2767 (
            .O(N__22698),
            .I(N__22695));
    LocalMux I__2766 (
            .O(N__22695),
            .I(N__22692));
    Odrv12 I__2765 (
            .O(N__22692),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    InMux I__2764 (
            .O(N__22689),
            .I(N__22683));
    InMux I__2763 (
            .O(N__22688),
            .I(N__22683));
    LocalMux I__2762 (
            .O(N__22683),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    InMux I__2761 (
            .O(N__22680),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__2760 (
            .O(N__22677),
            .I(N__22674));
    LocalMux I__2759 (
            .O(N__22674),
            .I(N__22670));
    InMux I__2758 (
            .O(N__22673),
            .I(N__22667));
    Odrv4 I__2757 (
            .O(N__22670),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    LocalMux I__2756 (
            .O(N__22667),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__2755 (
            .O(N__22662),
            .I(bfn_5_17_0_));
    CascadeMux I__2754 (
            .O(N__22659),
            .I(N__22656));
    InMux I__2753 (
            .O(N__22656),
            .I(N__22653));
    LocalMux I__2752 (
            .O(N__22653),
            .I(N__22649));
    InMux I__2751 (
            .O(N__22652),
            .I(N__22646));
    Odrv4 I__2750 (
            .O(N__22649),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    LocalMux I__2749 (
            .O(N__22646),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    InMux I__2748 (
            .O(N__22641),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__2747 (
            .O(N__22638),
            .I(N__22635));
    LocalMux I__2746 (
            .O(N__22635),
            .I(N__22631));
    InMux I__2745 (
            .O(N__22634),
            .I(N__22628));
    Odrv4 I__2744 (
            .O(N__22631),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    LocalMux I__2743 (
            .O(N__22628),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__2742 (
            .O(N__22623),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__2741 (
            .O(N__22620),
            .I(N__22616));
    CascadeMux I__2740 (
            .O(N__22619),
            .I(N__22613));
    LocalMux I__2739 (
            .O(N__22616),
            .I(N__22610));
    InMux I__2738 (
            .O(N__22613),
            .I(N__22607));
    Odrv4 I__2737 (
            .O(N__22610),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    LocalMux I__2736 (
            .O(N__22607),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    InMux I__2735 (
            .O(N__22602),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    InMux I__2734 (
            .O(N__22599),
            .I(N__22593));
    InMux I__2733 (
            .O(N__22598),
            .I(N__22593));
    LocalMux I__2732 (
            .O(N__22593),
            .I(N__22590));
    Odrv4 I__2731 (
            .O(N__22590),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__2730 (
            .O(N__22587),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    CascadeMux I__2729 (
            .O(N__22584),
            .I(N__22581));
    InMux I__2728 (
            .O(N__22581),
            .I(N__22578));
    LocalMux I__2727 (
            .O(N__22578),
            .I(N__22574));
    InMux I__2726 (
            .O(N__22577),
            .I(N__22571));
    Span4Mux_v I__2725 (
            .O(N__22574),
            .I(N__22565));
    LocalMux I__2724 (
            .O(N__22571),
            .I(N__22565));
    InMux I__2723 (
            .O(N__22570),
            .I(N__22562));
    Span4Mux_v I__2722 (
            .O(N__22565),
            .I(N__22559));
    LocalMux I__2721 (
            .O(N__22562),
            .I(N__22556));
    Span4Mux_h I__2720 (
            .O(N__22559),
            .I(N__22553));
    Span12Mux_s5_h I__2719 (
            .O(N__22556),
            .I(N__22550));
    Odrv4 I__2718 (
            .O(N__22553),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    Odrv12 I__2717 (
            .O(N__22550),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__2716 (
            .O(N__22545),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    CascadeMux I__2715 (
            .O(N__22542),
            .I(N__22538));
    InMux I__2714 (
            .O(N__22541),
            .I(N__22535));
    InMux I__2713 (
            .O(N__22538),
            .I(N__22532));
    LocalMux I__2712 (
            .O(N__22535),
            .I(N__22528));
    LocalMux I__2711 (
            .O(N__22532),
            .I(N__22525));
    InMux I__2710 (
            .O(N__22531),
            .I(N__22522));
    Span4Mux_h I__2709 (
            .O(N__22528),
            .I(N__22519));
    Span4Mux_s3_h I__2708 (
            .O(N__22525),
            .I(N__22514));
    LocalMux I__2707 (
            .O(N__22522),
            .I(N__22514));
    Span4Mux_v I__2706 (
            .O(N__22519),
            .I(N__22511));
    Span4Mux_v I__2705 (
            .O(N__22514),
            .I(N__22508));
    Span4Mux_v I__2704 (
            .O(N__22511),
            .I(N__22505));
    Span4Mux_v I__2703 (
            .O(N__22508),
            .I(N__22502));
    Odrv4 I__2702 (
            .O(N__22505),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    Odrv4 I__2701 (
            .O(N__22502),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__2700 (
            .O(N__22497),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__2699 (
            .O(N__22494),
            .I(N__22491));
    LocalMux I__2698 (
            .O(N__22491),
            .I(N__22486));
    InMux I__2697 (
            .O(N__22490),
            .I(N__22483));
    InMux I__2696 (
            .O(N__22489),
            .I(N__22480));
    Span4Mux_v I__2695 (
            .O(N__22486),
            .I(N__22475));
    LocalMux I__2694 (
            .O(N__22483),
            .I(N__22475));
    LocalMux I__2693 (
            .O(N__22480),
            .I(N__22472));
    Span4Mux_h I__2692 (
            .O(N__22475),
            .I(N__22469));
    Span4Mux_h I__2691 (
            .O(N__22472),
            .I(N__22466));
    Span4Mux_v I__2690 (
            .O(N__22469),
            .I(N__22463));
    Sp12to4 I__2689 (
            .O(N__22466),
            .I(N__22460));
    Odrv4 I__2688 (
            .O(N__22463),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    Odrv12 I__2687 (
            .O(N__22460),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__2686 (
            .O(N__22455),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__2685 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__2684 (
            .O(N__22449),
            .I(N__22444));
    InMux I__2683 (
            .O(N__22448),
            .I(N__22441));
    InMux I__2682 (
            .O(N__22447),
            .I(N__22438));
    Sp12to4 I__2681 (
            .O(N__22444),
            .I(N__22431));
    LocalMux I__2680 (
            .O(N__22441),
            .I(N__22431));
    LocalMux I__2679 (
            .O(N__22438),
            .I(N__22431));
    Span12Mux_v I__2678 (
            .O(N__22431),
            .I(N__22428));
    Odrv12 I__2677 (
            .O(N__22428),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    InMux I__2676 (
            .O(N__22425),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__2675 (
            .O(N__22422),
            .I(N__22417));
    InMux I__2674 (
            .O(N__22421),
            .I(N__22414));
    CascadeMux I__2673 (
            .O(N__22420),
            .I(N__22411));
    LocalMux I__2672 (
            .O(N__22417),
            .I(N__22408));
    LocalMux I__2671 (
            .O(N__22414),
            .I(N__22405));
    InMux I__2670 (
            .O(N__22411),
            .I(N__22402));
    Span4Mux_h I__2669 (
            .O(N__22408),
            .I(N__22397));
    Span4Mux_v I__2668 (
            .O(N__22405),
            .I(N__22397));
    LocalMux I__2667 (
            .O(N__22402),
            .I(N__22394));
    Span4Mux_v I__2666 (
            .O(N__22397),
            .I(N__22391));
    Span12Mux_s5_h I__2665 (
            .O(N__22394),
            .I(N__22388));
    Span4Mux_v I__2664 (
            .O(N__22391),
            .I(N__22385));
    Odrv12 I__2663 (
            .O(N__22388),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    Odrv4 I__2662 (
            .O(N__22385),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__2661 (
            .O(N__22380),
            .I(bfn_5_16_0_));
    InMux I__2660 (
            .O(N__22377),
            .I(N__22373));
    InMux I__2659 (
            .O(N__22376),
            .I(N__22370));
    LocalMux I__2658 (
            .O(N__22373),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    LocalMux I__2657 (
            .O(N__22370),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__2656 (
            .O(N__22365),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__2655 (
            .O(N__22362),
            .I(N__22358));
    InMux I__2654 (
            .O(N__22361),
            .I(N__22355));
    LocalMux I__2653 (
            .O(N__22358),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    LocalMux I__2652 (
            .O(N__22355),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    InMux I__2651 (
            .O(N__22350),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__2650 (
            .O(N__22347),
            .I(N__22344));
    LocalMux I__2649 (
            .O(N__22344),
            .I(N__22340));
    InMux I__2648 (
            .O(N__22343),
            .I(N__22337));
    Odrv12 I__2647 (
            .O(N__22340),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    LocalMux I__2646 (
            .O(N__22337),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    InMux I__2645 (
            .O(N__22332),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__2644 (
            .O(N__22329),
            .I(N__22323));
    InMux I__2643 (
            .O(N__22328),
            .I(N__22316));
    InMux I__2642 (
            .O(N__22327),
            .I(N__22316));
    InMux I__2641 (
            .O(N__22326),
            .I(N__22316));
    LocalMux I__2640 (
            .O(N__22323),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    LocalMux I__2639 (
            .O(N__22316),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    InMux I__2638 (
            .O(N__22311),
            .I(N__22308));
    LocalMux I__2637 (
            .O(N__22308),
            .I(N__22305));
    Odrv4 I__2636 (
            .O(N__22305),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__2635 (
            .O(N__22302),
            .I(N__22299));
    LocalMux I__2634 (
            .O(N__22299),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__2633 (
            .O(N__22296),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ));
    InMux I__2632 (
            .O(N__22293),
            .I(N__22290));
    LocalMux I__2631 (
            .O(N__22290),
            .I(N__22287));
    Odrv4 I__2630 (
            .O(N__22287),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    CascadeMux I__2629 (
            .O(N__22284),
            .I(N__22276));
    CascadeMux I__2628 (
            .O(N__22283),
            .I(N__22273));
    CascadeMux I__2627 (
            .O(N__22282),
            .I(N__22270));
    InMux I__2626 (
            .O(N__22281),
            .I(N__22267));
    InMux I__2625 (
            .O(N__22280),
            .I(N__22256));
    InMux I__2624 (
            .O(N__22279),
            .I(N__22256));
    InMux I__2623 (
            .O(N__22276),
            .I(N__22256));
    InMux I__2622 (
            .O(N__22273),
            .I(N__22256));
    InMux I__2621 (
            .O(N__22270),
            .I(N__22256));
    LocalMux I__2620 (
            .O(N__22267),
            .I(N__22252));
    LocalMux I__2619 (
            .O(N__22256),
            .I(N__22249));
    InMux I__2618 (
            .O(N__22255),
            .I(N__22246));
    Span4Mux_h I__2617 (
            .O(N__22252),
            .I(N__22243));
    Span4Mux_v I__2616 (
            .O(N__22249),
            .I(N__22238));
    LocalMux I__2615 (
            .O(N__22246),
            .I(N__22238));
    Span4Mux_v I__2614 (
            .O(N__22243),
            .I(N__22233));
    Span4Mux_h I__2613 (
            .O(N__22238),
            .I(N__22233));
    Span4Mux_v I__2612 (
            .O(N__22233),
            .I(N__22230));
    Odrv4 I__2611 (
            .O(N__22230),
            .I(\current_shift_inst.PI_CTRL.N_118 ));
    InMux I__2610 (
            .O(N__22227),
            .I(N__22224));
    LocalMux I__2609 (
            .O(N__22224),
            .I(N__22221));
    Span4Mux_h I__2608 (
            .O(N__22221),
            .I(N__22218));
    Sp12to4 I__2607 (
            .O(N__22218),
            .I(N__22215));
    Odrv12 I__2606 (
            .O(N__22215),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__2605 (
            .O(N__22212),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__2604 (
            .O(N__22209),
            .I(N__22205));
    InMux I__2603 (
            .O(N__22208),
            .I(N__22202));
    LocalMux I__2602 (
            .O(N__22205),
            .I(N__22196));
    LocalMux I__2601 (
            .O(N__22202),
            .I(N__22196));
    InMux I__2600 (
            .O(N__22201),
            .I(N__22193));
    Span4Mux_h I__2599 (
            .O(N__22196),
            .I(N__22190));
    LocalMux I__2598 (
            .O(N__22193),
            .I(N__22187));
    Span4Mux_v I__2597 (
            .O(N__22190),
            .I(N__22184));
    Span4Mux_h I__2596 (
            .O(N__22187),
            .I(N__22181));
    Span4Mux_v I__2595 (
            .O(N__22184),
            .I(N__22178));
    Span4Mux_v I__2594 (
            .O(N__22181),
            .I(N__22175));
    Odrv4 I__2593 (
            .O(N__22178),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    Odrv4 I__2592 (
            .O(N__22175),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__2591 (
            .O(N__22170),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__2590 (
            .O(N__22167),
            .I(N__22161));
    InMux I__2589 (
            .O(N__22166),
            .I(N__22158));
    InMux I__2588 (
            .O(N__22165),
            .I(N__22155));
    InMux I__2587 (
            .O(N__22164),
            .I(N__22152));
    LocalMux I__2586 (
            .O(N__22161),
            .I(N__22147));
    LocalMux I__2585 (
            .O(N__22158),
            .I(N__22147));
    LocalMux I__2584 (
            .O(N__22155),
            .I(N__22144));
    LocalMux I__2583 (
            .O(N__22152),
            .I(N__22141));
    Span4Mux_h I__2582 (
            .O(N__22147),
            .I(N__22138));
    Span4Mux_h I__2581 (
            .O(N__22144),
            .I(N__22135));
    Span12Mux_s5_h I__2580 (
            .O(N__22141),
            .I(N__22132));
    Span4Mux_v I__2579 (
            .O(N__22138),
            .I(N__22129));
    Span4Mux_v I__2578 (
            .O(N__22135),
            .I(N__22126));
    Odrv12 I__2577 (
            .O(N__22132),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2576 (
            .O(N__22129),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__2575 (
            .O(N__22126),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__2574 (
            .O(N__22119),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__2573 (
            .O(N__22116),
            .I(N__22113));
    LocalMux I__2572 (
            .O(N__22113),
            .I(N__22109));
    InMux I__2571 (
            .O(N__22112),
            .I(N__22105));
    Span4Mux_v I__2570 (
            .O(N__22109),
            .I(N__22102));
    InMux I__2569 (
            .O(N__22108),
            .I(N__22099));
    LocalMux I__2568 (
            .O(N__22105),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    Odrv4 I__2567 (
            .O(N__22102),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2566 (
            .O(N__22099),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2565 (
            .O(N__22092),
            .I(N__22089));
    LocalMux I__2564 (
            .O(N__22089),
            .I(N__22085));
    InMux I__2563 (
            .O(N__22088),
            .I(N__22081));
    Span4Mux_v I__2562 (
            .O(N__22085),
            .I(N__22078));
    InMux I__2561 (
            .O(N__22084),
            .I(N__22075));
    LocalMux I__2560 (
            .O(N__22081),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    Odrv4 I__2559 (
            .O(N__22078),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2558 (
            .O(N__22075),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2557 (
            .O(N__22068),
            .I(N__22065));
    LocalMux I__2556 (
            .O(N__22065),
            .I(N__22060));
    InMux I__2555 (
            .O(N__22064),
            .I(N__22057));
    InMux I__2554 (
            .O(N__22063),
            .I(N__22054));
    Span4Mux_v I__2553 (
            .O(N__22060),
            .I(N__22051));
    LocalMux I__2552 (
            .O(N__22057),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2551 (
            .O(N__22054),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    Odrv4 I__2550 (
            .O(N__22051),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2549 (
            .O(N__22044),
            .I(N__22041));
    LocalMux I__2548 (
            .O(N__22041),
            .I(N__22036));
    InMux I__2547 (
            .O(N__22040),
            .I(N__22033));
    InMux I__2546 (
            .O(N__22039),
            .I(N__22030));
    Span4Mux_v I__2545 (
            .O(N__22036),
            .I(N__22027));
    LocalMux I__2544 (
            .O(N__22033),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2543 (
            .O(N__22030),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    Odrv4 I__2542 (
            .O(N__22027),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    CascadeMux I__2541 (
            .O(N__22020),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__2540 (
            .O(N__22017),
            .I(N__22014));
    LocalMux I__2539 (
            .O(N__22014),
            .I(N__22009));
    InMux I__2538 (
            .O(N__22013),
            .I(N__22006));
    InMux I__2537 (
            .O(N__22012),
            .I(N__22003));
    Span4Mux_v I__2536 (
            .O(N__22009),
            .I(N__22000));
    LocalMux I__2535 (
            .O(N__22006),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2534 (
            .O(N__22003),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    Odrv4 I__2533 (
            .O(N__22000),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2532 (
            .O(N__21993),
            .I(N__21990));
    LocalMux I__2531 (
            .O(N__21990),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    InMux I__2530 (
            .O(N__21987),
            .I(N__21984));
    LocalMux I__2529 (
            .O(N__21984),
            .I(N__21979));
    InMux I__2528 (
            .O(N__21983),
            .I(N__21976));
    InMux I__2527 (
            .O(N__21982),
            .I(N__21973));
    Span4Mux_v I__2526 (
            .O(N__21979),
            .I(N__21970));
    LocalMux I__2525 (
            .O(N__21976),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2524 (
            .O(N__21973),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    Odrv4 I__2523 (
            .O(N__21970),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    CascadeMux I__2522 (
            .O(N__21963),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__2521 (
            .O(N__21960),
            .I(N__21957));
    LocalMux I__2520 (
            .O(N__21957),
            .I(N__21952));
    InMux I__2519 (
            .O(N__21956),
            .I(N__21949));
    InMux I__2518 (
            .O(N__21955),
            .I(N__21946));
    Span4Mux_v I__2517 (
            .O(N__21952),
            .I(N__21943));
    LocalMux I__2516 (
            .O(N__21949),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2515 (
            .O(N__21946),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    Odrv4 I__2514 (
            .O(N__21943),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2513 (
            .O(N__21936),
            .I(N__21918));
    InMux I__2512 (
            .O(N__21935),
            .I(N__21918));
    InMux I__2511 (
            .O(N__21934),
            .I(N__21918));
    InMux I__2510 (
            .O(N__21933),
            .I(N__21918));
    InMux I__2509 (
            .O(N__21932),
            .I(N__21913));
    InMux I__2508 (
            .O(N__21931),
            .I(N__21913));
    InMux I__2507 (
            .O(N__21930),
            .I(N__21904));
    InMux I__2506 (
            .O(N__21929),
            .I(N__21904));
    InMux I__2505 (
            .O(N__21928),
            .I(N__21904));
    InMux I__2504 (
            .O(N__21927),
            .I(N__21904));
    LocalMux I__2503 (
            .O(N__21918),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2502 (
            .O(N__21913),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2501 (
            .O(N__21904),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2500 (
            .O(N__21897),
            .I(N__21894));
    LocalMux I__2499 (
            .O(N__21894),
            .I(N__21891));
    Span4Mux_h I__2498 (
            .O(N__21891),
            .I(N__21888));
    Span4Mux_v I__2497 (
            .O(N__21888),
            .I(N__21885));
    Span4Mux_v I__2496 (
            .O(N__21885),
            .I(N__21882));
    Span4Mux_v I__2495 (
            .O(N__21882),
            .I(N__21879));
    Odrv4 I__2494 (
            .O(N__21879),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    CascadeMux I__2493 (
            .O(N__21876),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    CascadeMux I__2492 (
            .O(N__21873),
            .I(N__21870));
    InMux I__2491 (
            .O(N__21870),
            .I(N__21867));
    LocalMux I__2490 (
            .O(N__21867),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    CascadeMux I__2489 (
            .O(N__21864),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ));
    InMux I__2488 (
            .O(N__21861),
            .I(N__21858));
    LocalMux I__2487 (
            .O(N__21858),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    CascadeMux I__2486 (
            .O(N__21855),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__2485 (
            .O(N__21852),
            .I(N__21849));
    LocalMux I__2484 (
            .O(N__21849),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__2483 (
            .O(N__21846),
            .I(N__21843));
    LocalMux I__2482 (
            .O(N__21843),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ));
    InMux I__2481 (
            .O(N__21840),
            .I(N__21837));
    LocalMux I__2480 (
            .O(N__21837),
            .I(N__21834));
    Odrv4 I__2479 (
            .O(N__21834),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    InMux I__2478 (
            .O(N__21831),
            .I(N__21828));
    LocalMux I__2477 (
            .O(N__21828),
            .I(N__21824));
    InMux I__2476 (
            .O(N__21827),
            .I(N__21820));
    Span4Mux_v I__2475 (
            .O(N__21824),
            .I(N__21817));
    InMux I__2474 (
            .O(N__21823),
            .I(N__21814));
    LocalMux I__2473 (
            .O(N__21820),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2472 (
            .O(N__21817),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2471 (
            .O(N__21814),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2470 (
            .O(N__21807),
            .I(N__21804));
    LocalMux I__2469 (
            .O(N__21804),
            .I(N__21800));
    InMux I__2468 (
            .O(N__21803),
            .I(N__21796));
    Span4Mux_v I__2467 (
            .O(N__21800),
            .I(N__21793));
    InMux I__2466 (
            .O(N__21799),
            .I(N__21790));
    LocalMux I__2465 (
            .O(N__21796),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2464 (
            .O(N__21793),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2463 (
            .O(N__21790),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2462 (
            .O(N__21783),
            .I(N__21780));
    LocalMux I__2461 (
            .O(N__21780),
            .I(N__21775));
    InMux I__2460 (
            .O(N__21779),
            .I(N__21772));
    InMux I__2459 (
            .O(N__21778),
            .I(N__21769));
    Span4Mux_v I__2458 (
            .O(N__21775),
            .I(N__21766));
    LocalMux I__2457 (
            .O(N__21772),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2456 (
            .O(N__21769),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    Odrv4 I__2455 (
            .O(N__21766),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2454 (
            .O(N__21759),
            .I(N__21756));
    LocalMux I__2453 (
            .O(N__21756),
            .I(\pwm_generator_inst.counter_i_9 ));
    InMux I__2452 (
            .O(N__21753),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2451 (
            .O(N__21750),
            .I(N__21747));
    LocalMux I__2450 (
            .O(N__21747),
            .I(N__21744));
    Span12Mux_s1_v I__2449 (
            .O(N__21744),
            .I(N__21741));
    Span12Mux_h I__2448 (
            .O(N__21741),
            .I(N__21738));
    Span12Mux_v I__2447 (
            .O(N__21738),
            .I(N__21735));
    Odrv12 I__2446 (
            .O(N__21735),
            .I(pwm_output_c));
    CascadeMux I__2445 (
            .O(N__21732),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    CascadeMux I__2444 (
            .O(N__21729),
            .I(N__21726));
    InMux I__2443 (
            .O(N__21726),
            .I(N__21723));
    LocalMux I__2442 (
            .O(N__21723),
            .I(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ));
    CascadeMux I__2441 (
            .O(N__21720),
            .I(N__21717));
    InMux I__2440 (
            .O(N__21717),
            .I(N__21714));
    LocalMux I__2439 (
            .O(N__21714),
            .I(\pwm_generator_inst.un14_counter_8 ));
    InMux I__2438 (
            .O(N__21711),
            .I(N__21705));
    InMux I__2437 (
            .O(N__21710),
            .I(N__21705));
    LocalMux I__2436 (
            .O(N__21705),
            .I(N__21694));
    InMux I__2435 (
            .O(N__21704),
            .I(N__21677));
    InMux I__2434 (
            .O(N__21703),
            .I(N__21677));
    InMux I__2433 (
            .O(N__21702),
            .I(N__21677));
    InMux I__2432 (
            .O(N__21701),
            .I(N__21677));
    InMux I__2431 (
            .O(N__21700),
            .I(N__21677));
    InMux I__2430 (
            .O(N__21699),
            .I(N__21677));
    InMux I__2429 (
            .O(N__21698),
            .I(N__21677));
    InMux I__2428 (
            .O(N__21697),
            .I(N__21677));
    Span4Mux_v I__2427 (
            .O(N__21694),
            .I(N__21672));
    LocalMux I__2426 (
            .O(N__21677),
            .I(N__21672));
    Span4Mux_v I__2425 (
            .O(N__21672),
            .I(N__21669));
    Span4Mux_v I__2424 (
            .O(N__21669),
            .I(N__21666));
    Odrv4 I__2423 (
            .O(N__21666),
            .I(\pwm_generator_inst.N_17 ));
    InMux I__2422 (
            .O(N__21663),
            .I(N__21657));
    InMux I__2421 (
            .O(N__21662),
            .I(N__21657));
    LocalMux I__2420 (
            .O(N__21657),
            .I(N__21646));
    InMux I__2419 (
            .O(N__21656),
            .I(N__21629));
    InMux I__2418 (
            .O(N__21655),
            .I(N__21629));
    InMux I__2417 (
            .O(N__21654),
            .I(N__21629));
    InMux I__2416 (
            .O(N__21653),
            .I(N__21629));
    InMux I__2415 (
            .O(N__21652),
            .I(N__21629));
    InMux I__2414 (
            .O(N__21651),
            .I(N__21629));
    InMux I__2413 (
            .O(N__21650),
            .I(N__21629));
    InMux I__2412 (
            .O(N__21649),
            .I(N__21629));
    Span4Mux_v I__2411 (
            .O(N__21646),
            .I(N__21626));
    LocalMux I__2410 (
            .O(N__21629),
            .I(N__21623));
    Span4Mux_v I__2409 (
            .O(N__21626),
            .I(N__21620));
    Span12Mux_v I__2408 (
            .O(N__21623),
            .I(N__21617));
    Odrv4 I__2407 (
            .O(N__21620),
            .I(\pwm_generator_inst.N_16 ));
    Odrv12 I__2406 (
            .O(N__21617),
            .I(\pwm_generator_inst.N_16 ));
    CascadeMux I__2405 (
            .O(N__21612),
            .I(N__21608));
    InMux I__2404 (
            .O(N__21611),
            .I(N__21583));
    InMux I__2403 (
            .O(N__21608),
            .I(N__21583));
    CascadeMux I__2402 (
            .O(N__21607),
            .I(N__21579));
    CascadeMux I__2401 (
            .O(N__21606),
            .I(N__21575));
    CascadeMux I__2400 (
            .O(N__21605),
            .I(N__21571));
    CascadeMux I__2399 (
            .O(N__21604),
            .I(N__21567));
    CascadeMux I__2398 (
            .O(N__21603),
            .I(N__21559));
    InMux I__2397 (
            .O(N__21602),
            .I(N__21541));
    InMux I__2396 (
            .O(N__21601),
            .I(N__21541));
    InMux I__2395 (
            .O(N__21600),
            .I(N__21541));
    InMux I__2394 (
            .O(N__21599),
            .I(N__21541));
    InMux I__2393 (
            .O(N__21598),
            .I(N__21541));
    InMux I__2392 (
            .O(N__21597),
            .I(N__21541));
    InMux I__2391 (
            .O(N__21596),
            .I(N__21541));
    InMux I__2390 (
            .O(N__21595),
            .I(N__21541));
    InMux I__2389 (
            .O(N__21594),
            .I(N__21526));
    InMux I__2388 (
            .O(N__21593),
            .I(N__21526));
    InMux I__2387 (
            .O(N__21592),
            .I(N__21526));
    InMux I__2386 (
            .O(N__21591),
            .I(N__21526));
    InMux I__2385 (
            .O(N__21590),
            .I(N__21526));
    InMux I__2384 (
            .O(N__21589),
            .I(N__21526));
    InMux I__2383 (
            .O(N__21588),
            .I(N__21526));
    LocalMux I__2382 (
            .O(N__21583),
            .I(N__21523));
    InMux I__2381 (
            .O(N__21582),
            .I(N__21506));
    InMux I__2380 (
            .O(N__21579),
            .I(N__21506));
    InMux I__2379 (
            .O(N__21578),
            .I(N__21506));
    InMux I__2378 (
            .O(N__21575),
            .I(N__21506));
    InMux I__2377 (
            .O(N__21574),
            .I(N__21506));
    InMux I__2376 (
            .O(N__21571),
            .I(N__21506));
    InMux I__2375 (
            .O(N__21570),
            .I(N__21506));
    InMux I__2374 (
            .O(N__21567),
            .I(N__21506));
    InMux I__2373 (
            .O(N__21566),
            .I(N__21501));
    InMux I__2372 (
            .O(N__21565),
            .I(N__21501));
    InMux I__2371 (
            .O(N__21564),
            .I(N__21494));
    InMux I__2370 (
            .O(N__21563),
            .I(N__21494));
    InMux I__2369 (
            .O(N__21562),
            .I(N__21494));
    InMux I__2368 (
            .O(N__21559),
            .I(N__21491));
    InMux I__2367 (
            .O(N__21558),
            .I(N__21488));
    LocalMux I__2366 (
            .O(N__21541),
            .I(N__21485));
    LocalMux I__2365 (
            .O(N__21526),
            .I(N__21482));
    Span4Mux_v I__2364 (
            .O(N__21523),
            .I(N__21477));
    LocalMux I__2363 (
            .O(N__21506),
            .I(N__21477));
    LocalMux I__2362 (
            .O(N__21501),
            .I(N__21472));
    LocalMux I__2361 (
            .O(N__21494),
            .I(N__21472));
    LocalMux I__2360 (
            .O(N__21491),
            .I(N__21463));
    LocalMux I__2359 (
            .O(N__21488),
            .I(N__21463));
    Sp12to4 I__2358 (
            .O(N__21485),
            .I(N__21463));
    Sp12to4 I__2357 (
            .O(N__21482),
            .I(N__21463));
    Span4Mux_h I__2356 (
            .O(N__21477),
            .I(N__21460));
    Sp12to4 I__2355 (
            .O(N__21472),
            .I(N__21455));
    Span12Mux_v I__2354 (
            .O(N__21463),
            .I(N__21455));
    Odrv4 I__2353 (
            .O(N__21460),
            .I(N_19_1));
    Odrv12 I__2352 (
            .O(N__21455),
            .I(N_19_1));
    InMux I__2351 (
            .O(N__21450),
            .I(N__21447));
    LocalMux I__2350 (
            .O(N__21447),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ));
    CascadeMux I__2349 (
            .O(N__21444),
            .I(N__21441));
    InMux I__2348 (
            .O(N__21441),
            .I(N__21438));
    LocalMux I__2347 (
            .O(N__21438),
            .I(\pwm_generator_inst.threshold_9 ));
    InMux I__2346 (
            .O(N__21435),
            .I(N__21432));
    LocalMux I__2345 (
            .O(N__21432),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    CascadeMux I__2344 (
            .O(N__21429),
            .I(N__21426));
    InMux I__2343 (
            .O(N__21426),
            .I(N__21423));
    LocalMux I__2342 (
            .O(N__21423),
            .I(\pwm_generator_inst.threshold_2 ));
    InMux I__2341 (
            .O(N__21420),
            .I(N__21417));
    LocalMux I__2340 (
            .O(N__21417),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2339 (
            .O(N__21414),
            .I(N__21411));
    InMux I__2338 (
            .O(N__21411),
            .I(N__21408));
    LocalMux I__2337 (
            .O(N__21408),
            .I(N__21405));
    Odrv4 I__2336 (
            .O(N__21405),
            .I(\pwm_generator_inst.threshold_3 ));
    InMux I__2335 (
            .O(N__21402),
            .I(N__21399));
    LocalMux I__2334 (
            .O(N__21399),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2333 (
            .O(N__21396),
            .I(N__21393));
    InMux I__2332 (
            .O(N__21393),
            .I(N__21390));
    LocalMux I__2331 (
            .O(N__21390),
            .I(\pwm_generator_inst.threshold_4 ));
    InMux I__2330 (
            .O(N__21387),
            .I(N__21384));
    LocalMux I__2329 (
            .O(N__21384),
            .I(\pwm_generator_inst.counter_i_4 ));
    CascadeMux I__2328 (
            .O(N__21381),
            .I(N__21378));
    InMux I__2327 (
            .O(N__21378),
            .I(N__21375));
    LocalMux I__2326 (
            .O(N__21375),
            .I(\pwm_generator_inst.threshold_5 ));
    InMux I__2325 (
            .O(N__21372),
            .I(N__21369));
    LocalMux I__2324 (
            .O(N__21369),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2323 (
            .O(N__21366),
            .I(N__21363));
    InMux I__2322 (
            .O(N__21363),
            .I(N__21360));
    LocalMux I__2321 (
            .O(N__21360),
            .I(\pwm_generator_inst.un14_counter_6 ));
    InMux I__2320 (
            .O(N__21357),
            .I(N__21354));
    LocalMux I__2319 (
            .O(N__21354),
            .I(\pwm_generator_inst.counter_i_6 ));
    InMux I__2318 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__2317 (
            .O(N__21348),
            .I(\pwm_generator_inst.un14_counter_7 ));
    CascadeMux I__2316 (
            .O(N__21345),
            .I(N__21342));
    InMux I__2315 (
            .O(N__21342),
            .I(N__21339));
    LocalMux I__2314 (
            .O(N__21339),
            .I(\pwm_generator_inst.counter_i_7 ));
    InMux I__2313 (
            .O(N__21336),
            .I(N__21333));
    LocalMux I__2312 (
            .O(N__21333),
            .I(\pwm_generator_inst.counter_i_8 ));
    InMux I__2311 (
            .O(N__21330),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2310 (
            .O(N__21327),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2309 (
            .O(N__21324),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2308 (
            .O(N__21321),
            .I(bfn_3_19_0_));
    InMux I__2307 (
            .O(N__21318),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2306 (
            .O(N__21315),
            .I(N__21312));
    LocalMux I__2305 (
            .O(N__21312),
            .I(N__21309));
    Span4Mux_h I__2304 (
            .O(N__21309),
            .I(N__21306));
    Span4Mux_v I__2303 (
            .O(N__21306),
            .I(N__21303));
    Odrv4 I__2302 (
            .O(N__21303),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__2301 (
            .O(N__21300),
            .I(N__21297));
    InMux I__2300 (
            .O(N__21297),
            .I(N__21294));
    LocalMux I__2299 (
            .O(N__21294),
            .I(N__21291));
    Odrv4 I__2298 (
            .O(N__21291),
            .I(\pwm_generator_inst.threshold_0 ));
    InMux I__2297 (
            .O(N__21288),
            .I(N__21285));
    LocalMux I__2296 (
            .O(N__21285),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2295 (
            .O(N__21282),
            .I(N__21279));
    InMux I__2294 (
            .O(N__21279),
            .I(N__21276));
    LocalMux I__2293 (
            .O(N__21276),
            .I(\pwm_generator_inst.un14_counter_1 ));
    InMux I__2292 (
            .O(N__21273),
            .I(N__21270));
    LocalMux I__2291 (
            .O(N__21270),
            .I(\pwm_generator_inst.counter_i_1 ));
    InMux I__2290 (
            .O(N__21267),
            .I(N__21264));
    LocalMux I__2289 (
            .O(N__21264),
            .I(N__21261));
    Odrv4 I__2288 (
            .O(N__21261),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ));
    InMux I__2287 (
            .O(N__21258),
            .I(N__21255));
    LocalMux I__2286 (
            .O(N__21255),
            .I(N__21250));
    InMux I__2285 (
            .O(N__21254),
            .I(N__21247));
    InMux I__2284 (
            .O(N__21253),
            .I(N__21244));
    Span4Mux_h I__2283 (
            .O(N__21250),
            .I(N__21239));
    LocalMux I__2282 (
            .O(N__21247),
            .I(N__21239));
    LocalMux I__2281 (
            .O(N__21244),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    Odrv4 I__2280 (
            .O(N__21239),
            .I(\pwm_generator_inst.un15_threshold_1_axb_13 ));
    CascadeMux I__2279 (
            .O(N__21234),
            .I(N__21231));
    InMux I__2278 (
            .O(N__21231),
            .I(N__21228));
    LocalMux I__2277 (
            .O(N__21228),
            .I(N__21224));
    InMux I__2276 (
            .O(N__21227),
            .I(N__21221));
    Odrv4 I__2275 (
            .O(N__21224),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    LocalMux I__2274 (
            .O(N__21221),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ));
    InMux I__2273 (
            .O(N__21216),
            .I(N__21213));
    LocalMux I__2272 (
            .O(N__21213),
            .I(\pwm_generator_inst.un19_threshold_axb_3 ));
    InMux I__2271 (
            .O(N__21210),
            .I(N__21207));
    LocalMux I__2270 (
            .O(N__21207),
            .I(N__21203));
    InMux I__2269 (
            .O(N__21206),
            .I(N__21199));
    Span4Mux_v I__2268 (
            .O(N__21203),
            .I(N__21196));
    InMux I__2267 (
            .O(N__21202),
            .I(N__21193));
    LocalMux I__2266 (
            .O(N__21199),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    Odrv4 I__2265 (
            .O(N__21196),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    LocalMux I__2264 (
            .O(N__21193),
            .I(\pwm_generator_inst.un15_threshold_1_axb_10 ));
    InMux I__2263 (
            .O(N__21186),
            .I(N__21183));
    LocalMux I__2262 (
            .O(N__21183),
            .I(N__21180));
    Odrv4 I__2261 (
            .O(N__21180),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ));
    CascadeMux I__2260 (
            .O(N__21177),
            .I(N__21174));
    InMux I__2259 (
            .O(N__21174),
            .I(N__21171));
    LocalMux I__2258 (
            .O(N__21171),
            .I(N__21167));
    InMux I__2257 (
            .O(N__21170),
            .I(N__21164));
    Span4Mux_h I__2256 (
            .O(N__21167),
            .I(N__21161));
    LocalMux I__2255 (
            .O(N__21164),
            .I(N__21158));
    Sp12to4 I__2254 (
            .O(N__21161),
            .I(N__21155));
    Span4Mux_v I__2253 (
            .O(N__21158),
            .I(N__21152));
    Odrv12 I__2252 (
            .O(N__21155),
            .I(\pwm_generator_inst.O_10 ));
    Odrv4 I__2251 (
            .O(N__21152),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__2250 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__2249 (
            .O(N__21144),
            .I(\pwm_generator_inst.un19_threshold_axb_0 ));
    InMux I__2248 (
            .O(N__21141),
            .I(N__21138));
    LocalMux I__2247 (
            .O(N__21138),
            .I(N__21135));
    Odrv4 I__2246 (
            .O(N__21135),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ));
    InMux I__2245 (
            .O(N__21132),
            .I(N__21128));
    InMux I__2244 (
            .O(N__21131),
            .I(N__21125));
    LocalMux I__2243 (
            .O(N__21128),
            .I(N__21122));
    LocalMux I__2242 (
            .O(N__21125),
            .I(N__21119));
    Odrv4 I__2241 (
            .O(N__21122),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    Odrv4 I__2240 (
            .O(N__21119),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ));
    CascadeMux I__2239 (
            .O(N__21114),
            .I(N__21107));
    InMux I__2238 (
            .O(N__21113),
            .I(N__21104));
    CascadeMux I__2237 (
            .O(N__21112),
            .I(N__21100));
    CascadeMux I__2236 (
            .O(N__21111),
            .I(N__21092));
    InMux I__2235 (
            .O(N__21110),
            .I(N__21088));
    InMux I__2234 (
            .O(N__21107),
            .I(N__21085));
    LocalMux I__2233 (
            .O(N__21104),
            .I(N__21082));
    InMux I__2232 (
            .O(N__21103),
            .I(N__21077));
    InMux I__2231 (
            .O(N__21100),
            .I(N__21077));
    InMux I__2230 (
            .O(N__21099),
            .I(N__21070));
    InMux I__2229 (
            .O(N__21098),
            .I(N__21070));
    InMux I__2228 (
            .O(N__21097),
            .I(N__21070));
    InMux I__2227 (
            .O(N__21096),
            .I(N__21061));
    InMux I__2226 (
            .O(N__21095),
            .I(N__21061));
    InMux I__2225 (
            .O(N__21092),
            .I(N__21061));
    InMux I__2224 (
            .O(N__21091),
            .I(N__21061));
    LocalMux I__2223 (
            .O(N__21088),
            .I(N__21054));
    LocalMux I__2222 (
            .O(N__21085),
            .I(N__21054));
    Span4Mux_s3_h I__2221 (
            .O(N__21082),
            .I(N__21054));
    LocalMux I__2220 (
            .O(N__21077),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__2219 (
            .O(N__21070),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    LocalMux I__2218 (
            .O(N__21061),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    Odrv4 I__2217 (
            .O(N__21054),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ));
    InMux I__2216 (
            .O(N__21045),
            .I(N__21041));
    InMux I__2215 (
            .O(N__21044),
            .I(N__21037));
    LocalMux I__2214 (
            .O(N__21041),
            .I(N__21034));
    InMux I__2213 (
            .O(N__21040),
            .I(N__21031));
    LocalMux I__2212 (
            .O(N__21037),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    Odrv4 I__2211 (
            .O(N__21034),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    LocalMux I__2210 (
            .O(N__21031),
            .I(\pwm_generator_inst.un15_threshold_1_axb_12 ));
    InMux I__2209 (
            .O(N__21024),
            .I(N__21021));
    LocalMux I__2208 (
            .O(N__21021),
            .I(\pwm_generator_inst.un19_threshold_axb_2 ));
    InMux I__2207 (
            .O(N__21018),
            .I(N__21011));
    InMux I__2206 (
            .O(N__21017),
            .I(N__21001));
    InMux I__2205 (
            .O(N__21016),
            .I(N__21001));
    InMux I__2204 (
            .O(N__21015),
            .I(N__21001));
    InMux I__2203 (
            .O(N__21014),
            .I(N__21001));
    LocalMux I__2202 (
            .O(N__21011),
            .I(N__20998));
    InMux I__2201 (
            .O(N__21010),
            .I(N__20995));
    LocalMux I__2200 (
            .O(N__21001),
            .I(N__20988));
    Span4Mux_v I__2199 (
            .O(N__20998),
            .I(N__20988));
    LocalMux I__2198 (
            .O(N__20995),
            .I(N__20985));
    InMux I__2197 (
            .O(N__20994),
            .I(N__20980));
    InMux I__2196 (
            .O(N__20993),
            .I(N__20980));
    Sp12to4 I__2195 (
            .O(N__20988),
            .I(N__20977));
    Span4Mux_s3_h I__2194 (
            .O(N__20985),
            .I(N__20974));
    LocalMux I__2193 (
            .O(N__20980),
            .I(N__20971));
    Span12Mux_s3_h I__2192 (
            .O(N__20977),
            .I(N__20964));
    Sp12to4 I__2191 (
            .O(N__20974),
            .I(N__20964));
    Sp12to4 I__2190 (
            .O(N__20971),
            .I(N__20964));
    Odrv12 I__2189 (
            .O(N__20964),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ));
    InMux I__2188 (
            .O(N__20961),
            .I(bfn_3_18_0_));
    InMux I__2187 (
            .O(N__20958),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2186 (
            .O(N__20955),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2185 (
            .O(N__20952),
            .I(\pwm_generator_inst.counter_cry_2 ));
    InMux I__2184 (
            .O(N__20949),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2183 (
            .O(N__20946),
            .I(N__20943));
    LocalMux I__2182 (
            .O(N__20943),
            .I(N__20940));
    Odrv4 I__2181 (
            .O(N__20940),
            .I(\pwm_generator_inst.un19_threshold_axb_4 ));
    CascadeMux I__2180 (
            .O(N__20937),
            .I(N__20934));
    InMux I__2179 (
            .O(N__20934),
            .I(N__20931));
    LocalMux I__2178 (
            .O(N__20931),
            .I(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ));
    InMux I__2177 (
            .O(N__20928),
            .I(\pwm_generator_inst.un19_threshold_cry_3 ));
    InMux I__2176 (
            .O(N__20925),
            .I(N__20922));
    LocalMux I__2175 (
            .O(N__20922),
            .I(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ));
    InMux I__2174 (
            .O(N__20919),
            .I(\pwm_generator_inst.un19_threshold_cry_4 ));
    InMux I__2173 (
            .O(N__20916),
            .I(N__20913));
    LocalMux I__2172 (
            .O(N__20913),
            .I(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ));
    InMux I__2171 (
            .O(N__20910),
            .I(\pwm_generator_inst.un19_threshold_cry_5 ));
    InMux I__2170 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__2169 (
            .O(N__20904),
            .I(N__20901));
    Odrv4 I__2168 (
            .O(N__20901),
            .I(\pwm_generator_inst.un19_threshold_axb_7 ));
    CascadeMux I__2167 (
            .O(N__20898),
            .I(N__20895));
    InMux I__2166 (
            .O(N__20895),
            .I(N__20892));
    LocalMux I__2165 (
            .O(N__20892),
            .I(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ));
    InMux I__2164 (
            .O(N__20889),
            .I(\pwm_generator_inst.un19_threshold_cry_6 ));
    InMux I__2163 (
            .O(N__20886),
            .I(N__20883));
    LocalMux I__2162 (
            .O(N__20883),
            .I(\pwm_generator_inst.un19_threshold_axb_8 ));
    InMux I__2161 (
            .O(N__20880),
            .I(bfn_3_16_0_));
    InMux I__2160 (
            .O(N__20877),
            .I(N__20874));
    LocalMux I__2159 (
            .O(N__20874),
            .I(N__20871));
    Span4Mux_v I__2158 (
            .O(N__20871),
            .I(N__20868));
    Odrv4 I__2157 (
            .O(N__20868),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ));
    CascadeMux I__2156 (
            .O(N__20865),
            .I(N__20862));
    InMux I__2155 (
            .O(N__20862),
            .I(N__20859));
    LocalMux I__2154 (
            .O(N__20859),
            .I(N__20856));
    Odrv4 I__2153 (
            .O(N__20856),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ));
    InMux I__2152 (
            .O(N__20853),
            .I(\pwm_generator_inst.un19_threshold_cry_8 ));
    InMux I__2151 (
            .O(N__20850),
            .I(N__20847));
    LocalMux I__2150 (
            .O(N__20847),
            .I(N__20844));
    Odrv4 I__2149 (
            .O(N__20844),
            .I(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ));
    InMux I__2148 (
            .O(N__20841),
            .I(N__20838));
    LocalMux I__2147 (
            .O(N__20838),
            .I(N__20833));
    InMux I__2146 (
            .O(N__20837),
            .I(N__20828));
    InMux I__2145 (
            .O(N__20836),
            .I(N__20828));
    Odrv4 I__2144 (
            .O(N__20833),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    LocalMux I__2143 (
            .O(N__20828),
            .I(\pwm_generator_inst.un15_threshold_1_axb_16 ));
    InMux I__2142 (
            .O(N__20823),
            .I(N__20819));
    InMux I__2141 (
            .O(N__20822),
            .I(N__20816));
    LocalMux I__2140 (
            .O(N__20819),
            .I(N__20813));
    LocalMux I__2139 (
            .O(N__20816),
            .I(N__20810));
    Odrv4 I__2138 (
            .O(N__20813),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    Odrv4 I__2137 (
            .O(N__20810),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ));
    InMux I__2136 (
            .O(N__20805),
            .I(N__20802));
    LocalMux I__2135 (
            .O(N__20802),
            .I(\pwm_generator_inst.un19_threshold_axb_6 ));
    InMux I__2134 (
            .O(N__20799),
            .I(N__20796));
    LocalMux I__2133 (
            .O(N__20796),
            .I(N__20793));
    Odrv4 I__2132 (
            .O(N__20793),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ));
    CascadeMux I__2131 (
            .O(N__20790),
            .I(N__20787));
    InMux I__2130 (
            .O(N__20787),
            .I(N__20784));
    LocalMux I__2129 (
            .O(N__20784),
            .I(N__20780));
    InMux I__2128 (
            .O(N__20783),
            .I(N__20776));
    Span4Mux_v I__2127 (
            .O(N__20780),
            .I(N__20773));
    InMux I__2126 (
            .O(N__20779),
            .I(N__20770));
    LocalMux I__2125 (
            .O(N__20776),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    Odrv4 I__2124 (
            .O(N__20773),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    LocalMux I__2123 (
            .O(N__20770),
            .I(\pwm_generator_inst.un15_threshold_1_axb_15 ));
    InMux I__2122 (
            .O(N__20763),
            .I(N__20759));
    InMux I__2121 (
            .O(N__20762),
            .I(N__20756));
    LocalMux I__2120 (
            .O(N__20759),
            .I(N__20753));
    LocalMux I__2119 (
            .O(N__20756),
            .I(N__20750));
    Odrv12 I__2118 (
            .O(N__20753),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    Odrv4 I__2117 (
            .O(N__20750),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ));
    InMux I__2116 (
            .O(N__20745),
            .I(N__20742));
    LocalMux I__2115 (
            .O(N__20742),
            .I(\pwm_generator_inst.un19_threshold_axb_5 ));
    CascadeMux I__2114 (
            .O(N__20739),
            .I(N__20736));
    InMux I__2113 (
            .O(N__20736),
            .I(N__20733));
    LocalMux I__2112 (
            .O(N__20733),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ));
    InMux I__2111 (
            .O(N__20730),
            .I(N__20727));
    LocalMux I__2110 (
            .O(N__20727),
            .I(N__20724));
    Odrv4 I__2109 (
            .O(N__20724),
            .I(\pwm_generator_inst.un19_threshold_axb_1 ));
    InMux I__2108 (
            .O(N__20721),
            .I(N__20718));
    LocalMux I__2107 (
            .O(N__20718),
            .I(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ));
    InMux I__2106 (
            .O(N__20715),
            .I(\pwm_generator_inst.un19_threshold_cry_0 ));
    CascadeMux I__2105 (
            .O(N__20712),
            .I(N__20709));
    InMux I__2104 (
            .O(N__20709),
            .I(N__20706));
    LocalMux I__2103 (
            .O(N__20706),
            .I(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ));
    InMux I__2102 (
            .O(N__20703),
            .I(\pwm_generator_inst.un19_threshold_cry_1 ));
    InMux I__2101 (
            .O(N__20700),
            .I(N__20697));
    LocalMux I__2100 (
            .O(N__20697),
            .I(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ));
    InMux I__2099 (
            .O(N__20694),
            .I(\pwm_generator_inst.un19_threshold_cry_2 ));
    InMux I__2098 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__2097 (
            .O(N__20688),
            .I(N__20685));
    Odrv12 I__2096 (
            .O(N__20685),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ));
    InMux I__2095 (
            .O(N__20682),
            .I(N__20678));
    InMux I__2094 (
            .O(N__20681),
            .I(N__20675));
    LocalMux I__2093 (
            .O(N__20678),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    LocalMux I__2092 (
            .O(N__20675),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ));
    CascadeMux I__2091 (
            .O(N__20670),
            .I(N__20667));
    InMux I__2090 (
            .O(N__20667),
            .I(N__20662));
    InMux I__2089 (
            .O(N__20666),
            .I(N__20659));
    InMux I__2088 (
            .O(N__20665),
            .I(N__20656));
    LocalMux I__2087 (
            .O(N__20662),
            .I(N__20653));
    LocalMux I__2086 (
            .O(N__20659),
            .I(N__20650));
    LocalMux I__2085 (
            .O(N__20656),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__2084 (
            .O(N__20653),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    Odrv4 I__2083 (
            .O(N__20650),
            .I(\pwm_generator_inst.un15_threshold_1_axb_14 ));
    InMux I__2082 (
            .O(N__20643),
            .I(N__20638));
    InMux I__2081 (
            .O(N__20642),
            .I(N__20635));
    InMux I__2080 (
            .O(N__20641),
            .I(N__20632));
    LocalMux I__2079 (
            .O(N__20638),
            .I(N__20629));
    LocalMux I__2078 (
            .O(N__20635),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    LocalMux I__2077 (
            .O(N__20632),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    Odrv4 I__2076 (
            .O(N__20629),
            .I(\pwm_generator_inst.un15_threshold_1_axb_18 ));
    InMux I__2075 (
            .O(N__20622),
            .I(N__20618));
    InMux I__2074 (
            .O(N__20621),
            .I(N__20615));
    LocalMux I__2073 (
            .O(N__20618),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    LocalMux I__2072 (
            .O(N__20615),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ));
    CascadeMux I__2071 (
            .O(N__20610),
            .I(N__20607));
    InMux I__2070 (
            .O(N__20607),
            .I(N__20604));
    LocalMux I__2069 (
            .O(N__20604),
            .I(N__20601));
    Odrv4 I__2068 (
            .O(N__20601),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ));
    InMux I__2067 (
            .O(N__20598),
            .I(N__20595));
    LocalMux I__2066 (
            .O(N__20595),
            .I(N__20592));
    Odrv12 I__2065 (
            .O(N__20592),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ));
    InMux I__2064 (
            .O(N__20589),
            .I(N__20585));
    InMux I__2063 (
            .O(N__20588),
            .I(N__20582));
    LocalMux I__2062 (
            .O(N__20585),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    LocalMux I__2061 (
            .O(N__20582),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ));
    CascadeMux I__2060 (
            .O(N__20577),
            .I(N__20574));
    InMux I__2059 (
            .O(N__20574),
            .I(N__20570));
    InMux I__2058 (
            .O(N__20573),
            .I(N__20566));
    LocalMux I__2057 (
            .O(N__20570),
            .I(N__20563));
    InMux I__2056 (
            .O(N__20569),
            .I(N__20560));
    LocalMux I__2055 (
            .O(N__20566),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    Odrv4 I__2054 (
            .O(N__20563),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    LocalMux I__2053 (
            .O(N__20560),
            .I(\pwm_generator_inst.un15_threshold_1_axb_17 ));
    InMux I__2052 (
            .O(N__20553),
            .I(N__20550));
    LocalMux I__2051 (
            .O(N__20550),
            .I(\pwm_generator_inst.un1_duty_inputlt3 ));
    InMux I__2050 (
            .O(N__20547),
            .I(N__20543));
    InMux I__2049 (
            .O(N__20546),
            .I(N__20539));
    LocalMux I__2048 (
            .O(N__20543),
            .I(N__20536));
    InMux I__2047 (
            .O(N__20542),
            .I(N__20533));
    LocalMux I__2046 (
            .O(N__20539),
            .I(pwm_duty_input_3));
    Odrv4 I__2045 (
            .O(N__20536),
            .I(pwm_duty_input_3));
    LocalMux I__2044 (
            .O(N__20533),
            .I(pwm_duty_input_3));
    CascadeMux I__2043 (
            .O(N__20526),
            .I(N__20523));
    InMux I__2042 (
            .O(N__20523),
            .I(N__20520));
    LocalMux I__2041 (
            .O(N__20520),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ));
    InMux I__2040 (
            .O(N__20517),
            .I(N__20512));
    InMux I__2039 (
            .O(N__20516),
            .I(N__20509));
    InMux I__2038 (
            .O(N__20515),
            .I(N__20506));
    LocalMux I__2037 (
            .O(N__20512),
            .I(N__20503));
    LocalMux I__2036 (
            .O(N__20509),
            .I(N__20498));
    LocalMux I__2035 (
            .O(N__20506),
            .I(N__20498));
    Span4Mux_s1_h I__2034 (
            .O(N__20503),
            .I(N__20495));
    Odrv4 I__2033 (
            .O(N__20498),
            .I(pwm_duty_input_4));
    Odrv4 I__2032 (
            .O(N__20495),
            .I(pwm_duty_input_4));
    InMux I__2031 (
            .O(N__20490),
            .I(N__20487));
    LocalMux I__2030 (
            .O(N__20487),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ));
    InMux I__2029 (
            .O(N__20484),
            .I(N__20481));
    LocalMux I__2028 (
            .O(N__20481),
            .I(N__20478));
    Span4Mux_h I__2027 (
            .O(N__20478),
            .I(N__20475));
    Span4Mux_v I__2026 (
            .O(N__20475),
            .I(N__20472));
    Odrv4 I__2025 (
            .O(N__20472),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    CascadeMux I__2024 (
            .O(N__20469),
            .I(N__20466));
    InMux I__2023 (
            .O(N__20466),
            .I(N__20463));
    LocalMux I__2022 (
            .O(N__20463),
            .I(N__20460));
    Span4Mux_v I__2021 (
            .O(N__20460),
            .I(N__20457));
    Span4Mux_v I__2020 (
            .O(N__20457),
            .I(N__20454));
    Odrv4 I__2019 (
            .O(N__20454),
            .I(\pwm_generator_inst.un2_threshold_1_24 ));
    InMux I__2018 (
            .O(N__20451),
            .I(N__20448));
    LocalMux I__2017 (
            .O(N__20448),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ));
    InMux I__2016 (
            .O(N__20445),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    CascadeMux I__2015 (
            .O(N__20442),
            .I(N__20439));
    InMux I__2014 (
            .O(N__20439),
            .I(N__20436));
    LocalMux I__2013 (
            .O(N__20436),
            .I(N__20433));
    Span4Mux_h I__2012 (
            .O(N__20433),
            .I(N__20430));
    Span4Mux_v I__2011 (
            .O(N__20430),
            .I(N__20427));
    Odrv4 I__2010 (
            .O(N__20427),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__2009 (
            .O(N__20424),
            .I(N__20421));
    LocalMux I__2008 (
            .O(N__20421),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ));
    InMux I__2007 (
            .O(N__20418),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__2006 (
            .O(N__20415),
            .I(N__20412));
    InMux I__2005 (
            .O(N__20412),
            .I(N__20409));
    LocalMux I__2004 (
            .O(N__20409),
            .I(N__20406));
    Span4Mux_h I__2003 (
            .O(N__20406),
            .I(N__20403));
    Span4Mux_v I__2002 (
            .O(N__20403),
            .I(N__20400));
    Odrv4 I__2001 (
            .O(N__20400),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__2000 (
            .O(N__20397),
            .I(N__20394));
    LocalMux I__1999 (
            .O(N__20394),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ));
    InMux I__1998 (
            .O(N__20391),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    CascadeMux I__1997 (
            .O(N__20388),
            .I(N__20385));
    InMux I__1996 (
            .O(N__20385),
            .I(N__20382));
    LocalMux I__1995 (
            .O(N__20382),
            .I(N__20379));
    Span4Mux_h I__1994 (
            .O(N__20379),
            .I(N__20376));
    Span4Mux_v I__1993 (
            .O(N__20376),
            .I(N__20373));
    Odrv4 I__1992 (
            .O(N__20373),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__1991 (
            .O(N__20370),
            .I(N__20367));
    LocalMux I__1990 (
            .O(N__20367),
            .I(N__20364));
    Odrv4 I__1989 (
            .O(N__20364),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ));
    InMux I__1988 (
            .O(N__20361),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    CascadeMux I__1987 (
            .O(N__20358),
            .I(N__20355));
    InMux I__1986 (
            .O(N__20355),
            .I(N__20352));
    LocalMux I__1985 (
            .O(N__20352),
            .I(N__20349));
    Span4Mux_h I__1984 (
            .O(N__20349),
            .I(N__20346));
    Span4Mux_v I__1983 (
            .O(N__20346),
            .I(N__20343));
    Odrv4 I__1982 (
            .O(N__20343),
            .I(\pwm_generator_inst.un2_threshold_2_13 ));
    CascadeMux I__1981 (
            .O(N__20340),
            .I(N__20337));
    InMux I__1980 (
            .O(N__20337),
            .I(N__20334));
    LocalMux I__1979 (
            .O(N__20334),
            .I(N__20331));
    Odrv4 I__1978 (
            .O(N__20331),
            .I(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ));
    InMux I__1977 (
            .O(N__20328),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_12 ));
    CascadeMux I__1976 (
            .O(N__20325),
            .I(N__20322));
    InMux I__1975 (
            .O(N__20322),
            .I(N__20319));
    LocalMux I__1974 (
            .O(N__20319),
            .I(N__20316));
    Span12Mux_v I__1973 (
            .O(N__20316),
            .I(N__20313));
    Odrv12 I__1972 (
            .O(N__20313),
            .I(\pwm_generator_inst.un2_threshold_2_14 ));
    InMux I__1971 (
            .O(N__20310),
            .I(N__20307));
    LocalMux I__1970 (
            .O(N__20307),
            .I(N__20304));
    Odrv4 I__1969 (
            .O(N__20304),
            .I(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ));
    InMux I__1968 (
            .O(N__20301),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_13 ));
    InMux I__1967 (
            .O(N__20298),
            .I(N__20294));
    InMux I__1966 (
            .O(N__20297),
            .I(N__20291));
    LocalMux I__1965 (
            .O(N__20294),
            .I(N__20286));
    LocalMux I__1964 (
            .O(N__20291),
            .I(N__20286));
    Span4Mux_v I__1963 (
            .O(N__20286),
            .I(N__20277));
    InMux I__1962 (
            .O(N__20285),
            .I(N__20270));
    InMux I__1961 (
            .O(N__20284),
            .I(N__20270));
    InMux I__1960 (
            .O(N__20283),
            .I(N__20270));
    InMux I__1959 (
            .O(N__20282),
            .I(N__20263));
    InMux I__1958 (
            .O(N__20281),
            .I(N__20263));
    InMux I__1957 (
            .O(N__20280),
            .I(N__20263));
    Span4Mux_v I__1956 (
            .O(N__20277),
            .I(N__20256));
    LocalMux I__1955 (
            .O(N__20270),
            .I(N__20256));
    LocalMux I__1954 (
            .O(N__20263),
            .I(N__20256));
    Span4Mux_v I__1953 (
            .O(N__20256),
            .I(N__20253));
    Span4Mux_v I__1952 (
            .O(N__20253),
            .I(N__20250));
    Odrv4 I__1951 (
            .O(N__20250),
            .I(\pwm_generator_inst.un2_threshold_1_25 ));
    CascadeMux I__1950 (
            .O(N__20247),
            .I(N__20244));
    InMux I__1949 (
            .O(N__20244),
            .I(N__20241));
    LocalMux I__1948 (
            .O(N__20241),
            .I(N__20238));
    Span4Mux_h I__1947 (
            .O(N__20238),
            .I(N__20235));
    Span4Mux_v I__1946 (
            .O(N__20235),
            .I(N__20232));
    Odrv4 I__1945 (
            .O(N__20232),
            .I(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ));
    CascadeMux I__1944 (
            .O(N__20229),
            .I(N__20226));
    InMux I__1943 (
            .O(N__20226),
            .I(N__20223));
    LocalMux I__1942 (
            .O(N__20223),
            .I(N__20220));
    Odrv4 I__1941 (
            .O(N__20220),
            .I(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ));
    InMux I__1940 (
            .O(N__20217),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_14 ));
    InMux I__1939 (
            .O(N__20214),
            .I(N__20211));
    LocalMux I__1938 (
            .O(N__20211),
            .I(N__20208));
    Span4Mux_v I__1937 (
            .O(N__20208),
            .I(N__20205));
    Odrv4 I__1936 (
            .O(N__20205),
            .I(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ));
    InMux I__1935 (
            .O(N__20202),
            .I(N__20199));
    LocalMux I__1934 (
            .O(N__20199),
            .I(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ));
    InMux I__1933 (
            .O(N__20196),
            .I(bfn_2_17_0_));
    InMux I__1932 (
            .O(N__20193),
            .I(N__20190));
    LocalMux I__1931 (
            .O(N__20190),
            .I(N__20187));
    Span4Mux_h I__1930 (
            .O(N__20187),
            .I(N__20184));
    Span4Mux_v I__1929 (
            .O(N__20184),
            .I(N__20181));
    Odrv4 I__1928 (
            .O(N__20181),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    CascadeMux I__1927 (
            .O(N__20178),
            .I(N__20175));
    InMux I__1926 (
            .O(N__20175),
            .I(N__20172));
    LocalMux I__1925 (
            .O(N__20172),
            .I(N__20169));
    Span4Mux_v I__1924 (
            .O(N__20169),
            .I(N__20166));
    Span4Mux_v I__1923 (
            .O(N__20166),
            .I(N__20163));
    Odrv4 I__1922 (
            .O(N__20163),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    InMux I__1921 (
            .O(N__20160),
            .I(N__20157));
    LocalMux I__1920 (
            .O(N__20157),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ));
    InMux I__1919 (
            .O(N__20154),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__1918 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__1917 (
            .O(N__20148),
            .I(N__20145));
    Span4Mux_h I__1916 (
            .O(N__20145),
            .I(N__20142));
    Span4Mux_v I__1915 (
            .O(N__20142),
            .I(N__20139));
    Odrv4 I__1914 (
            .O(N__20139),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    CascadeMux I__1913 (
            .O(N__20136),
            .I(N__20133));
    InMux I__1912 (
            .O(N__20133),
            .I(N__20130));
    LocalMux I__1911 (
            .O(N__20130),
            .I(N__20127));
    Span4Mux_v I__1910 (
            .O(N__20127),
            .I(N__20124));
    Span4Mux_s3_h I__1909 (
            .O(N__20124),
            .I(N__20121));
    Span4Mux_v I__1908 (
            .O(N__20121),
            .I(N__20118));
    Odrv4 I__1907 (
            .O(N__20118),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__1906 (
            .O(N__20115),
            .I(N__20112));
    InMux I__1905 (
            .O(N__20112),
            .I(N__20109));
    LocalMux I__1904 (
            .O(N__20109),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ));
    InMux I__1903 (
            .O(N__20106),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    InMux I__1902 (
            .O(N__20103),
            .I(N__20100));
    LocalMux I__1901 (
            .O(N__20100),
            .I(N__20097));
    Span12Mux_h I__1900 (
            .O(N__20097),
            .I(N__20094));
    Odrv12 I__1899 (
            .O(N__20094),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    CascadeMux I__1898 (
            .O(N__20091),
            .I(N__20088));
    InMux I__1897 (
            .O(N__20088),
            .I(N__20085));
    LocalMux I__1896 (
            .O(N__20085),
            .I(N__20082));
    Span4Mux_v I__1895 (
            .O(N__20082),
            .I(N__20079));
    Span4Mux_v I__1894 (
            .O(N__20079),
            .I(N__20076));
    Odrv4 I__1893 (
            .O(N__20076),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    InMux I__1892 (
            .O(N__20073),
            .I(N__20070));
    LocalMux I__1891 (
            .O(N__20070),
            .I(N__20067));
    Odrv4 I__1890 (
            .O(N__20067),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ));
    InMux I__1889 (
            .O(N__20064),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__1888 (
            .O(N__20061),
            .I(N__20058));
    LocalMux I__1887 (
            .O(N__20058),
            .I(N__20055));
    Span4Mux_h I__1886 (
            .O(N__20055),
            .I(N__20052));
    Span4Mux_v I__1885 (
            .O(N__20052),
            .I(N__20049));
    Odrv4 I__1884 (
            .O(N__20049),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    CascadeMux I__1883 (
            .O(N__20046),
            .I(N__20043));
    InMux I__1882 (
            .O(N__20043),
            .I(N__20040));
    LocalMux I__1881 (
            .O(N__20040),
            .I(N__20037));
    Span4Mux_v I__1880 (
            .O(N__20037),
            .I(N__20034));
    Span4Mux_v I__1879 (
            .O(N__20034),
            .I(N__20031));
    Odrv4 I__1878 (
            .O(N__20031),
            .I(\pwm_generator_inst.un2_threshold_1_20 ));
    CascadeMux I__1877 (
            .O(N__20028),
            .I(N__20025));
    InMux I__1876 (
            .O(N__20025),
            .I(N__20022));
    LocalMux I__1875 (
            .O(N__20022),
            .I(N__20019));
    Odrv4 I__1874 (
            .O(N__20019),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ));
    InMux I__1873 (
            .O(N__20016),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__1872 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__1871 (
            .O(N__20010),
            .I(N__20007));
    Span4Mux_h I__1870 (
            .O(N__20007),
            .I(N__20004));
    Sp12to4 I__1869 (
            .O(N__20004),
            .I(N__20001));
    Odrv12 I__1868 (
            .O(N__20001),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    CascadeMux I__1867 (
            .O(N__19998),
            .I(N__19995));
    InMux I__1866 (
            .O(N__19995),
            .I(N__19992));
    LocalMux I__1865 (
            .O(N__19992),
            .I(N__19989));
    Span4Mux_v I__1864 (
            .O(N__19989),
            .I(N__19986));
    Span4Mux_v I__1863 (
            .O(N__19986),
            .I(N__19983));
    Odrv4 I__1862 (
            .O(N__19983),
            .I(\pwm_generator_inst.un2_threshold_1_21 ));
    InMux I__1861 (
            .O(N__19980),
            .I(N__19977));
    LocalMux I__1860 (
            .O(N__19977),
            .I(N__19974));
    Odrv4 I__1859 (
            .O(N__19974),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ));
    InMux I__1858 (
            .O(N__19971),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__1857 (
            .O(N__19968),
            .I(N__19965));
    LocalMux I__1856 (
            .O(N__19965),
            .I(N__19962));
    Span4Mux_s3_h I__1855 (
            .O(N__19962),
            .I(N__19959));
    Span4Mux_v I__1854 (
            .O(N__19959),
            .I(N__19956));
    Span4Mux_v I__1853 (
            .O(N__19956),
            .I(N__19953));
    Odrv4 I__1852 (
            .O(N__19953),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    CascadeMux I__1851 (
            .O(N__19950),
            .I(N__19947));
    InMux I__1850 (
            .O(N__19947),
            .I(N__19944));
    LocalMux I__1849 (
            .O(N__19944),
            .I(N__19941));
    Span4Mux_v I__1848 (
            .O(N__19941),
            .I(N__19938));
    Span4Mux_v I__1847 (
            .O(N__19938),
            .I(N__19935));
    Odrv4 I__1846 (
            .O(N__19935),
            .I(\pwm_generator_inst.un2_threshold_1_22 ));
    CascadeMux I__1845 (
            .O(N__19932),
            .I(N__19929));
    InMux I__1844 (
            .O(N__19929),
            .I(N__19926));
    LocalMux I__1843 (
            .O(N__19926),
            .I(N__19923));
    Odrv4 I__1842 (
            .O(N__19923),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ));
    InMux I__1841 (
            .O(N__19920),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__1840 (
            .O(N__19917),
            .I(N__19914));
    LocalMux I__1839 (
            .O(N__19914),
            .I(N__19911));
    Span4Mux_h I__1838 (
            .O(N__19911),
            .I(N__19908));
    Span4Mux_v I__1837 (
            .O(N__19908),
            .I(N__19905));
    Odrv4 I__1836 (
            .O(N__19905),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    CascadeMux I__1835 (
            .O(N__19902),
            .I(N__19899));
    InMux I__1834 (
            .O(N__19899),
            .I(N__19896));
    LocalMux I__1833 (
            .O(N__19896),
            .I(N__19893));
    Span4Mux_h I__1832 (
            .O(N__19893),
            .I(N__19890));
    Span4Mux_v I__1831 (
            .O(N__19890),
            .I(N__19887));
    Span4Mux_v I__1830 (
            .O(N__19887),
            .I(N__19884));
    Odrv4 I__1829 (
            .O(N__19884),
            .I(\pwm_generator_inst.un2_threshold_1_23 ));
    InMux I__1828 (
            .O(N__19881),
            .I(N__19878));
    LocalMux I__1827 (
            .O(N__19878),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ));
    InMux I__1826 (
            .O(N__19875),
            .I(bfn_2_16_0_));
    InMux I__1825 (
            .O(N__19872),
            .I(bfn_2_14_0_));
    InMux I__1824 (
            .O(N__19869),
            .I(\pwm_generator_inst.un15_threshold_1_cry_16 ));
    InMux I__1823 (
            .O(N__19866),
            .I(\pwm_generator_inst.un15_threshold_1_cry_17 ));
    InMux I__1822 (
            .O(N__19863),
            .I(\pwm_generator_inst.un15_threshold_1_cry_18 ));
    InMux I__1821 (
            .O(N__19860),
            .I(N__19857));
    LocalMux I__1820 (
            .O(N__19857),
            .I(N__19854));
    Span4Mux_h I__1819 (
            .O(N__19854),
            .I(N__19851));
    Span4Mux_v I__1818 (
            .O(N__19851),
            .I(N__19848));
    Odrv4 I__1817 (
            .O(N__19848),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__1816 (
            .O(N__19845),
            .I(N__19842));
    InMux I__1815 (
            .O(N__19842),
            .I(N__19839));
    LocalMux I__1814 (
            .O(N__19839),
            .I(N__19836));
    Span4Mux_h I__1813 (
            .O(N__19836),
            .I(N__19833));
    Span4Mux_v I__1812 (
            .O(N__19833),
            .I(N__19830));
    Span4Mux_v I__1811 (
            .O(N__19830),
            .I(N__19827));
    Odrv4 I__1810 (
            .O(N__19827),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__1809 (
            .O(N__19824),
            .I(N__19821));
    LocalMux I__1808 (
            .O(N__19821),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ));
    InMux I__1807 (
            .O(N__19818),
            .I(N__19815));
    LocalMux I__1806 (
            .O(N__19815),
            .I(N__19812));
    Span4Mux_h I__1805 (
            .O(N__19812),
            .I(N__19809));
    Span4Mux_v I__1804 (
            .O(N__19809),
            .I(N__19806));
    Odrv4 I__1803 (
            .O(N__19806),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__1802 (
            .O(N__19803),
            .I(N__19800));
    InMux I__1801 (
            .O(N__19800),
            .I(N__19797));
    LocalMux I__1800 (
            .O(N__19797),
            .I(N__19794));
    Span4Mux_v I__1799 (
            .O(N__19794),
            .I(N__19791));
    Span4Mux_v I__1798 (
            .O(N__19791),
            .I(N__19788));
    Odrv4 I__1797 (
            .O(N__19788),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    CascadeMux I__1796 (
            .O(N__19785),
            .I(N__19782));
    InMux I__1795 (
            .O(N__19782),
            .I(N__19779));
    LocalMux I__1794 (
            .O(N__19779),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ));
    InMux I__1793 (
            .O(N__19776),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__1792 (
            .O(N__19773),
            .I(N__19770));
    LocalMux I__1791 (
            .O(N__19770),
            .I(N__19767));
    Span12Mux_h I__1790 (
            .O(N__19767),
            .I(N__19764));
    Odrv12 I__1789 (
            .O(N__19764),
            .I(\pwm_generator_inst.O_7 ));
    CascadeMux I__1788 (
            .O(N__19761),
            .I(N__19758));
    InMux I__1787 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__1786 (
            .O(N__19755),
            .I(\pwm_generator_inst.un15_threshold_1_axb_7 ));
    InMux I__1785 (
            .O(N__19752),
            .I(N__19749));
    LocalMux I__1784 (
            .O(N__19749),
            .I(N__19746));
    Span4Mux_v I__1783 (
            .O(N__19746),
            .I(N__19743));
    Span4Mux_v I__1782 (
            .O(N__19743),
            .I(N__19740));
    Odrv4 I__1781 (
            .O(N__19740),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1780 (
            .O(N__19737),
            .I(N__19734));
    LocalMux I__1779 (
            .O(N__19734),
            .I(\pwm_generator_inst.un15_threshold_1_axb_8 ));
    InMux I__1778 (
            .O(N__19731),
            .I(N__19728));
    LocalMux I__1777 (
            .O(N__19728),
            .I(N__19725));
    Span4Mux_v I__1776 (
            .O(N__19725),
            .I(N__19722));
    Span4Mux_v I__1775 (
            .O(N__19722),
            .I(N__19719));
    Odrv4 I__1774 (
            .O(N__19719),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1773 (
            .O(N__19716),
            .I(N__19713));
    LocalMux I__1772 (
            .O(N__19713),
            .I(\pwm_generator_inst.un15_threshold_1_axb_9 ));
    InMux I__1771 (
            .O(N__19710),
            .I(\pwm_generator_inst.un15_threshold_1_cry_9 ));
    InMux I__1770 (
            .O(N__19707),
            .I(N__19703));
    InMux I__1769 (
            .O(N__19706),
            .I(N__19700));
    LocalMux I__1768 (
            .O(N__19703),
            .I(N__19697));
    LocalMux I__1767 (
            .O(N__19700),
            .I(N__19694));
    Span4Mux_h I__1766 (
            .O(N__19697),
            .I(N__19689));
    Span4Mux_v I__1765 (
            .O(N__19694),
            .I(N__19689));
    Span4Mux_v I__1764 (
            .O(N__19689),
            .I(N__19686));
    Odrv4 I__1763 (
            .O(N__19686),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__1762 (
            .O(N__19683),
            .I(\pwm_generator_inst.un15_threshold_1_cry_10 ));
    InMux I__1761 (
            .O(N__19680),
            .I(\pwm_generator_inst.un15_threshold_1_cry_11 ));
    InMux I__1760 (
            .O(N__19677),
            .I(\pwm_generator_inst.un15_threshold_1_cry_12 ));
    InMux I__1759 (
            .O(N__19674),
            .I(\pwm_generator_inst.un15_threshold_1_cry_13 ));
    InMux I__1758 (
            .O(N__19671),
            .I(\pwm_generator_inst.un15_threshold_1_cry_14 ));
    CascadeMux I__1757 (
            .O(N__19668),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ));
    CascadeMux I__1756 (
            .O(N__19665),
            .I(N__19662));
    InMux I__1755 (
            .O(N__19662),
            .I(N__19659));
    LocalMux I__1754 (
            .O(N__19659),
            .I(N__19655));
    InMux I__1753 (
            .O(N__19658),
            .I(N__19652));
    Odrv4 I__1752 (
            .O(N__19655),
            .I(\current_shift_inst.PI_CTRL.N_306 ));
    LocalMux I__1751 (
            .O(N__19652),
            .I(\current_shift_inst.PI_CTRL.N_306 ));
    InMux I__1750 (
            .O(N__19647),
            .I(N__19644));
    LocalMux I__1749 (
            .O(N__19644),
            .I(N__19641));
    Span4Mux_v I__1748 (
            .O(N__19641),
            .I(N__19638));
    Span4Mux_v I__1747 (
            .O(N__19638),
            .I(N__19635));
    Odrv4 I__1746 (
            .O(N__19635),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1745 (
            .O(N__19632),
            .I(N__19629));
    LocalMux I__1744 (
            .O(N__19629),
            .I(\pwm_generator_inst.un15_threshold_1_axb_0 ));
    InMux I__1743 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__1742 (
            .O(N__19623),
            .I(N__19620));
    Span4Mux_v I__1741 (
            .O(N__19620),
            .I(N__19617));
    Span4Mux_v I__1740 (
            .O(N__19617),
            .I(N__19614));
    Odrv4 I__1739 (
            .O(N__19614),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1738 (
            .O(N__19611),
            .I(N__19608));
    LocalMux I__1737 (
            .O(N__19608),
            .I(\pwm_generator_inst.un15_threshold_1_axb_1 ));
    InMux I__1736 (
            .O(N__19605),
            .I(N__19602));
    LocalMux I__1735 (
            .O(N__19602),
            .I(N__19599));
    Span4Mux_h I__1734 (
            .O(N__19599),
            .I(N__19596));
    Span4Mux_v I__1733 (
            .O(N__19596),
            .I(N__19593));
    Odrv4 I__1732 (
            .O(N__19593),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1731 (
            .O(N__19590),
            .I(N__19587));
    LocalMux I__1730 (
            .O(N__19587),
            .I(\pwm_generator_inst.un15_threshold_1_axb_2 ));
    InMux I__1729 (
            .O(N__19584),
            .I(N__19581));
    LocalMux I__1728 (
            .O(N__19581),
            .I(N__19578));
    Span4Mux_h I__1727 (
            .O(N__19578),
            .I(N__19575));
    Span4Mux_v I__1726 (
            .O(N__19575),
            .I(N__19572));
    Odrv4 I__1725 (
            .O(N__19572),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1724 (
            .O(N__19569),
            .I(N__19566));
    LocalMux I__1723 (
            .O(N__19566),
            .I(\pwm_generator_inst.un15_threshold_1_axb_3 ));
    InMux I__1722 (
            .O(N__19563),
            .I(N__19560));
    LocalMux I__1721 (
            .O(N__19560),
            .I(N__19557));
    Span4Mux_h I__1720 (
            .O(N__19557),
            .I(N__19554));
    Span4Mux_v I__1719 (
            .O(N__19554),
            .I(N__19551));
    Odrv4 I__1718 (
            .O(N__19551),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1717 (
            .O(N__19548),
            .I(N__19545));
    LocalMux I__1716 (
            .O(N__19545),
            .I(\pwm_generator_inst.un15_threshold_1_axb_4 ));
    InMux I__1715 (
            .O(N__19542),
            .I(N__19539));
    LocalMux I__1714 (
            .O(N__19539),
            .I(N__19536));
    Span4Mux_h I__1713 (
            .O(N__19536),
            .I(N__19533));
    Span4Mux_v I__1712 (
            .O(N__19533),
            .I(N__19530));
    Odrv4 I__1711 (
            .O(N__19530),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1710 (
            .O(N__19527),
            .I(N__19524));
    LocalMux I__1709 (
            .O(N__19524),
            .I(\pwm_generator_inst.un15_threshold_1_axb_5 ));
    InMux I__1708 (
            .O(N__19521),
            .I(N__19518));
    LocalMux I__1707 (
            .O(N__19518),
            .I(N__19515));
    Span12Mux_v I__1706 (
            .O(N__19515),
            .I(N__19512));
    Odrv12 I__1705 (
            .O(N__19512),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1704 (
            .O(N__19509),
            .I(N__19506));
    LocalMux I__1703 (
            .O(N__19506),
            .I(\pwm_generator_inst.un15_threshold_1_axb_6 ));
    CascadeMux I__1702 (
            .O(N__19503),
            .I(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ));
    InMux I__1701 (
            .O(N__19500),
            .I(N__19493));
    InMux I__1700 (
            .O(N__19499),
            .I(N__19493));
    InMux I__1699 (
            .O(N__19498),
            .I(N__19490));
    LocalMux I__1698 (
            .O(N__19493),
            .I(pwm_duty_input_8));
    LocalMux I__1697 (
            .O(N__19490),
            .I(pwm_duty_input_8));
    InMux I__1696 (
            .O(N__19485),
            .I(N__19478));
    InMux I__1695 (
            .O(N__19484),
            .I(N__19478));
    InMux I__1694 (
            .O(N__19483),
            .I(N__19475));
    LocalMux I__1693 (
            .O(N__19478),
            .I(N__19472));
    LocalMux I__1692 (
            .O(N__19475),
            .I(N__19469));
    Odrv4 I__1691 (
            .O(N__19472),
            .I(pwm_duty_input_9));
    Odrv4 I__1690 (
            .O(N__19469),
            .I(pwm_duty_input_9));
    CascadeMux I__1689 (
            .O(N__19464),
            .I(N__19460));
    InMux I__1688 (
            .O(N__19463),
            .I(N__19456));
    InMux I__1687 (
            .O(N__19460),
            .I(N__19451));
    InMux I__1686 (
            .O(N__19459),
            .I(N__19451));
    LocalMux I__1685 (
            .O(N__19456),
            .I(N__19448));
    LocalMux I__1684 (
            .O(N__19451),
            .I(pwm_duty_input_7));
    Odrv4 I__1683 (
            .O(N__19448),
            .I(pwm_duty_input_7));
    InMux I__1682 (
            .O(N__19443),
            .I(N__19436));
    InMux I__1681 (
            .O(N__19442),
            .I(N__19436));
    InMux I__1680 (
            .O(N__19441),
            .I(N__19433));
    LocalMux I__1679 (
            .O(N__19436),
            .I(pwm_duty_input_6));
    LocalMux I__1678 (
            .O(N__19433),
            .I(pwm_duty_input_6));
    CascadeMux I__1677 (
            .O(N__19428),
            .I(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ));
    InMux I__1676 (
            .O(N__19425),
            .I(N__19422));
    LocalMux I__1675 (
            .O(N__19422),
            .I(N__19417));
    InMux I__1674 (
            .O(N__19421),
            .I(N__19412));
    InMux I__1673 (
            .O(N__19420),
            .I(N__19412));
    Span4Mux_v I__1672 (
            .O(N__19417),
            .I(N__19409));
    LocalMux I__1671 (
            .O(N__19412),
            .I(pwm_duty_input_5));
    Odrv4 I__1670 (
            .O(N__19409),
            .I(pwm_duty_input_5));
    InMux I__1669 (
            .O(N__19404),
            .I(N__19400));
    InMux I__1668 (
            .O(N__19403),
            .I(N__19397));
    LocalMux I__1667 (
            .O(N__19400),
            .I(N__19392));
    LocalMux I__1666 (
            .O(N__19397),
            .I(N__19392));
    Odrv4 I__1665 (
            .O(N__19392),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__1664 (
            .O(N__19389),
            .I(N__19380));
    InMux I__1663 (
            .O(N__19388),
            .I(N__19380));
    InMux I__1662 (
            .O(N__19387),
            .I(N__19380));
    LocalMux I__1661 (
            .O(N__19380),
            .I(\current_shift_inst.PI_CTRL.N_120 ));
    CascadeMux I__1660 (
            .O(N__19377),
            .I(\current_shift_inst.PI_CTRL.N_31_cascade_ ));
    InMux I__1659 (
            .O(N__19374),
            .I(N__19370));
    InMux I__1658 (
            .O(N__19373),
            .I(N__19367));
    LocalMux I__1657 (
            .O(N__19370),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__1656 (
            .O(N__19367),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__1655 (
            .O(N__19362),
            .I(N__19358));
    InMux I__1654 (
            .O(N__19361),
            .I(N__19355));
    LocalMux I__1653 (
            .O(N__19358),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    LocalMux I__1652 (
            .O(N__19355),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    CascadeMux I__1651 (
            .O(N__19350),
            .I(N__19347));
    InMux I__1650 (
            .O(N__19347),
            .I(N__19344));
    LocalMux I__1649 (
            .O(N__19344),
            .I(\current_shift_inst.PI_CTRL.N_97 ));
    InMux I__1648 (
            .O(N__19341),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__1647 (
            .O(N__19338),
            .I(N__19334));
    InMux I__1646 (
            .O(N__19337),
            .I(N__19331));
    LocalMux I__1645 (
            .O(N__19334),
            .I(N__19328));
    LocalMux I__1644 (
            .O(N__19331),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    Odrv4 I__1643 (
            .O(N__19328),
            .I(\pwm_generator_inst.un2_threshold_2_1_15 ));
    InMux I__1642 (
            .O(N__19323),
            .I(N__19320));
    LocalMux I__1641 (
            .O(N__19320),
            .I(N__19317));
    Odrv4 I__1640 (
            .O(N__19317),
            .I(\pwm_generator_inst.un2_threshold_2_1_16 ));
    InMux I__1639 (
            .O(N__19314),
            .I(N__19311));
    LocalMux I__1638 (
            .O(N__19311),
            .I(N_6_0));
    InMux I__1637 (
            .O(N__19308),
            .I(N__19305));
    LocalMux I__1636 (
            .O(N__19305),
            .I(m38));
    InMux I__1635 (
            .O(N__19302),
            .I(N__19298));
    InMux I__1634 (
            .O(N__19301),
            .I(N__19295));
    LocalMux I__1633 (
            .O(N__19298),
            .I(N__19292));
    LocalMux I__1632 (
            .O(N__19295),
            .I(pwm_duty_input_0));
    Odrv4 I__1631 (
            .O(N__19292),
            .I(pwm_duty_input_0));
    InMux I__1630 (
            .O(N__19287),
            .I(N__19283));
    InMux I__1629 (
            .O(N__19286),
            .I(N__19280));
    LocalMux I__1628 (
            .O(N__19283),
            .I(N__19277));
    LocalMux I__1627 (
            .O(N__19280),
            .I(pwm_duty_input_1));
    Odrv4 I__1626 (
            .O(N__19277),
            .I(pwm_duty_input_1));
    InMux I__1625 (
            .O(N__19272),
            .I(N__19268));
    InMux I__1624 (
            .O(N__19271),
            .I(N__19265));
    LocalMux I__1623 (
            .O(N__19268),
            .I(N__19262));
    LocalMux I__1622 (
            .O(N__19265),
            .I(pwm_duty_input_2));
    Odrv4 I__1621 (
            .O(N__19262),
            .I(pwm_duty_input_2));
    InMux I__1620 (
            .O(N__19257),
            .I(N__19254));
    LocalMux I__1619 (
            .O(N__19254),
            .I(N__19251));
    Span4Mux_v I__1618 (
            .O(N__19251),
            .I(N__19248));
    Span4Mux_v I__1617 (
            .O(N__19248),
            .I(N__19245));
    Odrv4 I__1616 (
            .O(N__19245),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1615 (
            .O(N__19242),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    InMux I__1614 (
            .O(N__19239),
            .I(N__19236));
    LocalMux I__1613 (
            .O(N__19236),
            .I(N__19233));
    Span4Mux_v I__1612 (
            .O(N__19233),
            .I(N__19230));
    Span4Mux_v I__1611 (
            .O(N__19230),
            .I(N__19227));
    Odrv4 I__1610 (
            .O(N__19227),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1609 (
            .O(N__19224),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__1608 (
            .O(N__19221),
            .I(N__19218));
    LocalMux I__1607 (
            .O(N__19218),
            .I(N__19215));
    Span4Mux_v I__1606 (
            .O(N__19215),
            .I(N__19212));
    Span4Mux_v I__1605 (
            .O(N__19212),
            .I(N__19209));
    Odrv4 I__1604 (
            .O(N__19209),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1603 (
            .O(N__19206),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__1602 (
            .O(N__19203),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__1601 (
            .O(N__19200),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__1600 (
            .O(N__19197),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__1599 (
            .O(N__19194),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    InMux I__1598 (
            .O(N__19191),
            .I(bfn_1_17_0_));
    InMux I__1597 (
            .O(N__19188),
            .I(N__19185));
    LocalMux I__1596 (
            .O(N__19185),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__1595 (
            .O(N__19182),
            .I(\current_shift_inst.PI_CTRL.N_98_cascade_ ));
    InMux I__1594 (
            .O(N__19179),
            .I(N__19176));
    LocalMux I__1593 (
            .O(N__19176),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    IoInMux I__1592 (
            .O(N__19173),
            .I(N__19170));
    LocalMux I__1591 (
            .O(N__19170),
            .I(N__19167));
    IoSpan4Mux I__1590 (
            .O(N__19167),
            .I(N__19164));
    IoSpan4Mux I__1589 (
            .O(N__19164),
            .I(N__19161));
    Odrv4 I__1588 (
            .O(N__19161),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    IoInMux I__1587 (
            .O(N__19158),
            .I(N__19155));
    LocalMux I__1586 (
            .O(N__19155),
            .I(N__19152));
    Span4Mux_s3_v I__1585 (
            .O(N__19152),
            .I(N__19149));
    Span4Mux_h I__1584 (
            .O(N__19149),
            .I(N__19146));
    Sp12to4 I__1583 (
            .O(N__19146),
            .I(N__19143));
    Span12Mux_v I__1582 (
            .O(N__19143),
            .I(N__19140));
    Span12Mux_v I__1581 (
            .O(N__19140),
            .I(N__19137));
    Odrv12 I__1580 (
            .O(N__19137),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_1_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_18_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_1_18_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_17_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_17_22_0_));
    defparam IN_MUX_bfv_17_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_23_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_17_23_0_));
    defparam IN_MUX_bfv_5_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_15_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_5_16_0_));
    defparam IN_MUX_bfv_5_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_17_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_5_17_0_));
    defparam IN_MUX_bfv_5_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_5_18_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_3_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_15_0_));
    defparam IN_MUX_bfv_3_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_16_0_ (
            .carryinitin(\pwm_generator_inst.un19_threshold_cry_7 ),
            .carryinitout(bfn_3_16_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .carryinitout(bfn_2_13_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_13_0_));
    defparam IN_MUX_bfv_4_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_14_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_4_14_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_3_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_19_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_3_19_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_12_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_8_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_17_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_16_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_17_16_0_));
    defparam IN_MUX_bfv_17_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_17_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_17_17_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_16_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_6_0_));
    defparam IN_MUX_bfv_16_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .carryinitout(bfn_16_7_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_16_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_16_17_0_));
    defparam IN_MUX_bfv_18_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_22_0_));
    defparam IN_MUX_bfv_18_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_23_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_18_23_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_14_21_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19158),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19173),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \phase_controller_inst2.stoper_tr.un1_start_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__29912),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un1_start_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNI8ENL_0  (
            .USERSIGNALTOGLOBALBUFFER(N__38658),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_339_i_g ));
    ICE_GB \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0  (
            .USERSIGNALTOGLOBALBUFFER(N__47166),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_hc.un1_start_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__49882),
            .CLKHFEN(N__49884),
            .CLKHF(clk_12mhz));
    defparam rgb_drv.RGB2_CURRENT="0b111111";
    defparam rgb_drv.CURRENT_MODE="0b0";
    defparam rgb_drv.RGB0_CURRENT="0b111111";
    defparam rgb_drv.RGB1_CURRENT="0b111111";
    SB_RGBA_DRV rgb_drv (
            .RGBLEDEN(N__49883),
            .RGB2PWM(N__19314),
            .RGB1(rgb_g),
            .CURREN(N__49814),
            .RGB2(rgb_b),
            .RGB1PWM(N__19308),
            .RGB0PWM(N__50418),
            .RGB0(rgb_r));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_4_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_4_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_1_4_4 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_1_4_4  (
            .in0(N__23055),
            .in1(N__22281),
            .in2(N__22420),
            .in3(N__21018),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50915),
            .ce(),
            .sr(N__50338));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_5_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_5_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21315),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50914),
            .ce(),
            .sr(N__50345));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_1_5_2  (
            .in0(N__19388),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21897),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50914),
            .ce(),
            .sr(N__50345));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_1_5_4  (
            .in0(N__19389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22227),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50914),
            .ce(),
            .sr(N__50345));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__19179),
            .in2(_gnd_net_),
            .in3(N__19387),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50914),
            .ce(),
            .sr(N__50345));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_6_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_1_6_0 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_1_6_0  (
            .in0(N__21016),
            .in1(N__23036),
            .in2(N__22284),
            .in3(N__22452),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50913),
            .ce(),
            .sr(N__50352));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_1 .LUT_INIT=16'b0010001100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_1_6_1  (
            .in0(N__22164),
            .in1(N__19188),
            .in2(N__19665),
            .in3(N__22280),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50913),
            .ce(),
            .sr(N__50352));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_1_6_2  (
            .in0(N__21015),
            .in1(N__23035),
            .in2(N__22283),
            .in3(N__22494),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50913),
            .ce(),
            .sr(N__50352));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_6_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_6_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_1_6_5 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_1_6_5  (
            .in0(N__23033),
            .in1(N__22279),
            .in2(N__22584),
            .in3(N__21017),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50913),
            .ce(),
            .sr(N__50352));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_6 .LUT_INIT=16'b1111001100100010;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_1_6_6  (
            .in0(N__21014),
            .in1(N__23034),
            .in2(N__22282),
            .in3(N__22541),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50913),
            .ce(),
            .sr(N__50352));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_7 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_1_6_7  (
            .in0(N__22209),
            .in1(N__19404),
            .in2(_gnd_net_),
            .in3(N__19374),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50913),
            .ce(),
            .sr(N__50352));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_7_1 .LUT_INIT=16'b0000111100000111;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_1_7_1  (
            .in0(N__22167),
            .in1(N__19362),
            .in2(N__23054),
            .in3(N__21010),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_8_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_1_8_0  (
            .in0(_gnd_net_),
            .in1(N__22165),
            .in2(_gnd_net_),
            .in3(N__22201),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_8_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_8_1 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_1_8_1  (
            .in0(N__23037),
            .in1(N__19658),
            .in2(N__19182),
            .in3(N__22255),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_1_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23053),
            .lcout(N_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50905),
            .ce(),
            .sr(N__50374));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_12_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(N__21206),
            .in2(_gnd_net_),
            .in3(N__21170),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_1_15_1  (
            .in0(N__21253),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21227),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_1_15_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_1_15_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__20621),
            .in2(_gnd_net_),
            .in3(N__20642),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_1_15_3  (
            .in0(N__20665),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20681),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_1_15_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_1_15_5 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__20588),
            .in2(_gnd_net_),
            .in3(N__20573),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__19706),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__19257),
            .in2(_gnd_net_),
            .in3(N__19242),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__19239),
            .in2(_gnd_net_),
            .in3(N__19224),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__19221),
            .in2(_gnd_net_),
            .in3(N__19206),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__19824),
            .in2(_gnd_net_),
            .in3(N__19203),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__49785),
            .in2(N__19785),
            .in3(N__19200),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(N__20160),
            .in2(N__49815),
            .in3(N__19197),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(N__49789),
            .in2(N__20115),
            .in3(N__19194),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__20073),
            .in2(_gnd_net_),
            .in3(N__19191),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20028),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_LC_1_17_2  (
            .in0(_gnd_net_),
            .in1(N__19980),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__19881),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(N__20451),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__20424),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(N__20397),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(N__20370),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_18_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20340),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__20310),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_18_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_LC_1_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20229),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_18_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_1_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19341),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_22_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_1_22_4  (
            .in0(N__19338),
            .in1(N__20298),
            .in2(_gnd_net_),
            .in3(N__21558),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_23_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_23_2 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_1_23_2  (
            .in0(N__19337),
            .in1(N__20297),
            .in2(N__21603),
            .in3(N__19323),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.m5_LC_1_30_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m5_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m5_LC_1_30_1 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \phase_controller_inst1.stoper_hc.m5_LC_1_30_1  (
            .in0(N__50417),
            .in1(N__43689),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.m38_LC_1_30_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m38_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m38_LC_1_30_3 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.m38_LC_1_30_3  (
            .in0(N__50416),
            .in1(N__43688),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(m38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pwm_generator_inst.un1_duty_inputlto2_LC_2_5_6  (
            .in0(N__19301),
            .in1(N__19286),
            .in2(_gnd_net_),
            .in3(N__19271),
            .lcout(\pwm_generator_inst.un1_duty_inputlt3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_4_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__19459),
            .in2(_gnd_net_),
            .in3(N__19420),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_3_LC_2_6_2  (
            .in0(N__19499),
            .in1(N__19484),
            .in2(N__19503),
            .in3(N__19442),
            .lcout(\pwm_generator_inst.un2_duty_input_0_o3Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_6_4  (
            .in0(N__19500),
            .in1(N__19485),
            .in2(N__19464),
            .in3(N__19443),
            .lcout(),
            .ltout(\pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_5 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_6_5  (
            .in0(N__20546),
            .in1(N__20516),
            .in2(N__19428),
            .in3(N__19421),
            .lcout(\pwm_generator_inst.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_6_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_6_6 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_6_6  (
            .in0(N__19373),
            .in1(N__19403),
            .in2(N__19350),
            .in3(N__22208),
            .lcout(\current_shift_inst.PI_CTRL.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_7_0  (
            .in0(N__22489),
            .in1(N__22447),
            .in2(N__22542),
            .in3(N__20490),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(\current_shift_inst.PI_CTRL.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_7_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_7_1 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_7_1  (
            .in0(N__20993),
            .in1(N__23032),
            .in2(N__19377),
            .in3(N__22166),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_7_4  (
            .in0(N__23031),
            .in1(N__20994),
            .in2(_gnd_net_),
            .in3(N__19361),
            .lcout(\current_shift_inst.PI_CTRL.N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_8_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_8_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__22531),
            .in2(_gnd_net_),
            .in3(N__22422),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_8_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_2_8_4  (
            .in0(N__22448),
            .in1(N__22490),
            .in2(N__19668),
            .in3(N__22577),
            .lcout(\current_shift_inst.PI_CTRL.N_306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_12_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(N__19632),
            .in2(_gnd_net_),
            .in3(N__19647),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_12_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__19611),
            .in2(_gnd_net_),
            .in3(N__19626),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_12_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(N__19590),
            .in2(_gnd_net_),
            .in3(N__19605),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_12_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__19569),
            .in2(_gnd_net_),
            .in3(N__19584),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_12_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__19548),
            .in2(_gnd_net_),
            .in3(N__19563),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_12_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(N__19527),
            .in2(_gnd_net_),
            .in3(N__19542),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_12_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__19509),
            .in2(_gnd_net_),
            .in3(N__19521),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_12_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_12_7  (
            .in0(N__19773),
            .in1(_gnd_net_),
            .in2(N__19761),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__19737),
            .in2(_gnd_net_),
            .in3(N__19752),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__19716),
            .in2(_gnd_net_),
            .in3(N__19731),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(N__21202),
            .in2(_gnd_net_),
            .in3(N__19710),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_13_3 .LUT_INIT=16'b1001100100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_13_3  (
            .in0(N__21113),
            .in1(N__19707),
            .in2(_gnd_net_),
            .in3(N__19683),
            .lcout(\pwm_generator_inst.un19_threshold_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__21040),
            .in2(_gnd_net_),
            .in3(N__19680),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__21254),
            .in2(_gnd_net_),
            .in3(N__19677),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_13_6  (
            .in0(_gnd_net_),
            .in1(N__20666),
            .in2(_gnd_net_),
            .in3(N__19674),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(N__20779),
            .in2(_gnd_net_),
            .in3(N__19671),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__20836),
            .in2(_gnd_net_),
            .in3(N__19872),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__20569),
            .in2(_gnd_net_),
            .in3(N__19869),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__20641),
            .in2(_gnd_net_),
            .in3(N__19866),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un15_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un15_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_14_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19863),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_14_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(N__20837),
            .in2(_gnd_net_),
            .in3(N__20822),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_14_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_2_14_6  (
            .in0(N__21131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21044),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_14_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_14_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(N__20762),
            .in2(_gnd_net_),
            .in3(N__20783),
            .lcout(\pwm_generator_inst.un15_threshold_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_2_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_4_LC_2_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_4_LC_2_15_0  (
            .in0(_gnd_net_),
            .in1(N__19860),
            .in2(N__19845),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_4 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_2_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_2_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(N__19818),
            .in2(N__19803),
            .in3(N__19776),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_2_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_2_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_2_15_2  (
            .in0(_gnd_net_),
            .in1(N__20193),
            .in2(N__20178),
            .in3(N__20154),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_2_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_2_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__20151),
            .in2(N__20136),
            .in3(N__20106),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_2_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_2_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(N__20103),
            .in2(N__20091),
            .in3(N__20064),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_2_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_2_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_2_15_5  (
            .in0(_gnd_net_),
            .in1(N__20061),
            .in2(N__20046),
            .in3(N__20016),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_2_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_2_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__20013),
            .in2(N__19998),
            .in3(N__19971),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_2_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_2_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(N__19968),
            .in2(N__19950),
            .in3(N__19920),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_2_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_2_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__19917),
            .in2(N__19902),
            .in3(N__19875),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(bfn_2_16_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_2_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_2_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_2_16_1  (
            .in0(_gnd_net_),
            .in1(N__20484),
            .in2(N__20469),
            .in3(N__20445),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_2_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_2_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_2_16_2  (
            .in0(_gnd_net_),
            .in1(N__20280),
            .in2(N__20442),
            .in3(N__20418),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_2_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_2_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_2_16_3  (
            .in0(_gnd_net_),
            .in1(N__20283),
            .in2(N__20415),
            .in3(N__20391),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_2_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_2_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_2_16_4  (
            .in0(_gnd_net_),
            .in1(N__20281),
            .in2(N__20388),
            .in3(N__20361),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_2_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_2_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_2_16_5  (
            .in0(_gnd_net_),
            .in1(N__20284),
            .in2(N__20358),
            .in3(N__20328),
            .lcout(\pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_2_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_2_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_2_16_6  (
            .in0(_gnd_net_),
            .in1(N__20282),
            .in2(N__20325),
            .in3(N__20301),
            .lcout(\pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_2_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_2_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_2_16_7  (
            .in0(_gnd_net_),
            .in1(N__20285),
            .in2(N__20247),
            .in3(N__20217),
            .lcout(\pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_2_17_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_2_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_2_17_0  (
            .in0(N__20214),
            .in1(N__20202),
            .in2(_gnd_net_),
            .in3(N__20196),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_17_2 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_2_17_2  (
            .in0(N__20691),
            .in1(N__20682),
            .in2(N__20670),
            .in3(N__21097),
            .lcout(\pwm_generator_inst.un19_threshold_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_17_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_17_4 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_2_17_4  (
            .in0(N__20643),
            .in1(N__20622),
            .in2(N__20610),
            .in3(N__21099),
            .lcout(\pwm_generator_inst.un19_threshold_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_17_6 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_2_17_6  (
            .in0(N__20598),
            .in1(N__20589),
            .in2(N__20577),
            .in3(N__21098),
            .lcout(\pwm_generator_inst.un19_threshold_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_5 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \pwm_generator_inst.un2_duty_input_0_o3_LC_3_6_5  (
            .in0(N__20553),
            .in1(N__20547),
            .in2(N__20526),
            .in3(N__20515),
            .lcout(\pwm_generator_inst.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_7_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_7_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_3_7_2  (
            .in0(_gnd_net_),
            .in1(N__22421),
            .in2(_gnd_net_),
            .in3(N__22570),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_3_14_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_3_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_3_14_0 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_3_14_0  (
            .in0(N__21700),
            .in1(N__21652),
            .in2(N__21605),
            .in3(N__20700),
            .lcout(\pwm_generator_inst.threshold_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_3_14_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_3_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_3_14_1 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_3_14_1  (
            .in0(N__21651),
            .in1(N__21574),
            .in2(N__20712),
            .in3(N__21699),
            .lcout(\pwm_generator_inst.threshold_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_3_14_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_3_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_3_14_2 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_3_14_2  (
            .in0(N__21698),
            .in1(N__20721),
            .in2(N__21604),
            .in3(N__21650),
            .lcout(\pwm_generator_inst.un14_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_3_14_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_3_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_3_14_3 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_3_14_3  (
            .in0(N__21656),
            .in1(N__21582),
            .in2(N__20898),
            .in3(N__21704),
            .lcout(\pwm_generator_inst.un14_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_3_14_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_3_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_3_14_4 .LUT_INIT=16'b1111111101010011;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_3_14_4  (
            .in0(N__21703),
            .in1(N__21655),
            .in2(N__21607),
            .in3(N__20916),
            .lcout(\pwm_generator_inst.un14_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_3_14_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_3_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_3_14_5 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_3_14_5  (
            .in0(N__21653),
            .in1(N__21578),
            .in2(N__20937),
            .in3(N__21701),
            .lcout(\pwm_generator_inst.threshold_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_3_14_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_3_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_3_14_6 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_3_14_6  (
            .in0(N__21702),
            .in1(N__21654),
            .in2(N__21606),
            .in3(N__20925),
            .lcout(\pwm_generator_inst.threshold_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_3_14_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_3_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_3_14_7 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_3_14_7  (
            .in0(N__21649),
            .in1(N__21570),
            .in2(N__20739),
            .in3(N__21697),
            .lcout(\pwm_generator_inst.threshold_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_15_0  (
            .in0(_gnd_net_),
            .in1(N__21147),
            .in2(N__21114),
            .in3(N__21110),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93 ),
            .ltout(),
            .carryin(bfn_3_15_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_15_1  (
            .in0(_gnd_net_),
            .in1(N__20730),
            .in2(_gnd_net_),
            .in3(N__20715),
            .lcout(\pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_15_2  (
            .in0(_gnd_net_),
            .in1(N__21024),
            .in2(_gnd_net_),
            .in3(N__20703),
            .lcout(\pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_15_3  (
            .in0(_gnd_net_),
            .in1(N__21216),
            .in2(_gnd_net_),
            .in3(N__20694),
            .lcout(\pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_15_4  (
            .in0(_gnd_net_),
            .in1(N__20946),
            .in2(_gnd_net_),
            .in3(N__20928),
            .lcout(\pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_15_5  (
            .in0(_gnd_net_),
            .in1(N__20745),
            .in2(_gnd_net_),
            .in3(N__20919),
            .lcout(\pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_15_6  (
            .in0(_gnd_net_),
            .in1(N__20805),
            .in2(_gnd_net_),
            .in3(N__20910),
            .lcout(\pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_15_7  (
            .in0(_gnd_net_),
            .in1(N__20907),
            .in2(_gnd_net_),
            .in3(N__20889),
            .lcout(\pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un19_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un19_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_16_0  (
            .in0(_gnd_net_),
            .in1(N__20886),
            .in2(_gnd_net_),
            .in3(N__20880),
            .lcout(\pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033 ),
            .ltout(),
            .carryin(bfn_3_16_0_),
            .carryout(\pwm_generator_inst.un19_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_16_1 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_16_1  (
            .in0(N__20877),
            .in1(N__21103),
            .in2(N__20865),
            .in3(N__20853),
            .lcout(\pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_16_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_16_2 .LUT_INIT=16'b1001111110010000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_16_2  (
            .in0(N__20850),
            .in1(N__20841),
            .in2(N__21112),
            .in3(N__20823),
            .lcout(\pwm_generator_inst.un19_threshold_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_16_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_16_3 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_16_3  (
            .in0(N__21096),
            .in1(N__20799),
            .in2(N__20790),
            .in3(N__20763),
            .lcout(\pwm_generator_inst.un19_threshold_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_16_4 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_3_16_4  (
            .in0(N__21267),
            .in1(N__21258),
            .in2(N__21234),
            .in3(N__21095),
            .lcout(\pwm_generator_inst.un19_threshold_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_3_16_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_3_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_3_16_6 .LUT_INIT=16'b1001100111110000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_3_16_6  (
            .in0(N__21210),
            .in1(N__21186),
            .in2(N__21177),
            .in3(N__21091),
            .lcout(\pwm_generator_inst.un19_threshold_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_16_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_16_7 .LUT_INIT=16'b1010110001011100;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_3_16_7  (
            .in0(N__21141),
            .in1(N__21132),
            .in2(N__21111),
            .in3(N__21045),
            .lcout(\pwm_generator_inst.un19_threshold_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_3_17_1  (
            .in0(N__21435),
            .in1(N__21852),
            .in2(N__21873),
            .in3(N__21861),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_3_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_3_18_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_3_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_3_18_0  (
            .in0(N__21933),
            .in1(N__22088),
            .in2(_gnd_net_),
            .in3(N__20961),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_1_LC_3_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_3_18_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_3_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_3_18_1  (
            .in0(N__21927),
            .in1(N__22013),
            .in2(_gnd_net_),
            .in3(N__20958),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_2_LC_3_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_3_18_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_3_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_3_18_2  (
            .in0(N__21934),
            .in1(N__22112),
            .in2(_gnd_net_),
            .in3(N__20955),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_3_LC_3_18_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_3_18_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_3_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_3_18_3  (
            .in0(N__21928),
            .in1(N__22040),
            .in2(_gnd_net_),
            .in3(N__20952),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_4_LC_3_18_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_3_18_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_3_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_3_18_4  (
            .in0(N__21935),
            .in1(N__22064),
            .in2(_gnd_net_),
            .in3(N__20949),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_5_LC_3_18_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_3_18_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_3_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_3_18_5  (
            .in0(N__21929),
            .in1(N__21955),
            .in2(_gnd_net_),
            .in3(N__21330),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_6_LC_3_18_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_3_18_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_3_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_3_18_6  (
            .in0(N__21936),
            .in1(N__21983),
            .in2(_gnd_net_),
            .in3(N__21327),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_7_LC_3_18_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_3_18_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_3_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_3_18_7  (
            .in0(N__21930),
            .in1(N__21779),
            .in2(_gnd_net_),
            .in3(N__21324),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__50821),
            .ce(),
            .sr(N__50389));
    defparam \pwm_generator_inst.counter_8_LC_3_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_3_19_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_3_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_3_19_0  (
            .in0(N__21932),
            .in1(N__21803),
            .in2(_gnd_net_),
            .in3(N__21321),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_3_19_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__50811),
            .ce(),
            .sr(N__50393));
    defparam \pwm_generator_inst.counter_9_LC_3_19_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_3_19_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_3_19_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_3_19_1  (
            .in0(N__21827),
            .in1(N__21931),
            .in2(_gnd_net_),
            .in3(N__21318),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50811),
            .ce(),
            .sr(N__50393));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_4_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_4_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_4_10_6 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_4_10_6  (
            .in0(N__22329),
            .in1(N__31311),
            .in2(_gnd_net_),
            .in3(N__28628),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50894),
            .ce(),
            .sr(N__50358));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30696),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50877),
            .ce(),
            .sr(N__50369));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_13_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_4_13_0  (
            .in0(_gnd_net_),
            .in1(N__21288),
            .in2(N__21300),
            .in3(N__22092),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_4_13_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_13_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__21273),
            .in2(N__21282),
            .in3(N__22017),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_13_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__21420),
            .in2(N__21429),
            .in3(N__22116),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_13_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__21402),
            .in2(N__21414),
            .in3(N__22044),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_13_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__21387),
            .in2(N__21396),
            .in3(N__22068),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_13_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(N__21372),
            .in2(N__21381),
            .in3(N__21960),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_13_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__21357),
            .in2(N__21366),
            .in3(N__21987),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_13_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(N__21351),
            .in2(N__21345),
            .in3(N__21783),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_4_14_0  (
            .in0(_gnd_net_),
            .in1(N__21336),
            .in2(N__21720),
            .in3(N__21807),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_4_14_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__21759),
            .in2(N__21444),
            .in3(N__21831),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_4_14_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_4_14_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_4_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_4_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21753),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50854),
            .ce(),
            .sr(N__50375));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_4_15_1  (
            .in0(N__22815),
            .in1(N__22677),
            .in2(N__22659),
            .in3(N__23076),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_15_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(N__22343),
            .in2(_gnd_net_),
            .in3(N__22377),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_4_15_3  (
            .in0(N__22362),
            .in1(N__22794),
            .in2(N__21732),
            .in3(N__21840),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_15_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_15_6 .LUT_INIT=16'b1111000111111101;
    LogicCell40 \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_4_15_6  (
            .in0(N__21662),
            .in1(N__21611),
            .in2(N__21729),
            .in3(N__21710),
            .lcout(\pwm_generator_inst.un14_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_15_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_15_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_15_7  (
            .in0(N__21711),
            .in1(N__21663),
            .in2(N__21612),
            .in3(N__21450),
            .lcout(\pwm_generator_inst.threshold_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_4_16_0  (
            .in0(N__22751),
            .in1(N__22869),
            .in2(N__22733),
            .in3(N__22893),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_4_16_1  (
            .in0(_gnd_net_),
            .in1(N__22688),
            .in2(_gnd_net_),
            .in3(N__22709),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_4_16_2  (
            .in0(N__22854),
            .in1(N__22838),
            .in2(N__21876),
            .in3(N__22908),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_16_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_4_16_4  (
            .in0(N__22853),
            .in1(N__22839),
            .in2(N__22619),
            .in3(N__22634),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_4_16_6  (
            .in0(N__22689),
            .in1(N__22776),
            .in2(N__22713),
            .in3(N__22376),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_4_16_7  (
            .in0(N__22347),
            .in1(N__22361),
            .in2(N__21864),
            .in3(N__21846),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_17_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_4_17_2  (
            .in0(_gnd_net_),
            .in1(N__22907),
            .in2(_gnd_net_),
            .in3(N__22599),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_17_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_4_17_3  (
            .in0(N__22811),
            .in1(N__22790),
            .in2(N__21855),
            .in3(N__23072),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_4_17_4  (
            .in0(_gnd_net_),
            .in1(N__22652),
            .in2(_gnd_net_),
            .in3(N__22673),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_4_17_7  (
            .in0(N__22598),
            .in1(N__22868),
            .in2(N__22775),
            .in3(N__22892),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_18_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIVDL3_9_LC_4_18_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIVDL3_9_LC_4_18_2  (
            .in0(N__21823),
            .in1(N__21799),
            .in2(_gnd_net_),
            .in3(N__21778),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_4_18_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNISQD2_0_LC_4_18_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNISQD2_0_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__22108),
            .in2(_gnd_net_),
            .in3(N__22084),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_4_18_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_1_LC_4_18_5 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_1_LC_4_18_5  (
            .in0(N__22063),
            .in1(N__22039),
            .in2(N__22020),
            .in3(N__22012),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_4_18_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_4_18_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_5_LC_4_18_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_5_LC_4_18_6  (
            .in0(N__21993),
            .in1(N__21982),
            .in2(N__21963),
            .in3(N__21956),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_4_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_4_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36869),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50803),
            .ce(),
            .sr(N__50390));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_4_20_0  (
            .in0(_gnd_net_),
            .in1(N__23090),
            .in2(_gnd_net_),
            .in3(N__41795),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50795),
            .ce(),
            .sr(N__50394));
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_5_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_5_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_29_LC_5_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_29_LC_5_8_6  (
            .in0(N__25064),
            .in1(N__25041),
            .in2(_gnd_net_),
            .in3(N__32561),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50900),
            .ce(N__31703),
            .sr(N__50339));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_5_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_5_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_5_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23601),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50895),
            .ce(N__23281),
            .sr(N__50346));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22326),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_5_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_5_10_1 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_5_10_1  (
            .in0(N__22328),
            .in1(_gnd_net_),
            .in2(N__28629),
            .in3(N__31310),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_344_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_5_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_5_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__22327),
            .in2(_gnd_net_),
            .in3(N__28624),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_343_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_11_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_5_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37275),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50878),
            .ce(),
            .sr(N__50359));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_5_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36578),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50855),
            .ce(),
            .sr(N__50370));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_14_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_5_14_6  (
            .in0(N__22755),
            .in1(N__22620),
            .in2(N__22737),
            .in3(N__22638),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_5_14_7  (
            .in0(N__22311),
            .in1(N__22302),
            .in2(N__22296),
            .in3(N__22293),
            .lcout(\current_shift_inst.PI_CTRL.N_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_5_15_0  (
            .in0(_gnd_net_),
            .in1(N__23094),
            .in2(N__41805),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_15_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_5_15_1  (
            .in0(_gnd_net_),
            .in1(N__23352),
            .in2(N__41703),
            .in3(N__22212),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__23412),
            .in2(N__41631),
            .in3(N__22170),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(N__50940),
            .in2(N__42669),
            .in3(N__22119),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_5_15_4  (
            .in0(_gnd_net_),
            .in1(N__42568),
            .in2(N__23400),
            .in3(N__22545),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(N__23373),
            .in2(N__46899),
            .in3(N__22497),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_5_15_6  (
            .in0(_gnd_net_),
            .in1(N__46950),
            .in2(N__23481),
            .in3(N__22455),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(N__38202),
            .in2(N__42462),
            .in3(N__22425),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__50835),
            .ce(),
            .sr(N__50376));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(N__22962),
            .in2(N__42384),
            .in3(N__22380),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_16_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_5_16_1  (
            .in0(_gnd_net_),
            .in1(N__22971),
            .in2(N__42318),
            .in3(N__22365),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(N__23457),
            .in2(N__42243),
            .in3(N__22350),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(N__23421),
            .in2(N__46838),
            .in3(N__22332),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(N__23445),
            .in2(N__46248),
            .in3(N__22740),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(N__42984),
            .in2(N__23331),
            .in3(N__22716),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(N__22944),
            .in2(N__42915),
            .in3(N__22701),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_5_16_7  (
            .in0(_gnd_net_),
            .in1(N__22698),
            .in2(N__42846),
            .in3(N__22680),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__50822),
            .ce(),
            .sr(N__50380));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(N__23361),
            .in2(N__42786),
            .in3(N__22662),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__22926),
            .in2(N__42732),
            .in3(N__22641),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__22935),
            .in2(N__43527),
            .in3(N__22623),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_5_17_3  (
            .in0(_gnd_net_),
            .in1(N__23238),
            .in2(N__43473),
            .in3(N__22602),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_5_17_4  (
            .in0(_gnd_net_),
            .in1(N__43413),
            .in2(N__23385),
            .in3(N__22587),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_5_17_5  (
            .in0(_gnd_net_),
            .in1(N__22953),
            .in2(N__43362),
            .in3(N__22896),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__23112),
            .in2(N__43296),
            .in3(N__22881),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_5_17_7  (
            .in0(_gnd_net_),
            .in1(N__22878),
            .in2(N__43242),
            .in3(N__22857),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__50812),
            .ce(),
            .sr(N__50383));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_5_18_0  (
            .in0(_gnd_net_),
            .in1(N__22917),
            .in2(N__43173),
            .in3(N__22842),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_5_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(N__23433),
            .in2(N__43116),
            .in3(N__22827),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_5_18_2  (
            .in0(_gnd_net_),
            .in1(N__22824),
            .in2(N__43992),
            .in3(N__22797),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(N__23121),
            .in2(N__43932),
            .in3(N__22779),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(N__23103),
            .in2(N__43872),
            .in3(N__22758),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(N__23340),
            .in2(N__43812),
            .in3(N__23061),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_5_18_6  (
            .in0(N__46608),
            .in1(N__23466),
            .in2(_gnd_net_),
            .in3(N__23058),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50804),
            .ce(),
            .sr(N__50385));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36233),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50796),
            .ce(),
            .sr(N__50388));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_5_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_5_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36275),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50796),
            .ce(),
            .sr(N__50388));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36942),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50796),
            .ce(),
            .sr(N__50388));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_5_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_5_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36605),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50796),
            .ce(),
            .sr(N__50388));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37052),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50796),
            .ce(),
            .sr(N__50388));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_5_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36495),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50796),
            .ce(),
            .sr(N__50388));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_5_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36821),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50786),
            .ce(),
            .sr(N__50391));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_5_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_5_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37226),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50786),
            .ce(),
            .sr(N__50391));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_5_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_5_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36899),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50786),
            .ce(),
            .sr(N__50391));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_5_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_5_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37184),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50786),
            .ce(),
            .sr(N__50391));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_5_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_5_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36014),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50786),
            .ce(),
            .sr(N__50391));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_7_4_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_7_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_7_4_2  (
            .in0(N__25714),
            .in1(N__25698),
            .in2(_gnd_net_),
            .in3(N__32485),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_5_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_7_5_1  (
            .in0(N__32487),
            .in1(N__24610),
            .in2(_gnd_net_),
            .in3(N__24635),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_5_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_7_5_2  (
            .in0(N__25264),
            .in1(N__25240),
            .in2(_gnd_net_),
            .in3(N__32486),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_5_LC_7_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_5_LC_7_6_4  (
            .in0(N__32494),
            .in1(N__25906),
            .in2(_gnd_net_),
            .in3(N__25867),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50901),
            .ce(N__32169),
            .sr(N__50306));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_6_7  (
            .in0(N__28801),
            .in1(N__32493),
            .in2(_gnd_net_),
            .in3(N__28774),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_7_0  (
            .in0(N__26215),
            .in1(N__26245),
            .in2(_gnd_net_),
            .in3(N__32384),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_7_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_7_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_7_1  (
            .in0(N__32385),
            .in1(N__24932),
            .in2(_gnd_net_),
            .in3(N__24910),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_7_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_7_7_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_7_7_2  (
            .in0(N__26020),
            .in1(N__26050),
            .in2(_gnd_net_),
            .in3(N__32382),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_7_7_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_7_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_7_7_3  (
            .in0(N__32383),
            .in1(N__25316),
            .in2(_gnd_net_),
            .in3(N__25350),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_7_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_7_7_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_7_7_4  (
            .in0(N__25119),
            .in1(N__26158),
            .in2(N__25697),
            .in3(N__26095),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_7_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_7_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_7_7_5  (
            .in0(N__23607),
            .in1(N__23613),
            .in2(N__23130),
            .in3(N__23127),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_7_7_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_7_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_7_7_6  (
            .in0(N__26214),
            .in1(N__24789),
            .in2(N__32747),
            .in3(N__31801),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_7_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_7_8_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__25230),
            .in2(_gnd_net_),
            .in3(N__28764),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_8_2  (
            .in0(N__25033),
            .in1(N__25063),
            .in2(_gnd_net_),
            .in3(N__32364),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_7_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_7_8_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_7_8_3  (
            .in0(N__31401),
            .in1(N__23142),
            .in2(_gnd_net_),
            .in3(N__26367),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_7_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_7_8_4 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_7_8_4  (
            .in0(N__24600),
            .in1(N__23169),
            .in2(N__23163),
            .in3(N__23148),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_7_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_7_8_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_7_8_5  (
            .in0(N__24751),
            .in1(_gnd_net_),
            .in2(N__23160),
            .in3(N__24721),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_7_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_7_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_7_8_6  (
            .in0(N__24900),
            .in1(N__24862),
            .in2(N__25173),
            .in3(N__24963),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_7_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_7_8_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_7_8_7  (
            .in0(N__24684),
            .in1(N__25896),
            .in2(N__23157),
            .in3(N__23154),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_7_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_7_9_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_7_9_0  (
            .in0(N__24712),
            .in1(N__26011),
            .in2(N__25956),
            .in3(N__25747),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23574),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50879),
            .ce(N__23282),
            .sr(N__50332));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_7_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_7_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_7_10_0  (
            .in0(_gnd_net_),
            .in1(N__23548),
            .in2(N__23600),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_7_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_7_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__23573),
            .in2(N__23528),
            .in3(N__23136),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_7_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_7_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__23500),
            .in2(N__23553),
            .in3(N__23133),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_7_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_7_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(N__23824),
            .in2(N__23529),
            .in3(N__23199),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_7_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_7_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__23800),
            .in2(N__23505),
            .in3(N__23196),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_7_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_7_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__23776),
            .in2(N__23829),
            .in3(N__23193),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_7_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_7_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_7_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(N__23752),
            .in2(N__23805),
            .in3(N__23190),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_7_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_7_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_7_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__23728),
            .in2(N__23781),
            .in3(N__23187),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50868),
            .ce(N__23283),
            .sr(N__50340));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_7_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_7_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_7_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__23704),
            .in2(N__23757),
            .in3(N__23184),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_7_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__23680),
            .in2(N__23733),
            .in3(N__23181),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_7_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_7_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__23656),
            .in2(N__23709),
            .in3(N__23178),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_7_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_7_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__23632),
            .in2(N__23685),
            .in3(N__23175),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_7_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_7_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__24016),
            .in2(N__23661),
            .in3(N__23172),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_7_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_7_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__23992),
            .in2(N__23637),
            .in3(N__23226),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_7_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_7_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__23968),
            .in2(N__24021),
            .in3(N__23223),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_7_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_7_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__23944),
            .in2(N__23997),
            .in3(N__23220),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50856),
            .ce(N__23294),
            .sr(N__50347));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_7_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_7_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__23920),
            .in2(N__23973),
            .in3(N__23217),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_7_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_7_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__23896),
            .in2(N__23949),
            .in3(N__23214),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_7_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_7_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__23872),
            .in2(N__23925),
            .in3(N__23211),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_7_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__23848),
            .in2(N__23901),
            .in3(N__23208),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_7_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_7_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__24367),
            .in2(N__23877),
            .in3(N__23205),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_7_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__24343),
            .in2(N__23853),
            .in3(N__23202),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_7_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__24319),
            .in2(N__24372),
            .in3(N__23316),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_7_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_7_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__24298),
            .in2(N__24348),
            .in3(N__23313),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50845),
            .ce(N__23293),
            .sr(N__50353));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_7_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_7_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_7_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__24274),
            .in2(N__24324),
            .in3(N__23310),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50836),
            .ce(N__23295),
            .sr(N__50360));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_7_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_7_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__24300),
            .in2(N__24254),
            .in3(N__23307),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50836),
            .ce(N__23295),
            .sr(N__50360));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_7_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__24230),
            .in2(N__24279),
            .in3(N__23304),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50836),
            .ce(N__23295),
            .sr(N__50360));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_7_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_7_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__24074),
            .in2(N__24255),
            .in3(N__23301),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50836),
            .ce(N__23295),
            .sr(N__50360));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_7_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_7_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_7_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23298),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50836),
            .ce(N__23295),
            .sr(N__50360));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_7_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_7_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_7_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36165),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50813),
            .ce(N__36198),
            .sr(N__50371));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_7_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_7_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37023),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50805),
            .ce(),
            .sr(N__50373));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_7_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36725),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50805),
            .ce(),
            .sr(N__50373));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_7_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36443),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50805),
            .ce(),
            .sr(N__50373));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_7_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36399),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50797),
            .ce(),
            .sr(N__50377));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_7_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_7_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_7_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36983),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50797),
            .ce(),
            .sr(N__50377));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_7_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36362),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50797),
            .ce(),
            .sr(N__50377));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_7_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36524),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50797),
            .ce(),
            .sr(N__50377));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_7_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35966),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50787),
            .ce(),
            .sr(N__50381));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37149),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50787),
            .ce(),
            .sr(N__50381));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_7_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36648),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50787),
            .ce(),
            .sr(N__50381));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_7_18_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__36320),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50787),
            .ce(),
            .sr(N__50381));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_7_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_7_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_7_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37101),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50787),
            .ce(),
            .sr(N__50381));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_19_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_7_19_3  (
            .in0(N__33952),
            .in1(N__34339),
            .in2(N__35802),
            .in3(N__30329),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_19_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_7_19_6  (
            .in0(N__34338),
            .in1(N__33953),
            .in2(N__35886),
            .in3(N__33284),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36761),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50774),
            .ce(),
            .sr(N__50386));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_7_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_7_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_7_20_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_7_20_4  (
            .in0(N__41568),
            .in1(N__46329),
            .in2(_gnd_net_),
            .in3(N__46770),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50774),
            .ce(),
            .sr(N__50386));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_7_20_5 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_7_20_5  (
            .in0(N__46769),
            .in1(N__46607),
            .in2(N__46386),
            .in3(N__42519),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50774),
            .ce(),
            .sr(N__50386));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36684),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50774),
            .ce(),
            .sr(N__50386));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37316),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50774),
            .ce(),
            .sr(N__50386));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_5_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_8_5_5  (
            .in0(N__25786),
            .in1(N__25763),
            .in2(_gnd_net_),
            .in3(N__32492),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_6_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_6_2  (
            .in0(N__25199),
            .in1(N__25174),
            .in2(_gnd_net_),
            .in3(N__32489),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_8_6_4  (
            .in0(N__24824),
            .in1(N__24799),
            .in2(_gnd_net_),
            .in3(N__32491),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_8_6_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_8_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_8_6_6  (
            .in0(N__25871),
            .in1(N__25907),
            .in2(_gnd_net_),
            .in3(N__32490),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_6_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_6_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_6_7  (
            .in0(N__32488),
            .in1(N__28873),
            .in2(_gnd_net_),
            .in3(N__28847),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_8_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_8_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_31_LC_8_7_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_31_LC_8_7_1  (
            .in0(N__24612),
            .in1(N__24636),
            .in2(_gnd_net_),
            .in3(N__32433),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50887),
            .ce(N__32074),
            .sr(N__50307));
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_8_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_8_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_11_LC_8_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_11_LC_8_7_5  (
            .in0(N__24928),
            .in1(N__24911),
            .in2(_gnd_net_),
            .in3(N__32432),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50887),
            .ce(N__32074),
            .sr(N__50307));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_8_8_0  (
            .in0(N__24654),
            .in1(N__24685),
            .in2(_gnd_net_),
            .in3(N__32390),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_8_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_8_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_8_8_2  (
            .in0(N__27341),
            .in1(N__27312),
            .in2(_gnd_net_),
            .in3(N__32388),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_8_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_8_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_8_8_3  (
            .in0(N__32389),
            .in1(N__24882),
            .in2(_gnd_net_),
            .in3(N__24858),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_8_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_8_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_8_8_4  (
            .in0(N__32812),
            .in1(N__32223),
            .in2(N__31745),
            .in3(N__25357),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_8_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_8_5  (
            .in0(N__32387),
            .in1(_gnd_net_),
            .in2(N__24995),
            .in3(N__24964),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_8_6  (
            .in0(N__25087),
            .in1(N__25129),
            .in2(_gnd_net_),
            .in3(N__32386),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_7  (
            .in0(N__25032),
            .in1(N__26609),
            .in2(N__27317),
            .in3(N__28839),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_8_9_0  (
            .in0(N__24213),
            .in1(N__23593),
            .in2(_gnd_net_),
            .in3(N__23577),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_8_9_1  (
            .in0(N__24209),
            .in1(N__23572),
            .in2(_gnd_net_),
            .in3(N__23556),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_8_9_2  (
            .in0(N__24214),
            .in1(N__23549),
            .in2(_gnd_net_),
            .in3(N__23532),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_8_9_3  (
            .in0(N__24210),
            .in1(N__23527),
            .in2(_gnd_net_),
            .in3(N__23508),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_8_9_4  (
            .in0(N__24215),
            .in1(N__23501),
            .in2(_gnd_net_),
            .in3(N__23484),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_8_9_5  (
            .in0(N__24211),
            .in1(N__23825),
            .in2(_gnd_net_),
            .in3(N__23808),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_8_9_6  (
            .in0(N__24216),
            .in1(N__23801),
            .in2(_gnd_net_),
            .in3(N__23784),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_8_9_7  (
            .in0(N__24212),
            .in1(N__23777),
            .in2(_gnd_net_),
            .in3(N__23760),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__50869),
            .ce(N__24062),
            .sr(N__50323));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_8_10_0  (
            .in0(N__24167),
            .in1(N__23753),
            .in2(_gnd_net_),
            .in3(N__23736),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_8_10_1  (
            .in0(N__24171),
            .in1(N__23729),
            .in2(_gnd_net_),
            .in3(N__23712),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_8_10_2  (
            .in0(N__24164),
            .in1(N__23705),
            .in2(_gnd_net_),
            .in3(N__23688),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_8_10_3  (
            .in0(N__24168),
            .in1(N__23681),
            .in2(_gnd_net_),
            .in3(N__23664),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_8_10_4  (
            .in0(N__24165),
            .in1(N__23657),
            .in2(_gnd_net_),
            .in3(N__23640),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_8_10_5  (
            .in0(N__24169),
            .in1(N__23633),
            .in2(_gnd_net_),
            .in3(N__23616),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_8_10_6  (
            .in0(N__24166),
            .in1(N__24017),
            .in2(_gnd_net_),
            .in3(N__24000),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_8_10_7  (
            .in0(N__24170),
            .in1(N__23993),
            .in2(_gnd_net_),
            .in3(N__23976),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__50857),
            .ce(N__24060),
            .sr(N__50333));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_8_11_0  (
            .in0(N__24172),
            .in1(N__23969),
            .in2(_gnd_net_),
            .in3(N__23952),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_8_11_1  (
            .in0(N__24176),
            .in1(N__23945),
            .in2(_gnd_net_),
            .in3(N__23928),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_8_11_2  (
            .in0(N__24173),
            .in1(N__23921),
            .in2(_gnd_net_),
            .in3(N__23904),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_8_11_3  (
            .in0(N__24177),
            .in1(N__23897),
            .in2(_gnd_net_),
            .in3(N__23880),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_8_11_4  (
            .in0(N__24174),
            .in1(N__23873),
            .in2(_gnd_net_),
            .in3(N__23856),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_8_11_5  (
            .in0(N__24178),
            .in1(N__23849),
            .in2(_gnd_net_),
            .in3(N__23832),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_8_11_6  (
            .in0(N__24175),
            .in1(N__24368),
            .in2(_gnd_net_),
            .in3(N__24351),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_8_11_7  (
            .in0(N__24179),
            .in1(N__24344),
            .in2(_gnd_net_),
            .in3(N__24327),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__50846),
            .ce(N__24061),
            .sr(N__50341));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_8_12_0  (
            .in0(N__24203),
            .in1(N__24320),
            .in2(_gnd_net_),
            .in3(N__24303),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__50837),
            .ce(N__24063),
            .sr(N__50348));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_8_12_1  (
            .in0(N__24207),
            .in1(N__24299),
            .in2(_gnd_net_),
            .in3(N__24282),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__50837),
            .ce(N__24063),
            .sr(N__50348));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_8_12_2  (
            .in0(N__24204),
            .in1(N__24275),
            .in2(_gnd_net_),
            .in3(N__24258),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__50837),
            .ce(N__24063),
            .sr(N__50348));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_8_12_3  (
            .in0(N__24208),
            .in1(N__24253),
            .in2(_gnd_net_),
            .in3(N__24234),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__50837),
            .ce(N__24063),
            .sr(N__50348));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_8_12_4  (
            .in0(N__24205),
            .in1(N__24231),
            .in2(_gnd_net_),
            .in3(N__24219),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__50837),
            .ce(N__24063),
            .sr(N__50348));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_12_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_8_12_5  (
            .in0(N__24075),
            .in1(N__24206),
            .in2(_gnd_net_),
            .in3(N__24078),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50837),
            .ce(N__24063),
            .sr(N__50348));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31482),
            .lcout(\phase_controller_inst2.start_latched ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50823),
            .ce(),
            .sr(N__50354));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_8_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_8_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_8_14_4  (
            .in0(N__34315),
            .in1(N__35534),
            .in2(N__33963),
            .in3(N__30407),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_8_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_8_14_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_8_14_5  (
            .in0(N__38347),
            .in1(N__33859),
            .in2(N__38394),
            .in3(N__34316),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_8_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_8_15_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_8_15_5  (
            .in0(N__34198),
            .in1(N__33784),
            .in2(N__35937),
            .in3(N__33138),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_8_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_8_15_6 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_8_15_6  (
            .in0(N__33783),
            .in1(N__34197),
            .in2(N__35142),
            .in3(N__30065),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_8_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_8_16_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_8_16_0  (
            .in0(N__33781),
            .in1(N__34132),
            .in2(N__35196),
            .in3(N__30102),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_8_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_8_16_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_8_16_1  (
            .in0(N__34131),
            .in1(N__33018),
            .in2(_gnd_net_),
            .in3(N__24378),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_8_16_2  (
            .in0(N__49784),
            .in1(N__24384),
            .in2(_gnd_net_),
            .in3(N__31839),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_8_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_8_16_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_8_16_3  (
            .in0(N__34133),
            .in1(N__33782),
            .in2(N__38616),
            .in3(N__38571),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31869),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_16_6 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(N__34130),
            .in2(N__24426),
            .in3(N__33017),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__24423),
            .in2(N__25569),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_8_17_1  (
            .in0(_gnd_net_),
            .in1(N__29808),
            .in2(N__25398),
            .in3(N__28673),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_8_17_2  (
            .in0(N__28674),
            .in1(N__33484),
            .in2(N__25488),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_8_17_3  (
            .in0(_gnd_net_),
            .in1(N__25386),
            .in2(N__33670),
            .in3(N__24417),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_8_17_4  (
            .in0(_gnd_net_),
            .in1(N__33488),
            .in2(N__26514),
            .in3(N__24414),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_8_17_5  (
            .in0(_gnd_net_),
            .in1(N__33502),
            .in2(N__25410),
            .in3(N__24411),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(N__33489),
            .in2(N__24408),
            .in3(N__24399),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_8_17_7  (
            .in0(_gnd_net_),
            .in1(N__33503),
            .in2(N__24396),
            .in3(N__24387),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__24483),
            .in2(N__33762),
            .in3(N__24474),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__33581),
            .in2(N__25440),
            .in3(N__24471),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__25446),
            .in2(N__33763),
            .in3(N__24468),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_8_18_3  (
            .in0(_gnd_net_),
            .in1(N__33585),
            .in2(N__25479),
            .in3(N__24465),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_8_18_4  (
            .in0(_gnd_net_),
            .in1(N__24462),
            .in2(N__33764),
            .in3(N__24453),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_8_18_5  (
            .in0(_gnd_net_),
            .in1(N__33589),
            .in2(N__26481),
            .in3(N__24450),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_8_18_6  (
            .in0(_gnd_net_),
            .in1(N__25461),
            .in2(N__33765),
            .in3(N__24447),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_8_18_7  (
            .in0(_gnd_net_),
            .in1(N__33593),
            .in2(N__24444),
            .in3(N__24432),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__33690),
            .in2(N__25425),
            .in3(N__24429),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_8_19_1  (
            .in0(_gnd_net_),
            .in1(N__25455),
            .in2(N__33867),
            .in3(N__24540),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_8_19_2  (
            .in0(_gnd_net_),
            .in1(N__33694),
            .in2(N__26451),
            .in3(N__24537),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_8_19_3  (
            .in0(_gnd_net_),
            .in1(N__24534),
            .in2(N__33868),
            .in3(N__24522),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_8_19_4  (
            .in0(_gnd_net_),
            .in1(N__33698),
            .in2(N__24519),
            .in3(N__24510),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_8_19_5  (
            .in0(_gnd_net_),
            .in1(N__26697),
            .in2(N__33869),
            .in3(N__24507),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_8_19_6  (
            .in0(_gnd_net_),
            .in1(N__33702),
            .in2(N__24504),
            .in3(N__24495),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_8_19_7  (
            .in0(_gnd_net_),
            .in1(N__25470),
            .in2(N__33870),
            .in3(N__24492),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_8_20_0  (
            .in0(_gnd_net_),
            .in1(N__33746),
            .in2(N__33321),
            .in3(N__24489),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_8_20_1  (
            .in0(_gnd_net_),
            .in1(N__26727),
            .in2(N__33896),
            .in3(N__24486),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_8_20_2  (
            .in0(_gnd_net_),
            .in1(N__33750),
            .in2(N__26886),
            .in3(N__24573),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__26622),
            .in2(N__33897),
            .in3(N__24570),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__33754),
            .in2(N__26652),
            .in3(N__24567),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_8_20_5  (
            .in0(_gnd_net_),
            .in1(N__24555),
            .in2(N__33898),
            .in3(N__24564),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_8_20_6  (
            .in0(_gnd_net_),
            .in1(N__33758),
            .in2(N__24549),
            .in3(N__24561),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_20_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_8_20_7  (
            .in0(N__31935),
            .in1(N__25815),
            .in2(N__34750),
            .in3(N__24558),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_8_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_8_21_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_8_21_0  (
            .in0(N__34334),
            .in1(N__36078),
            .in2(N__33971),
            .in3(N__30788),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_8_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_8_21_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_8_21_4  (
            .in0(N__34333),
            .in1(N__30330),
            .in2(N__33970),
            .in3(N__35801),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_8_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_8_21_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_8_21_5  (
            .in0(N__30612),
            .in1(N__33895),
            .in2(N__28694),
            .in3(N__34335),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_9_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_3_LC_9_5_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_3_LC_9_5_2  (
            .in0(N__24759),
            .in1(N__24732),
            .in2(_gnd_net_),
            .in3(N__32666),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50896),
            .ce(N__31696),
            .sr(N__50283));
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_9_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_8_LC_9_5_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_8_LC_9_5_3  (
            .in0(N__32664),
            .in1(N__25265),
            .in2(_gnd_net_),
            .in3(N__25245),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50896),
            .ce(N__31696),
            .sr(N__50283));
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_31_LC_9_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_31_LC_9_5_6  (
            .in0(N__24634),
            .in1(N__24611),
            .in2(_gnd_net_),
            .in3(N__32665),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50896),
            .ce(N__31696),
            .sr(N__50283));
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_22_LC_9_6_1  (
            .in0(N__32660),
            .in1(N__26109),
            .in2(_gnd_net_),
            .in3(N__26124),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50888),
            .ce(N__31700),
            .sr(N__50293));
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_9_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_9_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_13_LC_9_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_13_LC_9_6_2  (
            .in0(N__24820),
            .in1(N__24804),
            .in2(_gnd_net_),
            .in3(N__32662),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50888),
            .ce(N__31700),
            .sr(N__50293));
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_9_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_9_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_21_LC_9_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_21_LC_9_6_4  (
            .in0(N__25092),
            .in1(N__25134),
            .in2(_gnd_net_),
            .in3(N__32663),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50888),
            .ce(N__31700),
            .sr(N__50293));
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_12_LC_9_6_6  (
            .in0(N__25195),
            .in1(N__25179),
            .in2(_gnd_net_),
            .in3(N__32661),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50888),
            .ce(N__31700),
            .sr(N__50293));
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_9_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_20_LC_9_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_20_LC_9_7_1  (
            .in0(N__25312),
            .in1(N__25362),
            .in2(_gnd_net_),
            .in3(N__32606),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50880),
            .ce(N__31702),
            .sr(N__50300));
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_27_LC_9_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_27_LC_9_7_3  (
            .in0(N__26394),
            .in1(N__26373),
            .in2(_gnd_net_),
            .in3(N__32607),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50880),
            .ce(N__31702),
            .sr(N__50300));
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_6_LC_9_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_6_LC_9_7_4  (
            .in0(N__32604),
            .in1(N__24692),
            .in2(_gnd_net_),
            .in3(N__24653),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50880),
            .ce(N__31702),
            .sr(N__50300));
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_9_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_10_LC_9_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_10_LC_9_7_5  (
            .in0(N__24881),
            .in1(N__24864),
            .in2(_gnd_net_),
            .in3(N__32605),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50880),
            .ce(N__31702),
            .sr(N__50300));
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_11_LC_9_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_11_LC_9_7_6  (
            .in0(N__32603),
            .in1(N__24933),
            .in2(_gnd_net_),
            .in3(N__24912),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50880),
            .ce(N__31702),
            .sr(N__50300));
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_9_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_9_LC_9_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_9_LC_9_7_7  (
            .in0(N__24996),
            .in1(N__24969),
            .in2(_gnd_net_),
            .in3(N__32608),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50880),
            .ce(N__31702),
            .sr(N__50300));
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_10_LC_9_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_10_LC_9_8_1  (
            .in0(N__24880),
            .in1(N__24863),
            .in2(_gnd_net_),
            .in3(N__32564),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50870),
            .ce(N__32176),
            .sr(N__50308));
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_13_LC_9_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_13_LC_9_8_6  (
            .in0(N__32639),
            .in1(N__24825),
            .in2(_gnd_net_),
            .in3(N__24800),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50870),
            .ce(N__32176),
            .sr(N__50308));
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_9_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_9_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_17_LC_9_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_17_LC_9_8_7  (
            .in0(N__31762),
            .in1(N__31740),
            .in2(_gnd_net_),
            .in3(N__32565),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50870),
            .ce(N__32176),
            .sr(N__50308));
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_9_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_3_LC_9_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_3_LC_9_9_0  (
            .in0(N__32667),
            .in1(N__24758),
            .in2(_gnd_net_),
            .in3(N__24731),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50858),
            .ce(N__32134),
            .sr(N__50316));
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_9_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_9_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_30_LC_9_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_30_LC_9_9_2  (
            .in0(N__27340),
            .in1(N__27316),
            .in2(_gnd_net_),
            .in3(N__32650),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50858),
            .ce(N__32134),
            .sr(N__50316));
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_6_LC_9_9_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_6_LC_9_9_3  (
            .in0(N__32644),
            .in1(_gnd_net_),
            .in2(N__24696),
            .in3(N__24652),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50858),
            .ce(N__32134),
            .sr(N__50316));
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_9_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_9_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_7_LC_9_9_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_7_LC_9_9_4  (
            .in0(N__28806),
            .in1(N__32648),
            .in2(_gnd_net_),
            .in3(N__28778),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50858),
            .ce(N__32134),
            .sr(N__50316));
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_9_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_9_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_8_LC_9_9_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_8_LC_9_9_5  (
            .in0(N__25269),
            .in1(_gnd_net_),
            .in2(N__32694),
            .in3(N__25244),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50858),
            .ce(N__32134),
            .sr(N__50316));
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_1_LC_9_9_6  (
            .in0(N__25791),
            .in1(N__25762),
            .in2(_gnd_net_),
            .in3(N__32649),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50858),
            .ce(N__32134),
            .sr(N__50316));
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_12_LC_9_10_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_12_LC_9_10_0  (
            .in0(N__25203),
            .in1(N__25178),
            .in2(_gnd_net_),
            .in3(N__32654),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_9_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_9_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_21_LC_9_10_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_21_LC_9_10_2  (
            .in0(N__32659),
            .in1(N__25130),
            .in2(_gnd_net_),
            .in3(N__25091),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_29_LC_9_10_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_29_LC_9_10_3  (
            .in0(N__32653),
            .in1(N__25068),
            .in2(_gnd_net_),
            .in3(N__25040),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_9_LC_9_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_9_LC_9_10_4  (
            .in0(N__24991),
            .in1(N__24965),
            .in2(_gnd_net_),
            .in3(N__32656),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_15_LC_9_10_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_15_LC_9_10_5  (
            .in0(N__32651),
            .in1(N__26250),
            .in2(_gnd_net_),
            .in3(N__26222),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_9_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_9_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_25_LC_9_10_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_25_LC_9_10_6  (
            .in0(N__28878),
            .in1(N__28846),
            .in2(_gnd_net_),
            .in3(N__32655),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_9_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_9_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_24_LC_9_10_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_24_LC_9_10_7  (
            .in0(N__32652),
            .in1(_gnd_net_),
            .in2(N__25728),
            .in3(N__25696),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50847),
            .ce(N__32177),
            .sr(N__50324));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_11_0  (
            .in0(N__25380),
            .in1(N__28218),
            .in2(N__28247),
            .in3(N__25371),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_9_11_2  (
            .in0(N__32611),
            .in1(N__25991),
            .in2(_gnd_net_),
            .in3(N__25966),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_4 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_9_11_4  (
            .in0(N__25379),
            .in1(N__28217),
            .in2(N__28248),
            .in3(N__25370),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_9_11_5  (
            .in0(N__26393),
            .in1(N__26368),
            .in2(_gnd_net_),
            .in3(N__32612),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_12_0  (
            .in0(N__28322),
            .in1(N__25283),
            .in2(N__28350),
            .in3(N__25293),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_9_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_20_LC_9_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_20_LC_9_12_2  (
            .in0(N__25361),
            .in1(N__25320),
            .in2(_gnd_net_),
            .in3(N__32658),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50824),
            .ce(N__32178),
            .sr(N__50342));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_12_5 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_9_12_5  (
            .in0(N__25292),
            .in1(N__28349),
            .in2(N__25284),
            .in3(N__28323),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_9_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_2_LC_9_12_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_2_LC_9_12_7  (
            .in0(N__32657),
            .in1(N__25987),
            .in2(_gnd_net_),
            .in3(N__25970),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50824),
            .ce(N__32178),
            .sr(N__50342));
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_9_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_9_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_26_LC_9_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_26_LC_9_13_2  (
            .in0(N__26610),
            .in1(N__26319),
            .in2(_gnd_net_),
            .in3(N__32693),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50814),
            .ce(N__31704),
            .sr(N__50349));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_14_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_9_14_0  (
            .in0(N__34288),
            .in1(N__35094),
            .in2(N__33976),
            .in3(N__31910),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_9_14_2  (
            .in0(N__34289),
            .in1(N__35438),
            .in2(N__33977),
            .in3(N__30182),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_15_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_9_15_1  (
            .in0(N__33787),
            .in1(N__34247),
            .in2(N__35195),
            .in3(N__30101),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_9_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_9_15_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_9_15_2  (
            .in0(N__49726),
            .in1(N__28672),
            .in2(_gnd_net_),
            .in3(N__25544),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_15_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_9_15_3  (
            .in0(N__33785),
            .in1(N__34248),
            .in2(N__31917),
            .in3(N__35093),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_15_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_9_15_6  (
            .in0(N__34246),
            .in1(N__33786),
            .in2(N__35237),
            .in3(N__30134),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_15_7 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_9_15_7  (
            .in0(N__29816),
            .in1(N__29772),
            .in2(N__29712),
            .in3(N__34245),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_16_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_9_16_4  (
            .in0(N__34177),
            .in1(N__35315),
            .in2(N__33855),
            .in3(N__32981),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36164),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50788),
            .ce(N__36196),
            .sr(N__50364));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_9_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_9_16_7 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_9_16_7  (
            .in0(N__35351),
            .in1(N__34176),
            .in2(N__29688),
            .in3(N__33661),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_9_17_0  (
            .in0(N__34183),
            .in1(N__38064),
            .in2(N__33789),
            .in3(N__38031),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_1 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_9_17_1  (
            .in0(N__30372),
            .in1(N__33628),
            .in2(N__35748),
            .in3(N__34191),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_9_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_9_17_2 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_9_17_2  (
            .in0(N__33627),
            .in1(N__38112),
            .in2(N__34287),
            .in3(N__30218),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_17_3 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_9_17_3  (
            .in0(N__37940),
            .in1(N__33629),
            .in2(N__37983),
            .in3(N__34190),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_9_17_4  (
            .in0(N__34180),
            .in1(N__35316),
            .in2(N__33788),
            .in3(N__32988),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_17_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_9_17_5  (
            .in0(N__30027),
            .in1(N__33621),
            .in2(N__35058),
            .in3(N__34182),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_9_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_9_17_6 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_9_17_6  (
            .in0(N__33626),
            .in1(N__30249),
            .in2(N__34286),
            .in3(N__35487),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_17_7 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_9_17_7  (
            .in0(N__35238),
            .in1(N__33622),
            .in2(N__30138),
            .in3(N__34181),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__25565),
            .in2(N__25548),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(N__29809),
            .in2(N__29790),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(N__33490),
            .in2(N__26736),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_9_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__25530),
            .in2(N__33671),
            .in3(N__25524),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_9_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__33494),
            .in2(N__26706),
            .in3(N__25521),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_9_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__25518),
            .in2(N__33672),
            .in3(N__25512),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__33498),
            .in2(N__25509),
            .in3(N__25497),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__26673),
            .in2(N__33673),
            .in3(N__25494),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__33674),
            .in2(N__26634),
            .in3(N__25491),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25614),
            .in2(N__33863),
            .in3(N__25605),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__33678),
            .in2(N__26466),
            .in3(N__25602),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__26745),
            .in2(N__33864),
            .in3(N__25599),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__33682),
            .in2(N__26811),
            .in3(N__25596),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__25593),
            .in2(N__33865),
            .in3(N__25584),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__33686),
            .in2(N__26895),
            .in3(N__25581),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__26436),
            .in2(N__33866),
            .in3(N__25578),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__33706),
            .in2(N__26496),
            .in3(N__25575),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__26790),
            .in2(N__33871),
            .in3(N__25572),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__33710),
            .in2(N__26904),
            .in3(N__25650),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__26685),
            .in2(N__33872),
            .in3(N__25647),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__33714),
            .in2(N__26802),
            .in3(N__25644),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__26769),
            .in2(N__33873),
            .in3(N__25641),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__33718),
            .in2(N__25638),
            .in3(N__25629),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__26715),
            .in2(N__33874),
            .in3(N__25626),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__33875),
            .in2(N__26919),
            .in3(N__25623),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__26817),
            .in2(N__33967),
            .in3(N__25620),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__33879),
            .in2(N__27006),
            .in3(N__25617),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__26664),
            .in2(N__33968),
            .in3(N__25830),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__33883),
            .in2(N__26874),
            .in3(N__25827),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__27012),
            .in2(N__33969),
            .in3(N__25824),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_9_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_9_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__33887),
            .in2(N__28644),
            .in3(N__25821),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_9_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_9_21_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_9_21_7  (
            .in0(N__33888),
            .in1(N__34336),
            .in2(_gnd_net_),
            .in3(N__25818),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_4.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_9_30_4 (
            .in0(N__25809),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_er_LC_10_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_er_LC_10_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_er_LC_10_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_er_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29084),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50889),
            .ce(N__26277),
            .sr(N__50262));
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_1_LC_10_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_1_LC_10_5_4  (
            .in0(N__25787),
            .in1(N__25764),
            .in2(_gnd_net_),
            .in3(N__32682),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50881),
            .ce(N__31694),
            .sr(N__50269));
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_10_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_10_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_24_LC_10_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_24_LC_10_5_5  (
            .in0(N__32681),
            .in1(N__25724),
            .in2(_gnd_net_),
            .in3(N__25695),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50881),
            .ce(N__31694),
            .sr(N__50269));
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_2_LC_10_5_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_2_LC_10_5_6  (
            .in0(N__25995),
            .in1(N__25971),
            .in2(_gnd_net_),
            .in3(N__32683),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50881),
            .ce(N__31694),
            .sr(N__50269));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_6_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_6_0  (
            .in0(N__29300),
            .in1(N__25929),
            .in2(N__25920),
            .in3(N__29642),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_10_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_10_6_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_10_6_1  (
            .in0(N__25928),
            .in1(N__29301),
            .in2(N__29643),
            .in3(N__25916),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_23_LC_10_6_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_23_LC_10_6_3  (
            .in0(N__26172),
            .in1(N__32679),
            .in2(_gnd_net_),
            .in3(N__26187),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50872),
            .ce(N__31695),
            .sr(N__50275));
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_4_LC_10_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_4_LC_10_6_6  (
            .in0(N__32678),
            .in1(N__26057),
            .in2(_gnd_net_),
            .in3(N__26031),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50872),
            .ce(N__31695),
            .sr(N__50275));
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_5_LC_10_6_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_5_LC_10_6_7  (
            .in0(N__25908),
            .in1(N__25872),
            .in2(_gnd_net_),
            .in3(N__32680),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50872),
            .ce(N__31695),
            .sr(N__50275));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_7_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_10_7_0  (
            .in0(N__29351),
            .in1(N__25851),
            .in2(N__25842),
            .in3(N__29327),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_7_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_10_7_1  (
            .in0(N__25850),
            .in1(N__29352),
            .in2(N__29328),
            .in3(N__25838),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_10_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_10_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_14_LC_10_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_14_LC_10_7_5  (
            .in0(N__32745),
            .in1(N__32768),
            .in2(_gnd_net_),
            .in3(N__32610),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50860),
            .ce(N__31697),
            .sr(N__50284));
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_10_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_10_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_15_LC_10_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_15_LC_10_7_6  (
            .in0(N__32609),
            .in1(N__26246),
            .in2(_gnd_net_),
            .in3(N__26223),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50860),
            .ce(N__31697),
            .sr(N__50284));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_10_8_0  (
            .in0(N__28272),
            .in1(N__28295),
            .in2(N__26136),
            .in3(N__26070),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_10_8_1  (
            .in0(N__26069),
            .in1(N__28271),
            .in2(N__28299),
            .in3(N__26132),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_10_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_10_8_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_10_8_2  (
            .in0(N__32674),
            .in1(N__26167),
            .in2(_gnd_net_),
            .in3(N__26183),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(elapsed_time_ns_1_RNI1CPBB_0_23_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_23_LC_10_8_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_23_LC_10_8_3  (
            .in0(N__26168),
            .in1(_gnd_net_),
            .in2(N__26139),
            .in3(N__32676),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50849),
            .ce(N__32171),
            .sr(N__50294));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_8_4  (
            .in0(N__32673),
            .in1(N__26107),
            .in2(_gnd_net_),
            .in3(N__26120),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(elapsed_time_ns_1_RNI0BPBB_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_22_LC_10_8_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_22_LC_10_8_5  (
            .in0(N__26108),
            .in1(_gnd_net_),
            .in2(N__26073),
            .in3(N__32675),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50849),
            .ce(N__32171),
            .sr(N__50294));
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_4_LC_10_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_4_LC_10_8_7  (
            .in0(N__26061),
            .in1(N__26027),
            .in2(_gnd_net_),
            .in3(N__32677),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50849),
            .ce(N__32171),
            .sr(N__50294));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_9_0 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_9_0  (
            .in0(N__28035),
            .in1(N__26304),
            .in2(N__28065),
            .in3(N__26295),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_9_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_10_9_1  (
            .in0(N__31810),
            .in1(N__31778),
            .in2(_gnd_net_),
            .in3(N__32670),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_10_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_10_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_16_LC_10_9_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_16_LC_10_9_2  (
            .in0(N__32672),
            .in1(_gnd_net_),
            .in2(N__26307),
            .in3(N__31811),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50838),
            .ce(N__32133),
            .sr(N__50301));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_9_4 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_9_4  (
            .in0(N__28034),
            .in1(N__26303),
            .in2(N__28064),
            .in3(N__26294),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_5  (
            .in0(N__31741),
            .in1(N__31766),
            .in2(_gnd_net_),
            .in3(N__32671),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_10_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_10_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_10_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_10_10_0  (
            .in0(N__31224),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.start_latched ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50826),
            .ce(),
            .sr(N__50309));
    defparam \phase_controller_inst1.stoper_tr.running_LC_10_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_10_10_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_10_10_1  (
            .in0(N__29074),
            .in1(N__26266),
            .in2(_gnd_net_),
            .in3(N__26286),
            .lcout(\phase_controller_inst1.running ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50826),
            .ce(),
            .sr(N__50309));
    defparam \phase_controller_inst1.stoper_hc.m42_LC_10_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m42_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m42_LC_10_10_2 .LUT_INIT=16'b1101110101011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.m42_LC_10_10_2  (
            .in0(N__31223),
            .in1(N__29073),
            .in2(N__26268),
            .in3(N__27726),
            .lcout(\phase_controller_inst1.N_43 ),
            .ltout(\phase_controller_inst1.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_sbtinv_LC_10_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_sbtinv_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_sbtinv_LC_10_10_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_sbtinv_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26280),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.N_43_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.m41_LC_10_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m41_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m41_LC_10_10_4 .LUT_INIT=16'b0101110111011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.m41_LC_10_10_4  (
            .in0(N__31222),
            .in1(N__29072),
            .in2(N__26267),
            .in3(N__27725),
            .lcout(\phase_controller_inst1.N_42 ),
            .ltout(\phase_controller_inst1.N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_10_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_10_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_10_10_5 .LUT_INIT=16'b0011000000000011;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_10_10_5  (
            .in0(_gnd_net_),
            .in1(N__32172),
            .in2(N__26424),
            .in3(N__27707),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50826),
            .ce(),
            .sr(N__50309));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_11_0 .LUT_INIT=16'b0010001010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_10_11_0  (
            .in0(N__26418),
            .in1(N__28446),
            .in2(N__26409),
            .in3(N__28470),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_11_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_10_11_1  (
            .in0(N__31402),
            .in1(N__32622),
            .in2(_gnd_net_),
            .in3(N__31358),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(elapsed_time_ns_1_RNI6HPBB_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_28_LC_10_11_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_28_LC_10_11_2  (
            .in0(N__32623),
            .in1(_gnd_net_),
            .in2(N__26421),
            .in3(N__31403),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50816),
            .ce(N__32135),
            .sr(N__50317));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_11_4 .LUT_INIT=16'b1011001010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_10_11_4  (
            .in0(N__26417),
            .in1(N__28445),
            .in2(N__26408),
            .in3(N__28469),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_7 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_7  (
            .in0(N__26562),
            .in1(N__28391),
            .in2(N__26546),
            .in3(N__28422),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_12_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_12_0  (
            .in0(N__26571),
            .in1(N__28493),
            .in2(N__26331),
            .in3(N__28194),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_12_1 .LUT_INIT=16'b1101111100001101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_10_12_1  (
            .in0(N__28193),
            .in1(N__26570),
            .in2(N__28497),
            .in3(N__26327),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_10_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_10_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_27_LC_10_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_27_LC_10_12_3  (
            .in0(N__26389),
            .in1(N__26369),
            .in2(_gnd_net_),
            .in3(N__32626),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50807),
            .ce(N__32170),
            .sr(N__50325));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_12_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_10_12_4  (
            .in0(N__32624),
            .in1(N__26604),
            .in2(_gnd_net_),
            .in3(N__26318),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_10_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_10_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_26_LC_10_12_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_26_LC_10_12_5  (
            .in0(N__26605),
            .in1(_gnd_net_),
            .in2(N__26574),
            .in3(N__32625),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50807),
            .ce(N__32170),
            .sr(N__50325));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_12_7 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_10_12_7  (
            .in0(N__26561),
            .in1(N__28392),
            .in2(N__26547),
            .in3(N__28418),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_13_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_10_13_3  (
            .in0(N__34282),
            .in1(N__35273),
            .in2(N__33989),
            .in3(N__32924),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_14_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_10_14_2  (
            .in0(N__38517),
            .in1(N__35050),
            .in2(_gnd_net_),
            .in3(N__30016),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_10_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_10_14_3 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_10_14_3  (
            .in0(N__30183),
            .in1(N__33915),
            .in2(N__35439),
            .in3(N__34285),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_10_14_4  (
            .in0(N__34284),
            .in1(N__35483),
            .in2(N__33978),
            .in3(N__30247),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_14_5 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_10_14_5  (
            .in0(N__35051),
            .in1(N__34283),
            .in2(N__30023),
            .in3(N__33911),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_15_1 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_10_15_1  (
            .in0(N__33959),
            .in1(N__34213),
            .in2(N__30536),
            .in3(N__35393),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_15_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_10_15_2  (
            .in0(N__34212),
            .in1(N__33962),
            .in2(N__38355),
            .in3(N__38387),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_10_15_4  (
            .in0(N__38499),
            .in1(N__35344),
            .in2(_gnd_net_),
            .in3(N__29680),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_15_5 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_10_15_5  (
            .in0(N__33960),
            .in1(N__33083),
            .in2(N__35844),
            .in3(N__34215),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_10_15_6  (
            .in0(N__38500),
            .in1(N__35224),
            .in2(_gnd_net_),
            .in3(N__30133),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_15_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_10_15_7  (
            .in0(N__33961),
            .in1(N__34214),
            .in2(N__35936),
            .in3(N__33137),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_10_16_0  (
            .in0(N__34192),
            .in1(N__38612),
            .in2(N__33981),
            .in3(N__38570),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_16_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_10_16_1  (
            .in0(N__35574),
            .in1(N__34195),
            .in2(N__30288),
            .in3(N__33920),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_10_16_2  (
            .in0(N__34196),
            .in1(N__36125),
            .in2(N__33980),
            .in3(N__31109),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_10_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_10_16_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_10_16_5  (
            .in0(N__30064),
            .in1(N__33927),
            .in2(N__35138),
            .in3(N__34193),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_10_16_6  (
            .in0(N__34194),
            .in1(N__35573),
            .in2(N__33979),
            .in3(N__30283),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_17_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_10_17_0  (
            .in0(N__34179),
            .in1(N__38060),
            .in2(N__33916),
            .in3(N__38030),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_17_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_10_17_1  (
            .in0(N__33793),
            .in1(N__34178),
            .in2(N__35355),
            .in3(N__29684),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_10_17_2  (
            .in0(N__38101),
            .in1(N__38528),
            .in2(_gnd_net_),
            .in3(N__30217),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_10_17_3  (
            .in0(N__38529),
            .in1(N__35791),
            .in2(_gnd_net_),
            .in3(N__30322),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_10_17_5  (
            .in0(N__38527),
            .in1(N__35482),
            .in2(_gnd_net_),
            .in3(N__30248),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_10_17_7  (
            .in0(N__38526),
            .in1(N__35182),
            .in2(_gnd_net_),
            .in3(N__30100),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_0 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_10_18_0  (
            .in0(N__30581),
            .in1(N__33935),
            .in2(N__35654),
            .in3(N__34244),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_18_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_10_18_1  (
            .in0(N__34243),
            .in1(N__35744),
            .in2(N__33983),
            .in3(N__30371),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_10_18_2  (
            .in0(N__38530),
            .in1(N__35131),
            .in2(_gnd_net_),
            .in3(N__30066),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_18_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_10_18_3  (
            .in0(N__34241),
            .in1(N__35274),
            .in2(N__33982),
            .in3(N__32931),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_4 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_10_18_4  (
            .in0(N__30287),
            .in1(N__34240),
            .in2(_gnd_net_),
            .in3(N__35567),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_10_18_5  (
            .in0(N__35690),
            .in1(N__38532),
            .in2(_gnd_net_),
            .in3(N__33350),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_18_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_10_18_6  (
            .in0(N__30414),
            .in1(N__33931),
            .in2(N__35538),
            .in3(N__34242),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_10_18_7  (
            .in0(N__35431),
            .in1(N__38531),
            .in2(_gnd_net_),
            .in3(N__30181),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_0 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_10_19_0  (
            .in0(N__33285),
            .in1(N__33941),
            .in2(N__35882),
            .in3(N__34320),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_19_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_10_19_1  (
            .in0(N__34318),
            .in1(N__37982),
            .in2(N__33985),
            .in3(N__37944),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_10_19_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_10_19_2  (
            .in0(N__26784),
            .in1(N__26775),
            .in2(_gnd_net_),
            .in3(N__34716),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_3 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_10_19_3  (
            .in0(N__33937),
            .in1(N__35843),
            .in2(N__34341),
            .in3(N__33087),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_19_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_10_19_4  (
            .in0(N__26763),
            .in1(N__26754),
            .in2(_gnd_net_),
            .in3(N__34717),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_19_5 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_10_19_5  (
            .in0(N__34324),
            .in1(N__35694),
            .in2(N__33357),
            .in3(N__33945),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_19_6 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_10_19_6  (
            .in0(N__35394),
            .in1(N__34319),
            .in2(N__30540),
            .in3(N__33936),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_10_19_7  (
            .in0(N__34317),
            .in1(N__38111),
            .in2(N__33984),
            .in3(N__30219),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_20_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_10_20_1  (
            .in0(N__33948),
            .in1(N__34326),
            .in2(N__35613),
            .in3(N__30896),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_20_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_10_20_2  (
            .in0(N__34327),
            .in1(N__33946),
            .in2(N__36126),
            .in3(N__31113),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_10_20_3  (
            .in0(N__34704),
            .in1(N__26865),
            .in2(_gnd_net_),
            .in3(N__26859),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_10_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_10_20_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_10_20_4  (
            .in0(N__26850),
            .in1(N__26838),
            .in2(_gnd_net_),
            .in3(N__34702),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_10_20_5  (
            .in0(N__34705),
            .in1(N__26832),
            .in2(_gnd_net_),
            .in3(N__26823),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_20_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_10_20_6  (
            .in0(N__34325),
            .in1(N__33947),
            .in2(N__35658),
            .in3(N__30582),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_10_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_10_20_7 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_10_20_7  (
            .in0(N__34703),
            .in1(_gnd_net_),
            .in2(N__27033),
            .in3(N__27021),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_0 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_10_21_0  (
            .in0(N__33987),
            .in1(N__34329),
            .in2(N__30792),
            .in3(N__36077),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_10_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_10_21_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_10_21_1  (
            .in0(N__34328),
            .in1(N__33988),
            .in2(N__30903),
            .in3(N__35612),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_11_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_11_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_11_5_0  (
            .in0(_gnd_net_),
            .in1(N__26997),
            .in2(N__26991),
            .in3(N__29008),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_11_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_11_5_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_11_5_1  (
            .in0(N__28977),
            .in1(N__26982),
            .in2(N__26976),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_11_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_11_5_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_11_5_2  (
            .in0(N__28941),
            .in1(N__26967),
            .in2(N__26958),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_11_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_11_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__26949),
            .in2(N__26943),
            .in3(N__28923),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_11_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_11_5_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_11_5_4  (
            .in0(N__28905),
            .in1(N__26934),
            .in2(N__26928),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_11_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_11_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__27180),
            .in2(N__27168),
            .in3(N__29277),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_11_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_11_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(N__27159),
            .in2(N__28740),
            .in3(N__29256),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_11_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_11_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__27153),
            .in2(N__27144),
            .in3(N__29235),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_11_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_11_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__27135),
            .in2(N__27123),
            .in3(N__29214),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_11_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_11_6_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_11_6_1  (
            .in0(N__29196),
            .in1(N__27111),
            .in2(N__27099),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_11_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_11_6_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_11_6_2  (
            .in0(N__29178),
            .in1(N__27090),
            .in2(N__27078),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_11_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_11_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__27069),
            .in2(N__27060),
            .in3(N__29160),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_11_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_11_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__27051),
            .in2(N__27042),
            .in3(N__29142),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_11_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_11_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__27252),
            .in2(N__27246),
            .in3(N__29445),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_11_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_11_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_11_6_6  (
            .in0(_gnd_net_),
            .in1(N__27234),
            .in2(N__27228),
            .in3(N__29427),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_11_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_11_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__31638),
            .in2(N__31566),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_11_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_11_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__28731),
            .in2(N__28725),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_11_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_11_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__27219),
            .in2(N__27210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_11_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_11_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__27201),
            .in2(N__27189),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_11_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_11_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__29091),
            .in2(N__28887),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_11_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_11_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__29019),
            .in2(N__28716),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_11_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_11_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__27408),
            .in2(N__27387),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_11_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_11_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__27375),
            .in2(N__27351),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.un4_running_cry_30_THRU_LUT4_0_LC_11_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.un4_running_cry_30_THRU_LUT4_0_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.un4_running_cry_30_THRU_LUT4_0_LC_11_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.un4_running_cry_30_THRU_LUT4_0_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27411),
            .lcout(\phase_controller_inst2.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_11_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_11_8_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_11_8_0  (
            .in0(N__29511),
            .in1(N__27398),
            .in2(N__29490),
            .in3(N__31347),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_11_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_11_8_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_11_8_1  (
            .in0(N__31346),
            .in1(N__29489),
            .in2(N__27402),
            .in3(N__29510),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_11_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_11_8_5 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_11_8_5  (
            .in0(N__27278),
            .in1(N__29846),
            .in2(N__27369),
            .in3(N__29465),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_11_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_11_8_6 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_11_8_6  (
            .in0(N__29466),
            .in1(N__27365),
            .in2(N__29847),
            .in3(N__27279),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_11_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_11_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_30_LC_11_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_30_LC_11_8_7  (
            .in0(N__27342),
            .in1(N__27321),
            .in2(_gnd_net_),
            .in3(N__32640),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50839),
            .ce(N__31698),
            .sr(N__50285));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__27270),
            .in2(N__27261),
            .in3(N__27703),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__27561),
            .in2(N__27549),
            .in3(N__28011),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__27540),
            .in2(N__27531),
            .in3(N__27978),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__27522),
            .in2(N__27516),
            .in3(N__27960),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__27507),
            .in2(N__27495),
            .in3(N__27942),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_11_9_5  (
            .in0(N__27924),
            .in1(N__27486),
            .in2(N__27477),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__27465),
            .in2(N__27456),
            .in3(N__27906),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__27447),
            .in2(N__27438),
            .in3(N__27888),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__27429),
            .in2(N__27420),
            .in3(N__27870),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__27687),
            .in2(N__27675),
            .in3(N__28173),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__27666),
            .in2(N__27654),
            .in3(N__28155),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_10_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_11_10_3  (
            .in0(N__28137),
            .in1(N__27645),
            .in2(N__27636),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_11_10_4  (
            .in0(N__28119),
            .in1(N__27627),
            .in2(N__27615),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_11_10_5  (
            .in0(N__28101),
            .in1(N__32706),
            .in2(N__27603),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_11_10_6  (
            .in0(N__28083),
            .in1(N__27582),
            .in2(N__27594),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(N__27576),
            .in2(N__27570),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__31491),
            .in2(N__31551),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__27852),
            .in2(N__27840),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__27825),
            .in2(N__27813),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__27798),
            .in2(N__27789),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__27777),
            .in2(N__27771),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__27762),
            .in2(N__27756),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__27744),
            .in2(N__27738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.un4_running_cry_30_THRU_LUT4_0_LC_11_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.un4_running_cry_30_THRU_LUT4_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.un4_running_cry_30_THRU_LUT4_0_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.un4_running_cry_30_THRU_LUT4_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27729),
            .lcout(\phase_controller_inst1.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_11_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_11_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_11_12_0  (
            .in0(N__27717),
            .in1(N__27708),
            .in2(N__27992),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.N_42_i ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_11_12_1  (
            .in0(N__32104),
            .in1(N__28010),
            .in2(_gnd_net_),
            .in3(N__27996),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_12_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_11_12_2  (
            .in0(N__32108),
            .in1(N__27977),
            .in2(N__27993),
            .in3(N__27963),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_11_12_3  (
            .in0(N__32105),
            .in1(N__27959),
            .in2(_gnd_net_),
            .in3(N__27945),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_11_12_4  (
            .in0(N__32109),
            .in1(N__27941),
            .in2(_gnd_net_),
            .in3(N__27927),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_11_12_5  (
            .in0(N__32106),
            .in1(N__27923),
            .in2(_gnd_net_),
            .in3(N__27909),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_11_12_6  (
            .in0(N__32110),
            .in1(N__27905),
            .in2(_gnd_net_),
            .in3(N__27891),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_11_12_7  (
            .in0(N__32107),
            .in1(N__27887),
            .in2(_gnd_net_),
            .in3(N__27873),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__50799),
            .ce(),
            .sr(N__50318));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_11_13_0  (
            .in0(N__32087),
            .in1(N__27869),
            .in2(_gnd_net_),
            .in3(N__27855),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_11_13_1  (
            .in0(N__32111),
            .in1(N__28172),
            .in2(_gnd_net_),
            .in3(N__28158),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_11_13_2  (
            .in0(N__32084),
            .in1(N__28154),
            .in2(_gnd_net_),
            .in3(N__28140),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_11_13_3  (
            .in0(N__32112),
            .in1(N__28136),
            .in2(_gnd_net_),
            .in3(N__28122),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_11_13_4  (
            .in0(N__32085),
            .in1(N__28118),
            .in2(_gnd_net_),
            .in3(N__28104),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_11_13_5  (
            .in0(N__32113),
            .in1(N__28100),
            .in2(_gnd_net_),
            .in3(N__28086),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_11_13_6  (
            .in0(N__32086),
            .in1(N__28082),
            .in2(_gnd_net_),
            .in3(N__28068),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_11_13_7  (
            .in0(N__32114),
            .in1(N__28052),
            .in2(_gnd_net_),
            .in3(N__28038),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__50790),
            .ce(),
            .sr(N__50326));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_11_14_0  (
            .in0(N__32115),
            .in1(N__28028),
            .in2(_gnd_net_),
            .in3(N__28014),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_11_14_1  (
            .in0(N__32144),
            .in1(N__31505),
            .in2(_gnd_net_),
            .in3(N__28356),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_11_14_2  (
            .in0(N__32116),
            .in1(N__31529),
            .in2(_gnd_net_),
            .in3(N__28353),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_11_14_3  (
            .in0(N__32145),
            .in1(N__28340),
            .in2(_gnd_net_),
            .in3(N__28326),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_11_14_4  (
            .in0(N__32117),
            .in1(N__28316),
            .in2(_gnd_net_),
            .in3(N__28302),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_11_14_5  (
            .in0(N__32146),
            .in1(N__28289),
            .in2(_gnd_net_),
            .in3(N__28275),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_11_14_6  (
            .in0(N__32118),
            .in1(N__28265),
            .in2(_gnd_net_),
            .in3(N__28251),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_11_14_7  (
            .in0(N__32147),
            .in1(N__28235),
            .in2(_gnd_net_),
            .in3(N__28221),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__50781),
            .ce(),
            .sr(N__50334));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_11_15_0  (
            .in0(N__32140),
            .in1(N__28211),
            .in2(_gnd_net_),
            .in3(N__28197),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_11_15_1  (
            .in0(N__32148),
            .in1(N__28192),
            .in2(_gnd_net_),
            .in3(N__28176),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_11_15_2  (
            .in0(N__32141),
            .in1(N__28487),
            .in2(_gnd_net_),
            .in3(N__28473),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_11_15_3  (
            .in0(N__32149),
            .in1(N__28463),
            .in2(_gnd_net_),
            .in3(N__28449),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_11_15_4  (
            .in0(N__32142),
            .in1(N__28439),
            .in2(_gnd_net_),
            .in3(N__28425),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_11_15_5  (
            .in0(N__32150),
            .in1(N__28417),
            .in2(_gnd_net_),
            .in3(N__28398),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_11_15_6  (
            .in0(N__32143),
            .in1(N__28384),
            .in2(_gnd_net_),
            .in3(N__28395),
            .lcout(\phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50775),
            .ce(),
            .sr(N__50343));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_11_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_11_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(N__28681),
            .in2(N__31838),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_11_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_11_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__49666),
            .in2(N__29745),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_11_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_11_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__28362),
            .in2(N__49769),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_11_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_11_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(N__49670),
            .in2(N__32952),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_11_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_11_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__32901),
            .in2(N__49770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_11_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_11_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__49674),
            .in2(N__28536),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_11_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_11_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__28524),
            .in2(N__49771),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_11_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_11_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__49678),
            .in2(N__38544),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_11_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(N__49691),
            .in2(N__28518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_11_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_11_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(N__31884),
            .in2(N__49775),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_11_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_11_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(N__49679),
            .in2(N__28509),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_11_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_11_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__37995),
            .in2(N__49772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_11_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_11_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__49683),
            .in2(N__30381),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_11_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_11_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__28557),
            .in2(N__49773),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_11_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_11_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__49687),
            .in2(N__28551),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_11_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_11_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__38319),
            .in2(N__49774),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_11_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_11_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__28542),
            .in2(N__49776),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_11_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_11_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__49698),
            .in2(N__37908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_11_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_11_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__30507),
            .in2(N__49777),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_11_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_11_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__49702),
            .in2(N__33114),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_11_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_11_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__33258),
            .in2(N__49778),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_11_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_11_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__49706),
            .in2(N__33060),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_11_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_11_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__28578),
            .in2(N__49779),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_11_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_11_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__49710),
            .in2(N__30342),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_11_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_11_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__28572),
            .in2(N__49780),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_11_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_11_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__49714),
            .in2(N__30552),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_11_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_11_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__30870),
            .in2(N__49781),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_11_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_11_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__49718),
            .in2(N__28566),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_11_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_11_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__31083),
            .in2(N__49782),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_11_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_11_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__49722),
            .in2(N__30753),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_11_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_11_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__29730),
            .in2(N__49783),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_11_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_11_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__34340),
            .in2(_gnd_net_),
            .in3(N__28707),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_11_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_11_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_11_20_0  (
            .in0(N__42836),
            .in1(N__42977),
            .in2(N__46839),
            .in3(N__42236),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_11_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_11_20_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_11_20_1  (
            .in0(N__28701),
            .in1(N__38133),
            .in2(N__28704),
            .in3(N__31323),
            .lcout(\current_shift_inst.PI_CTRL.N_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_11_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_11_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_11_20_7  (
            .in0(N__42905),
            .in1(N__46235),
            .in2(N__43865),
            .in3(N__42308),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_21_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_11_21_5  (
            .in0(N__28695),
            .in1(N__34337),
            .in2(N__33986),
            .in3(N__30605),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_23_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_23_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_11_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31289),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31269),
            .ce(),
            .sr(N__50382));
    defparam \phase_controller_inst2.S2_LC_11_27_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_11_27_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_11_27_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.S2_LC_11_27_0  (
            .in0(N__37416),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50751),
            .ce(N__43676),
            .sr(N__50392));
    defparam \phase_controller_inst2.stoper_hc.m10_1_LC_12_3_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m10_1_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m10_1_LC_12_3_2 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \phase_controller_inst2.stoper_hc.m10_1_LC_12_3_2  (
            .in0(N__34859),
            .in1(N__37387),
            .in2(_gnd_net_),
            .in3(N__31470),
            .lcout(\phase_controller_inst2.stoper_hc.m10Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.m3_LC_12_3_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m3_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m3_LC_12_3_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.m3_LC_12_3_6  (
            .in0(N__44126),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31469),
            .lcout(\phase_controller_inst2.m3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_2_LC_12_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_12_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_12_4_6 .LUT_INIT=16'b0100000011101010;
    LogicCell40 \phase_controller_inst2.state_2_LC_12_4_6  (
            .in0(N__37388),
            .in1(N__41862),
            .in2(N__34812),
            .in3(N__34863),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50871),
            .ce(N__43628),
            .sr(N__50248));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_5_3 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_5_3  (
            .in0(N__29954),
            .in1(N__28992),
            .in2(_gnd_net_),
            .in3(N__29012),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50859),
            .ce(),
            .sr(N__50253));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_12_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_12_6_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_12_6_1  (
            .in0(N__29120),
            .in1(N__29585),
            .in2(N__29613),
            .in3(N__29102),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_12_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_12_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_25_LC_12_6_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_25_LC_12_6_3  (
            .in0(N__28877),
            .in1(N__32692),
            .in2(_gnd_net_),
            .in3(N__28851),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50848),
            .ce(N__31693),
            .sr(N__50263));
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_12_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_12_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_7_LC_12_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_7_LC_12_6_7  (
            .in0(N__28802),
            .in1(N__32691),
            .in2(_gnd_net_),
            .in3(N__28779),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50848),
            .ce(N__31693),
            .sr(N__50263));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_12_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_12_7_0 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_12_7_0  (
            .in0(N__31427),
            .in1(N__29373),
            .in2(N__29400),
            .in3(N__31418),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_12_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_12_7_1 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_12_7_1  (
            .in0(N__29372),
            .in1(N__31428),
            .in2(N__31419),
            .in3(N__29399),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_7_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_12_7_2  (
            .in0(N__29036),
            .in1(N__29537),
            .in2(N__29052),
            .in3(N__29559),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_12_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_12_7_4 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_12_7_4  (
            .in0(N__29121),
            .in1(N__29612),
            .in2(N__29586),
            .in3(N__29103),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.m3_LC_12_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m3_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m3_LC_12_7_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.m3_LC_12_7_5  (
            .in0(N__29085),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31221),
            .lcout(\phase_controller_inst1.m3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.m37_LC_12_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m37_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m37_LC_12_7_6 .LUT_INIT=16'b0111010111110101;
    LogicCell40 \phase_controller_inst2.stoper_hc.m37_LC_12_7_6  (
            .in0(N__31471),
            .in1(N__44081),
            .in2(N__44137),
            .in3(N__31439),
            .lcout(\phase_controller_inst2.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_12_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_12_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_12_7_7 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_12_7_7  (
            .in0(N__29558),
            .in1(N__29048),
            .in2(N__29538),
            .in3(N__29037),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_12_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_12_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_c_inv_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(N__29013),
            .in2(N__28955),
            .in3(N__28988),
            .lcout(\phase_controller_inst2.stoper_tr.N_38_i ),
            .ltout(),
            .carryin(bfn_12_8_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_12_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_12_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_12_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_12_8_1  (
            .in0(N__29943),
            .in1(N__28973),
            .in2(_gnd_net_),
            .in3(N__28959),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_12_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_12_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_12_8_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_12_8_2  (
            .in0(N__29947),
            .in1(N__28940),
            .in2(N__28956),
            .in3(N__28926),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_12_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_12_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_12_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_12_8_3  (
            .in0(N__29944),
            .in1(N__28922),
            .in2(_gnd_net_),
            .in3(N__28908),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_12_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_12_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_12_8_4  (
            .in0(N__29948),
            .in1(N__28904),
            .in2(_gnd_net_),
            .in3(N__28890),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_12_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_12_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_12_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_12_8_5  (
            .in0(N__29945),
            .in1(N__29273),
            .in2(_gnd_net_),
            .in3(N__29259),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_12_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_12_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_12_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_12_8_6  (
            .in0(N__29949),
            .in1(N__29252),
            .in2(_gnd_net_),
            .in3(N__29238),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_12_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_12_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_12_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_12_8_7  (
            .in0(N__29946),
            .in1(N__29231),
            .in2(_gnd_net_),
            .in3(N__29217),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7 ),
            .clk(N__50825),
            .ce(),
            .sr(N__50276));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_12_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_12_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_12_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_12_9_0  (
            .in0(N__29953),
            .in1(N__29213),
            .in2(_gnd_net_),
            .in3(N__29199),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_12_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_12_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_12_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_12_9_1  (
            .in0(N__29980),
            .in1(N__29195),
            .in2(_gnd_net_),
            .in3(N__29181),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_12_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_12_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_12_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_12_9_2  (
            .in0(N__29950),
            .in1(N__29177),
            .in2(_gnd_net_),
            .in3(N__29163),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_12_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_12_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_12_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_12_9_3  (
            .in0(N__29981),
            .in1(N__29159),
            .in2(_gnd_net_),
            .in3(N__29145),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_12_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_12_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_12_9_4  (
            .in0(N__29951),
            .in1(N__29138),
            .in2(_gnd_net_),
            .in3(N__29124),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_12_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_12_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_12_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_12_9_5  (
            .in0(N__29982),
            .in1(N__29444),
            .in2(_gnd_net_),
            .in3(N__29430),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_12_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_12_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_12_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_12_9_6  (
            .in0(N__29952),
            .in1(N__29423),
            .in2(_gnd_net_),
            .in3(N__29409),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_12_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_12_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_12_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_12_9_7  (
            .in0(N__29983),
            .in1(N__31598),
            .in2(_gnd_net_),
            .in3(N__29406),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15 ),
            .clk(N__50815),
            .ce(),
            .sr(N__50286));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_12_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_12_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_12_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_12_10_0  (
            .in0(N__29984),
            .in1(N__31616),
            .in2(_gnd_net_),
            .in3(N__29403),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_12_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_12_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_12_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_12_10_1  (
            .in0(N__29988),
            .in1(N__29390),
            .in2(_gnd_net_),
            .in3(N__29376),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_12_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_12_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_12_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_12_10_2  (
            .in0(N__29985),
            .in1(N__29371),
            .in2(_gnd_net_),
            .in3(N__29355),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_12_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_12_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_12_10_3  (
            .in0(N__29989),
            .in1(N__29345),
            .in2(_gnd_net_),
            .in3(N__29331),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_12_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_12_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_12_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_12_10_4  (
            .in0(N__29986),
            .in1(N__29318),
            .in2(_gnd_net_),
            .in3(N__29304),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_12_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_12_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_12_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_12_10_5  (
            .in0(N__29990),
            .in1(N__29294),
            .in2(_gnd_net_),
            .in3(N__29280),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_12_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_12_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_12_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_12_10_6  (
            .in0(N__29987),
            .in1(N__29630),
            .in2(_gnd_net_),
            .in3(N__29616),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_12_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_12_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_12_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_12_10_7  (
            .in0(N__29991),
            .in1(N__29608),
            .in2(_gnd_net_),
            .in3(N__29589),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23 ),
            .clk(N__50806),
            .ce(),
            .sr(N__50295));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_12_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_12_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_12_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_12_11_0  (
            .in0(N__29955),
            .in1(N__29581),
            .in2(_gnd_net_),
            .in3(N__29562),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_12_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_12_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_12_11_1  (
            .in0(N__29959),
            .in1(N__29557),
            .in2(_gnd_net_),
            .in3(N__29541),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_12_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_12_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_12_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_12_11_2  (
            .in0(N__29956),
            .in1(N__29528),
            .in2(_gnd_net_),
            .in3(N__29514),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_12_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_12_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_12_11_3  (
            .in0(N__29960),
            .in1(N__29509),
            .in2(_gnd_net_),
            .in3(N__29493),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_12_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_12_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_12_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_12_11_4  (
            .in0(N__29957),
            .in1(N__29485),
            .in2(_gnd_net_),
            .in3(N__29469),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_12_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_12_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_12_11_5  (
            .in0(N__29961),
            .in1(N__29464),
            .in2(_gnd_net_),
            .in3(N__29448),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29 ),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_12_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_12_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_12_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_12_11_6  (
            .in0(N__29958),
            .in1(N__29837),
            .in2(_gnd_net_),
            .in3(N__29850),
            .lcout(\phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50798),
            .ce(),
            .sr(N__50302));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39783),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50789),
            .ce(N__36197),
            .sr(N__50310));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29760),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_12_3 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_12_12_3  (
            .in0(N__29702),
            .in1(N__34330),
            .in2(N__29768),
            .in3(N__29823),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_12_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_12_12_4  (
            .in0(N__38432),
            .in1(N__29701),
            .in2(_gnd_net_),
            .in3(N__29761),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__34331),
            .in2(_gnd_net_),
            .in3(N__30598),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_12_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_12_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__29718),
            .in2(N__31865),
            .in3(N__31861),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_12_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_12_13_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33033),
            .in3(N__29649),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_12_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_12_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__32937),
            .in2(_gnd_net_),
            .in3(N__29646),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_12_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_12_13_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32883),
            .in3(N__30141),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_12_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_12_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__32889),
            .in2(_gnd_net_),
            .in3(N__30105),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_12_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_12_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__33045),
            .in2(_gnd_net_),
            .in3(N__30072),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_12_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_12_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__34947),
            .in2(_gnd_net_),
            .in3(N__30069),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_12_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_12_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__32847),
            .in2(_gnd_net_),
            .in3(N__30033),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_12_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_12_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__33039),
            .in2(_gnd_net_),
            .in3(N__30030),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_12_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_12_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__33156),
            .in2(_gnd_net_),
            .in3(N__29997),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_12_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_12_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__33195),
            .in2(_gnd_net_),
            .in3(N__29994),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_12_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_12_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__33099),
            .in2(_gnd_net_),
            .in3(N__30252),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_12_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_12_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__33093),
            .in2(_gnd_net_),
            .in3(N__30222),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_12_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_12_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__38073),
            .in2(_gnd_net_),
            .in3(N__30189),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_12_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_12_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__38121),
            .in2(_gnd_net_),
            .in3(N__30186),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_12_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_12_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__33024),
            .in2(_gnd_net_),
            .in3(N__30156),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_12_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_12_15_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33183),
            .in3(N__30153),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_12_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_12_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__33162),
            .in2(_gnd_net_),
            .in3(N__30150),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_12_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_12_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__33168),
            .in2(_gnd_net_),
            .in3(N__30147),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_12_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_12_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__33150),
            .in2(_gnd_net_),
            .in3(N__30144),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_12_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_12_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__33174),
            .in2(_gnd_net_),
            .in3(N__30333),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_12_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_12_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__33246),
            .in2(_gnd_net_),
            .in3(N__30303),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_12_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_12_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__33303),
            .in2(_gnd_net_),
            .in3(N__30300),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_12_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_12_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__33189),
            .in2(_gnd_net_),
            .in3(N__30297),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_12_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_12_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__33297),
            .in2(_gnd_net_),
            .in3(N__30294),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_12_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_12_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__33144),
            .in2(_gnd_net_),
            .in3(N__30291),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_12_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_12_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__33291),
            .in2(_gnd_net_),
            .in3(N__30261),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_12_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_12_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__36090),
            .in2(_gnd_net_),
            .in3(N__30258),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_12_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_12_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__30255),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_12_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_12_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30615),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_12_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_12_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_12_16_6  (
            .in0(N__34225),
            .in1(N__35641),
            .in2(_gnd_net_),
            .in3(N__30568),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_12_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_12_16_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_12_16_7  (
            .in0(N__38524),
            .in1(N__35386),
            .in2(_gnd_net_),
            .in3(N__30523),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_17_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_12_17_0  (
            .in0(N__30498),
            .in1(N__30486),
            .in2(_gnd_net_),
            .in3(N__34726),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_17_1 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_17_1  (
            .in0(N__34727),
            .in1(N__30477),
            .in2(_gnd_net_),
            .in3(N__30468),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_17_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_12_17_2  (
            .in0(N__30456),
            .in1(N__30444),
            .in2(_gnd_net_),
            .in3(N__34728),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_17_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_12_17_3  (
            .in0(N__34729),
            .in1(N__30435),
            .in2(_gnd_net_),
            .in3(N__30423),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_12_17_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_12_17_4  (
            .in0(N__38522),
            .in1(N__35527),
            .in2(_gnd_net_),
            .in3(N__30406),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_12_17_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_12_17_5  (
            .in0(N__35737),
            .in1(N__38523),
            .in2(_gnd_net_),
            .in3(N__30364),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_17_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_17_6  (
            .in0(N__30816),
            .in1(N__30804),
            .in2(_gnd_net_),
            .in3(N__34730),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_12_17_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_12_17_7  (
            .in0(N__36067),
            .in1(N__34314),
            .in2(_gnd_net_),
            .in3(N__30769),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_18_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_18_0  (
            .in0(N__34699),
            .in1(N__30741),
            .in2(_gnd_net_),
            .in3(N__30732),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_12_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_12_18_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_12_18_1  (
            .in0(N__30720),
            .in1(N__30711),
            .in2(_gnd_net_),
            .in3(N__34697),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_12_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_12_18_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30699),
            .in3(N__33233),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50765),
            .ce(),
            .sr(N__50355));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_12_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_12_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34698),
            .lcout(\current_shift_inst.N_1275_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_18_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_18_6  (
            .in0(N__34700),
            .in1(N__30660),
            .in2(_gnd_net_),
            .in3(N__30648),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_18_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_18_7  (
            .in0(N__30636),
            .in1(N__30627),
            .in2(_gnd_net_),
            .in3(N__34701),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_19_0 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_19_0  (
            .in0(N__34708),
            .in1(N__31047),
            .in2(_gnd_net_),
            .in3(N__31035),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_19_1 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_19_1  (
            .in0(N__31023),
            .in1(N__31011),
            .in2(_gnd_net_),
            .in3(N__34709),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_19_2 .LUT_INIT=16'b0000010110101111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_19_2  (
            .in0(N__34710),
            .in1(_gnd_net_),
            .in2(N__30999),
            .in3(N__30984),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_19_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_19_3  (
            .in0(N__30969),
            .in1(N__30960),
            .in2(_gnd_net_),
            .in3(N__34711),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_12_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_12_19_4 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_12_19_4  (
            .in0(N__34712),
            .in1(N__30948),
            .in2(_gnd_net_),
            .in3(N__30936),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_12_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_12_19_5 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_12_19_5  (
            .in0(N__30924),
            .in1(N__30912),
            .in2(_gnd_net_),
            .in3(N__34707),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_12_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_12_19_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_12_19_6  (
            .in0(N__34312),
            .in1(N__35602),
            .in2(_gnd_net_),
            .in3(N__30889),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_12_19_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_12_19_7  (
            .in0(N__30861),
            .in1(N__30849),
            .in2(_gnd_net_),
            .in3(N__34706),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_20_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_12_20_0  (
            .in0(N__30840),
            .in1(N__30828),
            .in2(_gnd_net_),
            .in3(N__34719),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_20_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_12_20_1  (
            .in0(N__34720),
            .in1(N__31182),
            .in2(_gnd_net_),
            .in3(N__31170),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_20_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_20_2  (
            .in0(N__31158),
            .in1(N__31146),
            .in2(_gnd_net_),
            .in3(N__34718),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_20_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_20_3  (
            .in0(N__34721),
            .in1(N__31134),
            .in2(_gnd_net_),
            .in3(N__31122),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_12_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_12_20_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_12_20_5  (
            .in0(N__36121),
            .in1(N__34313),
            .in2(_gnd_net_),
            .in3(N__31108),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34722),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_21_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_21_1  (
            .in0(N__31071),
            .in1(N__31062),
            .in2(_gnd_net_),
            .in3(N__34740),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_12_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_12_21_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_12_21_2  (
            .in0(N__43514),
            .in1(N__42719),
            .in2(N__43358),
            .in3(N__42772),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_12_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_12_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_12_21_3  (
            .in0(N__43915),
            .in1(N__43978),
            .in2(N__43802),
            .in3(N__43165),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_12_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_12_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_12_21_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_12_21_4  (
            .in0(N__43231),
            .in1(N__43466),
            .in2(N__31050),
            .in3(N__31317),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_12_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_12_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_12_21_5  (
            .in0(N__43282),
            .in1(N__46585),
            .in2(N__31332),
            .in3(N__31329),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_12_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_12_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_12_22_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__43106),
            .in2(_gnd_net_),
            .in3(N__43402),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_tr_LC_12_23_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_23_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_12_23_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31288),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__31268),
            .ce(),
            .sr(N__50378));
    defparam \phase_controller_inst2.S1_LC_12_26_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_12_26_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_12_26_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_12_26_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41918),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50750),
            .ce(N__43663),
            .sr(N__50387));
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_4.C_ON=1'b0;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_4 (
            .in0(N__50415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_red_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_0_LC_13_2_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_0_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_0_LC_13_2_0 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_0_LC_13_2_0  (
            .in0(N__37463),
            .in1(N__37533),
            .in2(N__38845),
            .in3(N__40642),
            .lcout(\phase_controller_inst1.stoper_hc.m19_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_1_LC_13_3_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_1_LC_13_3_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_1_LC_13_3_7 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_er_RNISS5N_1_LC_13_3_7  (
            .in0(N__37472),
            .in1(N__37534),
            .in2(N__38856),
            .in3(N__40635),
            .lcout(\phase_controller_inst1.stoper_hc.m34_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_tr_LC_13_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_13_4_2 .LUT_INIT=16'b0111000001110111;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_13_4_2  (
            .in0(N__37584),
            .in1(N__34933),
            .in2(N__31213),
            .in3(N__31230),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50882),
            .ce(N__43627),
            .sr(N__50244));
    defparam \phase_controller_inst2.start_timer_tr_LC_13_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_13_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_13_4_4 .LUT_INIT=16'b0010101000111111;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_13_4_4  (
            .in0(N__42152),
            .in1(N__34906),
            .in2(N__44208),
            .in3(N__31188),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50882),
            .ce(N__43627),
            .sr(N__50244));
    defparam \phase_controller_inst2.state_1_LC_13_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_13_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_13_4_6 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \phase_controller_inst2.state_1_LC_13_4_6  (
            .in0(N__34878),
            .in1(N__34864),
            .in2(N__37401),
            .in3(N__34907),
            .lcout(\phase_controller_inst2.N_139_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50882),
            .ce(N__43627),
            .sr(N__50244));
    defparam \phase_controller_inst2.stoper_hc.m20_ns_1_LC_13_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m20_ns_1_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m20_ns_1_LC_13_5_7 .LUT_INIT=16'b0000001110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.m20_ns_1_LC_13_5_7  (
            .in0(N__42115),
            .in1(N__41908),
            .in2(N__44204),
            .in3(N__34904),
            .lcout(\phase_controller_inst2.stoper_hc.m20_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_13_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_13_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_28_LC_13_6_0 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_28_LC_13_6_0  (
            .in0(N__34995),
            .in1(N__48171),
            .in2(N__51520),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50861),
            .ce(N__49248),
            .sr(N__50254));
    defparam \phase_controller_inst2.stoper_hc.m38_LC_13_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m38_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m38_LC_13_7_2 .LUT_INIT=16'b1111010101110101;
    LogicCell40 \phase_controller_inst2.stoper_hc.m38_LC_13_7_2  (
            .in0(N__31472),
            .in1(N__44082),
            .in2(N__44144),
            .in3(N__31443),
            .lcout(\phase_controller_inst2.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_13_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_13_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_13_7_4  (
            .in0(N__32669),
            .in1(N__32252),
            .in2(_gnd_net_),
            .in3(N__32232),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_7_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_13_7_5  (
            .in0(N__32767),
            .in1(N__32748),
            .in2(_gnd_net_),
            .in3(N__32668),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_13_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_18_LC_13_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_18_LC_13_8_2  (
            .in0(N__32248),
            .in1(N__32231),
            .in2(_gnd_net_),
            .in3(N__32563),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50840),
            .ce(N__31699),
            .sr(N__50270));
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_19_LC_13_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_19_LC_13_8_4  (
            .in0(N__32821),
            .in1(N__32562),
            .in2(_gnd_net_),
            .in3(N__32841),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50840),
            .ce(N__31699),
            .sr(N__50270));
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_13_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_28_LC_13_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_28_LC_13_9_4  (
            .in0(N__32689),
            .in1(N__31407),
            .in2(_gnd_net_),
            .in3(N__31365),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50827),
            .ce(N__31701),
            .sr(N__50277));
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_16_LC_13_9_5  (
            .in0(N__31815),
            .in1(N__31782),
            .in2(_gnd_net_),
            .in3(N__32690),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50827),
            .ce(N__31701),
            .sr(N__50277));
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_13_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.target_time_17_LC_13_9_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_time_17_LC_13_9_6  (
            .in0(N__32688),
            .in1(N__31767),
            .in2(_gnd_net_),
            .in3(N__31746),
            .lcout(\phase_controller_inst2.stoper_tr.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50827),
            .ce(N__31701),
            .sr(N__50277));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_10_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_10_0  (
            .in0(N__41300),
            .in1(N__41552),
            .in2(N__31650),
            .in3(N__31662),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_10_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_13_10_1  (
            .in0(N__31661),
            .in1(N__41301),
            .in2(N__41553),
            .in3(N__31646),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_13_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_29_LC_13_10_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_29_LC_13_10_3  (
            .in0(N__34973),
            .in1(_gnd_net_),
            .in2(N__51516),
            .in3(N__45057),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50817),
            .ce(N__49241),
            .sr(N__50287));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_10_4 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_13_10_4  (
            .in0(N__31594),
            .in1(N__31578),
            .in2(N__31617),
            .in3(N__31626),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_10_5 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_13_10_5  (
            .in0(N__31625),
            .in1(N__31615),
            .in2(N__31599),
            .in3(N__31577),
            .lcout(\phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_13_11_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_13_11_0  (
            .in0(N__31536),
            .in1(N__31511),
            .in2(N__32784),
            .in3(N__32187),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_13_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_13_11_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_13_11_1  (
            .in0(N__32186),
            .in1(N__31535),
            .in2(N__31515),
            .in3(N__32780),
            .lcout(\phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_13_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_13_11_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_13_11_2  (
            .in0(N__32822),
            .in1(N__32684),
            .in2(_gnd_net_),
            .in3(N__32837),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_19_LC_13_11_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_19_LC_13_11_3  (
            .in0(N__32686),
            .in1(_gnd_net_),
            .in2(N__32826),
            .in3(N__32823),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50808),
            .ce(N__32139),
            .sr(N__50296));
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_13_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_13_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_14_LC_13_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_14_LC_13_11_6  (
            .in0(N__32772),
            .in1(N__32746),
            .in2(_gnd_net_),
            .in3(N__32687),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50808),
            .ce(N__32139),
            .sr(N__50296));
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.target_time_18_LC_13_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_time_18_LC_13_11_7  (
            .in0(N__32685),
            .in1(N__32253),
            .in2(_gnd_net_),
            .in3(N__32230),
            .lcout(\phase_controller_inst1.stoper_tr.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50808),
            .ce(N__32139),
            .sr(N__50296));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__34332),
            .in2(_gnd_net_),
            .in3(N__33975),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_12_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_13_12_3  (
            .in0(N__35086),
            .in1(N__38431),
            .in2(_gnd_net_),
            .in3(N__31909),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33001),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_12_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_13_12_5  (
            .in0(N__33002),
            .in1(_gnd_net_),
            .in2(N__31842),
            .in3(N__38430),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36160),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50800),
            .ce(N__36195),
            .sr(N__50303));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39456),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50800),
            .ce(N__36195),
            .sr(N__50303));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_13_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_13_13_0  (
            .in0(N__35296),
            .in1(N__38447),
            .in2(_gnd_net_),
            .in3(N__32968),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35295),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_13_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_13_13_2  (
            .in0(N__35260),
            .in1(N__38448),
            .in2(_gnd_net_),
            .in3(N__32917),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35210),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35259),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_13_6 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_13_13_6  (
            .in0(N__32874),
            .in1(N__32862),
            .in2(_gnd_net_),
            .in3(N__34752),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35113),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_14_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_13_14_0  (
            .in0(N__38497),
            .in1(N__35917),
            .in2(_gnd_net_),
            .in3(N__33130),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35508),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35464),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.m16_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m16_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m16_LC_13_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.m16_LC_13_14_3  (
            .in0(N__34911),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42132),
            .lcout(\phase_controller_inst2.stoper_hc.mZ0Z16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_14_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_13_14_4  (
            .in0(N__38498),
            .in1(N__35833),
            .in2(_gnd_net_),
            .in3(N__33076),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_13_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_13_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35164),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35072),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35327),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35413),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38047),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_13_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_13_15_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_13_15_2  (
            .in0(N__35677),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37960),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35823),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_5  (
            .in0(N__35907),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_13_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35376),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35035),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35863),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35588),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_13_16_2  (
            .in0(N__34311),
            .in1(N__35683),
            .in2(N__33990),
            .in3(N__33343),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35718),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_13_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_13_16_4  (
            .in0(N__35632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35555),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_13_16_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_13_16_6  (
            .in0(N__35864),
            .in1(N__38525),
            .in2(_gnd_net_),
            .in3(N__33269),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35767),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_13_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_13_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__33240),
            .in2(N__33234),
            .in3(N__33232),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__33213),
            .in2(_gnd_net_),
            .in3(N__33207),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_17_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__33204),
            .in2(_gnd_net_),
            .in3(N__33198),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_17_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__34425),
            .in2(_gnd_net_),
            .in3(N__34419),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_17_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__34416),
            .in2(_gnd_net_),
            .in3(N__34410),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_17_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__34407),
            .in2(_gnd_net_),
            .in3(N__34395),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_17_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(N__34392),
            .in2(_gnd_net_),
            .in3(N__34386),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_17_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__34383),
            .in2(_gnd_net_),
            .in3(N__34371),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_18_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__34368),
            .in2(_gnd_net_),
            .in3(N__34362),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_18_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__34359),
            .in2(_gnd_net_),
            .in3(N__34353),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_18_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__34350),
            .in2(_gnd_net_),
            .in3(N__34344),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_18_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__34506),
            .in2(_gnd_net_),
            .in3(N__34500),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_18_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__34497),
            .in2(_gnd_net_),
            .in3(N__34491),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_18_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__34488),
            .in2(_gnd_net_),
            .in3(N__34482),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_13_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_13_18_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__34479),
            .in2(_gnd_net_),
            .in3(N__34473),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_13_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_13_18_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__34470),
            .in2(_gnd_net_),
            .in3(N__34464),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_13_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_13_19_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__34461),
            .in2(_gnd_net_),
            .in3(N__34452),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_13_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_13_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__34449),
            .in2(_gnd_net_),
            .in3(N__34443),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_13_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_13_19_2 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34440),
            .in3(N__34428),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_13_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_13_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__34599),
            .in2(_gnd_net_),
            .in3(N__34590),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_13_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_13_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__34587),
            .in2(_gnd_net_),
            .in3(N__34581),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__34578),
            .in2(_gnd_net_),
            .in3(N__34572),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_13_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_13_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__34569),
            .in2(_gnd_net_),
            .in3(N__34563),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_13_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_13_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__34560),
            .in2(_gnd_net_),
            .in3(N__34554),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_20_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__34551),
            .in2(_gnd_net_),
            .in3(N__34542),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__34539),
            .in2(_gnd_net_),
            .in3(N__34533),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_13_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_13_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__34530),
            .in2(_gnd_net_),
            .in3(N__34521),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_13_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_13_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__34518),
            .in2(_gnd_net_),
            .in3(N__34509),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_13_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_13_20_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__34773),
            .in2(_gnd_net_),
            .in3(N__34764),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_13_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_13_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_13_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__34761),
            .in2(_gnd_net_),
            .in3(N__34755),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_13_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_13_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__34751),
            .in2(_gnd_net_),
            .in3(N__34602),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_13_21_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_13_21_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_13_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_13_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42018),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50758),
            .ce(),
            .sr(N__50365));
    defparam \phase_controller_inst2.stoper_hc.running_LC_13_21_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_13_21_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_13_21_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_13_21_4  (
            .in0(N__42045),
            .in1(N__42083),
            .in2(_gnd_net_),
            .in3(N__41984),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50758),
            .ce(),
            .sr(N__50365));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_13_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_13_21_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37115),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_13_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_13_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_13_22_5 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_13_22_5  (
            .in0(N__46589),
            .in1(N__46378),
            .in2(N__42402),
            .in3(N__46780),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50757),
            .ce(),
            .sr(N__50372));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_23_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_23_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_13_23_0  (
            .in0(N__42017),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42049),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNI3USR_LC_14_2_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNI3USR_LC_14_2_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNI3USR_LC_14_2_7 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_er_RNI3USR_LC_14_2_7  (
            .in0(N__34937),
            .in1(N__38832),
            .in2(N__40643),
            .in3(N__37575),
            .lcout(\phase_controller_inst1.stoper_hc.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNI61TR_LC_14_3_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNI61TR_LC_14_3_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNI61TR_LC_14_3_1 .LUT_INIT=16'b0000000110001001;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_er_RNI61TR_LC_14_3_1  (
            .in0(N__38820),
            .in1(N__38773),
            .in2(N__34938),
            .in3(N__40631),
            .lcout(\phase_controller_inst1.stoper_hc.m12_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI72V01_LC_14_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI72V01_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI72V01_LC_14_4_2 .LUT_INIT=16'b0101001100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_er_RNI72V01_LC_14_4_2  (
            .in0(N__34808),
            .in1(N__44203),
            .in2(N__41858),
            .in3(N__34905),
            .lcout(\phase_controller_inst2.stoper_hc.N_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.m21_LC_14_4_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.m21_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.m21_LC_14_4_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.m21_LC_14_4_5  (
            .in0(N__34865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41892),
            .lcout(\phase_controller_inst2.m21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI23UO1_LC_14_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI23UO1_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI23UO1_LC_14_5_3 .LUT_INIT=16'b0100000001001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_er_RNI23UO1_LC_14_5_3  (
            .in0(N__34804),
            .in1(N__41891),
            .in2(N__41857),
            .in3(N__34872),
            .lcout(\phase_controller_inst2.time_passed_er_RNI23UO1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI0D511_0_LC_14_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI0D511_0_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI0D511_0_LC_14_5_7 .LUT_INIT=16'b0001001111010011;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_er_RNI0D511_0_LC_14_5_7  (
            .in0(N__34803),
            .in1(N__37402),
            .in2(N__41856),
            .in3(N__34866),
            .lcout(\phase_controller_inst2.stoper_hc.m28_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI7HLK_LC_14_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI7HLK_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_RNI7HLK_LC_14_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_er_RNI7HLK_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__34799),
            .in2(_gnd_net_),
            .in3(N__41843),
            .lcout(\phase_controller_inst2.stoper_hc.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_LC_14_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_LC_14_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_er_LC_14_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_er_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42069),
            .lcout(\phase_controller_inst2.stoper_hc.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50862),
            .ce(N__35004),
            .sr(N__50255));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_8_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_8_0  (
            .in0(N__35016),
            .in1(N__37697),
            .in2(N__37830),
            .in3(N__37720),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_14_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_24_LC_14_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_24_LC_14_8_2  (
            .in0(N__39535),
            .in1(N__44679),
            .in2(_gnd_net_),
            .in3(N__51299),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50850),
            .ce(N__48826),
            .sr(N__50264));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_14_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_14_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_14_9_0  (
            .in0(N__51285),
            .in1(N__34974),
            .in2(_gnd_net_),
            .in3(N__45055),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_9_1 .LUT_INIT=16'b1111001101110001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_9_1  (
            .in0(N__37722),
            .in1(N__37696),
            .in2(N__37826),
            .in3(N__35015),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_14_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_14_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_14_9_2  (
            .in0(N__51284),
            .in1(N__48163),
            .in2(_gnd_net_),
            .in3(N__34994),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_sbtinv_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_sbtinv_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_sbtinv_LC_14_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_sbtinv_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41988),
            .lcout(\phase_controller_inst2.stoper_hc.N_266_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_9_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_9_7  (
            .in0(N__44678),
            .in1(N__39539),
            .in2(_gnd_net_),
            .in3(N__51283),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_28_LC_14_10_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_28_LC_14_10_2  (
            .in0(N__34990),
            .in1(N__48170),
            .in2(_gnd_net_),
            .in3(N__51300),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50828),
            .ce(N__48862),
            .sr(N__50278));
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_14_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_29_LC_14_10_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_29_LC_14_10_4  (
            .in0(N__34972),
            .in1(N__45056),
            .in2(_gnd_net_),
            .in3(N__51301),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50828),
            .ce(N__48862),
            .sr(N__50278));
    defparam \delay_measurement_inst.start_timer_hc_LC_14_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_14_11_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_14_11_1  (
            .in0(N__38272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34956),
            .ce(),
            .sr(N__50288));
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_14_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38271),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34956),
            .ce(),
            .sr(N__50288));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38592),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_14_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__39749),
            .in2(N__39455),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__39728),
            .in2(N__39782),
            .in3(N__35277),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__39750),
            .in2(N__39707),
            .in3(N__35241),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__39729),
            .in2(N__39680),
            .in3(N__35199),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__39653),
            .in2(N__39708),
            .in3(N__35148),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(N__39632),
            .in2(N__39681),
            .in3(N__35145),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__39654),
            .in2(N__39611),
            .in3(N__35097),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(N__39633),
            .in2(N__40026),
            .in3(N__35061),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50791),
            .ce(N__36194),
            .sr(N__50311));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__39989),
            .in2(N__39612),
            .in3(N__35019),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__39968),
            .in2(N__40025),
            .in3(N__35541),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__39990),
            .in2(N__39948),
            .in3(N__35490),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__39969),
            .in2(N__39920),
            .in3(N__35448),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__39947),
            .in2(N__39893),
            .in3(N__35445),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__39866),
            .in2(N__39921),
            .in3(N__35442),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__39842),
            .in2(N__39894),
            .in3(N__35400),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__39867),
            .in2(N__39815),
            .in3(N__35397),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50782),
            .ce(N__36193),
            .sr(N__50319));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__40238),
            .in2(N__39846),
            .in3(N__35358),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__40217),
            .in2(N__39816),
            .in3(N__35889),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__40239),
            .in2(N__40194),
            .in3(N__35847),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__40218),
            .in2(N__40167),
            .in3(N__35805),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__40193),
            .in2(N__40139),
            .in3(N__35751),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__40166),
            .in2(N__40112),
            .in3(N__35697),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__40082),
            .in2(N__40140),
            .in3(N__35661),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__40052),
            .in2(N__40113),
            .in3(N__35616),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50776),
            .ce(N__36192),
            .sr(N__50327));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__40406),
            .in2(N__40086),
            .in3(N__35577),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50771),
            .ce(N__36191),
            .sr(N__50335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__40382),
            .in2(N__40056),
            .in3(N__35544),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50771),
            .ce(N__36191),
            .sr(N__50335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__40362),
            .in2(N__40410),
            .in3(N__36204),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50771),
            .ce(N__36191),
            .sr(N__50335));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__40383),
            .in2(N__40341),
            .in3(N__36201),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50771),
            .ce(N__36191),
            .sr(N__50335));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36168),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36103),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36058),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_14_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__36027),
            .in2(_gnd_net_),
            .in3(N__36033),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_14_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__36021),
            .in2(_gnd_net_),
            .in3(N__35979),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_14_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__35976),
            .in2(_gnd_net_),
            .in3(N__35940),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_14_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__36456),
            .in2(_gnd_net_),
            .in3(N__36417),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_14_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_14_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_14_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__36414),
            .in2(_gnd_net_),
            .in3(N__36408),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_14_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_14_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_14_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__36405),
            .in2(_gnd_net_),
            .in3(N__36372),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_14_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_14_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_14_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(N__36369),
            .in2(_gnd_net_),
            .in3(N__36330),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_14_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_14_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(N__36327),
            .in2(_gnd_net_),
            .in3(N__36300),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__50770),
            .ce(),
            .sr(N__50344));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_14_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_14_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__36297),
            .in2(_gnd_net_),
            .in3(N__36291),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_14_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_14_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__36288),
            .in2(_gnd_net_),
            .in3(N__36249),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_14_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__36246),
            .in2(_gnd_net_),
            .in3(N__36207),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_14_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__36774),
            .in2(_gnd_net_),
            .in3(N__36735),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_14_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_14_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__36732),
            .in2(_gnd_net_),
            .in3(N__36693),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_14_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__36690),
            .in2(_gnd_net_),
            .in3(N__36657),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_14_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__36654),
            .in2(_gnd_net_),
            .in3(N__36621),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_14_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__36618),
            .in2(_gnd_net_),
            .in3(N__36588),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__50768),
            .ce(),
            .sr(N__50350));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_14_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_14_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__36585),
            .in2(_gnd_net_),
            .in3(N__36540),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_14_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_14_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__36537),
            .in2(_gnd_net_),
            .in3(N__36504),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_14_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_14_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__36501),
            .in2(_gnd_net_),
            .in3(N__36459),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_14_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_14_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__37065),
            .in2(_gnd_net_),
            .in3(N__37032),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_14_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_14_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__37029),
            .in2(_gnd_net_),
            .in3(N__36993),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_14_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_14_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_14_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__36990),
            .in2(_gnd_net_),
            .in3(N__36951),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_14_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_14_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_14_20_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__36948),
            .in2(_gnd_net_),
            .in3(N__36915),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_14_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_14_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_14_20_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__36912),
            .in2(_gnd_net_),
            .in3(N__36879),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__50766),
            .ce(),
            .sr(N__50356));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_14_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_14_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_14_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__36876),
            .in2(_gnd_net_),
            .in3(N__36831),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_14_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_14_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_14_21_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__36828),
            .in2(_gnd_net_),
            .in3(N__36783),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_14_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_14_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_14_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__36780),
            .in2(_gnd_net_),
            .in3(N__37284),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_14_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_14_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_14_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__37281),
            .in2(_gnd_net_),
            .in3(N__37239),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_14_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_14_21_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__37236),
            .in2(_gnd_net_),
            .in3(N__37197),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_14_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_14_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_14_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__37194),
            .in2(_gnd_net_),
            .in3(N__37158),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_14_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_14_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_14_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__37155),
            .in2(_gnd_net_),
            .in3(N__37119),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_14_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_14_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_14_21_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__37116),
            .in2(_gnd_net_),
            .in3(N__37104),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50762),
            .ce(),
            .sr(N__50361));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_14_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_14_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_14_22_5 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_14_22_5  (
            .in0(N__46750),
            .in1(N__46597),
            .in2(N__42600),
            .in3(N__46379),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50759),
            .ce(),
            .sr(N__50366));
    defparam \phase_controller_inst1.S2_LC_14_25_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_14_25_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_14_25_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37479),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50756),
            .ce(N__43659),
            .sr(N__50379));
    defparam \phase_controller_inst1.state_3_LC_15_2_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_15_2_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_15_2_4 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \phase_controller_inst1.state_3_LC_15_2_4  (
            .in0(N__38787),
            .in1(N__37580),
            .in2(N__38855),
            .in3(N__37074),
            .lcout(\phase_controller_inst1.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50907),
            .ce(N__43599),
            .sr(N__50229));
    defparam \phase_controller_inst1.state_1_LC_15_2_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_15_2_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_15_2_6 .LUT_INIT=16'b1110111111100000;
    LogicCell40 \phase_controller_inst1.state_1_LC_15_2_6  (
            .in0(N__37541),
            .in1(N__37579),
            .in2(N__37471),
            .in3(N__37605),
            .lcout(\phase_controller_inst1.N_175_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50907),
            .ce(N__43599),
            .sr(N__50229));
    defparam \phase_controller_inst1.state_2_LC_15_2_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_15_2_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_15_2_7 .LUT_INIT=16'b0011001110100000;
    LogicCell40 \phase_controller_inst1.state_2_LC_15_2_7  (
            .in0(N__38833),
            .in1(N__37542),
            .in2(N__40644),
            .in3(N__37462),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50907),
            .ce(N__43599),
            .sr(N__50229));
    defparam \phase_controller_inst1.stoper_hc.m7_LC_15_3_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m7_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m7_LC_15_3_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.m7_LC_15_3_2  (
            .in0(_gnd_net_),
            .in1(N__37599),
            .in2(_gnd_net_),
            .in3(N__38770),
            .lcout(\phase_controller_inst1.stoper_hc.N_8_0 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNINITI1_LC_15_3_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNINITI1_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_RNINITI1_LC_15_3_3 .LUT_INIT=16'b1100110100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_er_RNINITI1_LC_15_3_3  (
            .in0(N__37574),
            .in1(N__38844),
            .in2(N__37551),
            .in3(N__37548),
            .lcout(\phase_controller_inst1.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.m13_LC_15_3_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.m13_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.m13_LC_15_3_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.m13_LC_15_3_5  (
            .in0(N__38772),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37540),
            .lcout(\phase_controller_inst1.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_RNI9RLH_LC_15_3_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_RNI9RLH_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.S1_RNI9RLH_LC_15_3_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \phase_controller_inst1.S1_RNI9RLH_LC_15_3_7  (
            .in0(N__38771),
            .in1(N__43626),
            .in2(_gnd_net_),
            .in3(N__37328),
            .lcout(S1_RNI9RLH),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_4_LC_15_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_15_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_4_LC_15_4_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \phase_controller_inst1.state_4_LC_15_4_0  (
            .in0(N__37497),
            .in1(N__38702),
            .in2(N__37491),
            .in3(N__37470),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50897),
            .ce(N__43607),
            .sr(N__50237));
    defparam \phase_controller_inst2.state_4_LC_15_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_4_LC_15_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_4_LC_15_4_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \phase_controller_inst2.state_4_LC_15_4_2  (
            .in0(N__38714),
            .in1(N__37422),
            .in2(N__37415),
            .in3(N__37353),
            .lcout(\phase_controller_inst2.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50897),
            .ce(N__43607),
            .sr(N__50237));
    defparam \phase_controller_inst1.S1_LC_15_4_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_15_4_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_15_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38775),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50897),
            .ce(N__43607),
            .sr(N__50237));
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_15_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_15_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__40575),
            .in2(N__37640),
            .in3(N__40586),
            .lcout(\phase_controller_inst1.stoper_hc.N_45_i ),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_15_5_1  (
            .in0(N__48712),
            .in1(N__39024),
            .in2(_gnd_net_),
            .in3(N__37644),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_15_5_2  (
            .in0(N__48809),
            .in1(N__39003),
            .in2(N__37641),
            .in3(N__37626),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_15_5_3  (
            .in0(N__48713),
            .in1(N__38985),
            .in2(_gnd_net_),
            .in3(N__37623),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_15_5_4  (
            .in0(N__48810),
            .in1(N__38964),
            .in2(_gnd_net_),
            .in3(N__37620),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_15_5_5  (
            .in0(N__48714),
            .in1(N__38931),
            .in2(_gnd_net_),
            .in3(N__37617),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_15_5_6  (
            .in0(N__48811),
            .in1(N__38898),
            .in2(_gnd_net_),
            .in3(N__37614),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_15_5_7  (
            .in0(N__48715),
            .in1(N__38877),
            .in2(_gnd_net_),
            .in3(N__37611),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__50890),
            .ce(),
            .sr(N__50240));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_15_6_0  (
            .in0(N__48723),
            .in1(N__39189),
            .in2(_gnd_net_),
            .in3(N__37608),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_15_6_1  (
            .in0(N__48716),
            .in1(N__39171),
            .in2(_gnd_net_),
            .in3(N__37671),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_15_6_2  (
            .in0(N__48720),
            .in1(N__39150),
            .in2(_gnd_net_),
            .in3(N__37668),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_15_6_3  (
            .in0(N__48717),
            .in1(N__39129),
            .in2(_gnd_net_),
            .in3(N__37665),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_15_6_4  (
            .in0(N__48721),
            .in1(N__39102),
            .in2(_gnd_net_),
            .in3(N__37662),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_15_6_5  (
            .in0(N__48718),
            .in1(N__39078),
            .in2(_gnd_net_),
            .in3(N__37659),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_15_6_6  (
            .in0(N__48722),
            .in1(N__39045),
            .in2(_gnd_net_),
            .in3(N__37656),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_15_6_7  (
            .in0(N__48719),
            .in1(N__40795),
            .in2(_gnd_net_),
            .in3(N__37653),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__50883),
            .ce(),
            .sr(N__50245));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_15_7_0  (
            .in0(N__48838),
            .in1(N__40811),
            .in2(_gnd_net_),
            .in3(N__37650),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_15_7_1  (
            .in0(N__48751),
            .in1(N__39331),
            .in2(_gnd_net_),
            .in3(N__37647),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_15_7_2  (
            .in0(N__48839),
            .in1(N__39352),
            .in2(_gnd_net_),
            .in3(N__37737),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_15_7_3  (
            .in0(N__48752),
            .in1(N__39389),
            .in2(_gnd_net_),
            .in3(N__37734),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_15_7_4  (
            .in0(N__48840),
            .in1(N__39412),
            .in2(_gnd_net_),
            .in3(N__37731),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_15_7_5  (
            .in0(N__48753),
            .in1(N__40859),
            .in2(_gnd_net_),
            .in3(N__37728),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_15_7_6  (
            .in0(N__48841),
            .in1(N__40880),
            .in2(_gnd_net_),
            .in3(N__37725),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_15_7_7  (
            .in0(N__48754),
            .in1(N__37721),
            .in2(_gnd_net_),
            .in3(N__37701),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__50873),
            .ce(),
            .sr(N__50249));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_15_8_0  (
            .in0(N__48842),
            .in1(N__37698),
            .in2(_gnd_net_),
            .in3(N__37680),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_15_8_1  (
            .in0(N__48833),
            .in1(N__40691),
            .in2(_gnd_net_),
            .in3(N__37677),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_15_8_2  (
            .in0(N__48843),
            .in1(N__40670),
            .in2(_gnd_net_),
            .in3(N__37674),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_15_8_3  (
            .in0(N__48834),
            .in1(N__37879),
            .in2(_gnd_net_),
            .in3(N__37803),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_15_8_4  (
            .in0(N__48844),
            .in1(N__37858),
            .in2(_gnd_net_),
            .in3(N__37800),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_15_8_5  (
            .in0(N__48835),
            .in1(N__37791),
            .in2(_gnd_net_),
            .in3(N__37797),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_15_8_6  (
            .in0(N__37775),
            .in1(N__48836),
            .in2(_gnd_net_),
            .in3(N__37794),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50863),
            .ce(),
            .sr(N__50256));
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_15_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_31_LC_15_9_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_31_LC_15_9_2  (
            .in0(N__51386),
            .in1(N__49201),
            .in2(_gnd_net_),
            .in3(N__49164),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50851),
            .ce(N__48837),
            .sr(N__50265));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_15_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_15_9_3 .LUT_INIT=16'b1011000011111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_15_9_3  (
            .in0(N__37745),
            .in1(N__37790),
            .in2(N__37776),
            .in3(N__37754),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_15_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_15_9_4 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_15_9_4  (
            .in0(N__37789),
            .in1(N__37774),
            .in2(N__37758),
            .in3(N__37746),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_15_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_30_LC_15_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_30_LC_15_9_5  (
            .in0(N__42187),
            .in1(N__44985),
            .in2(_gnd_net_),
            .in3(N__51387),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50851),
            .ce(N__48837),
            .sr(N__50265));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_9_6 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_15_9_6  (
            .in0(N__48126),
            .in1(N__49200),
            .in2(N__47781),
            .in3(N__39285),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_15_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_15_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_13_LC_15_9_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_13_LC_15_9_7  (
            .in0(_gnd_net_),
            .in1(N__44481),
            .in2(N__37893),
            .in3(N__44349),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50851),
            .ce(N__48837),
            .sr(N__50265));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_10_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_15_10_0  (
            .in0(N__37880),
            .in1(N__37890),
            .in2(N__37842),
            .in3(N__37862),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_15_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_15_10_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_15_10_1  (
            .in0(N__37889),
            .in1(N__37881),
            .in2(N__37863),
            .in3(N__37841),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_15_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_15_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_6_LC_15_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_6_LC_15_10_6  (
            .in0(N__47853),
            .in1(N__39477),
            .in2(_gnd_net_),
            .in3(N__51298),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50841),
            .ce(N__48866),
            .sr(N__50271));
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_15_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_15_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_7_LC_15_11_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_7_LC_15_11_1  (
            .in0(N__51389),
            .in1(N__39517),
            .in2(_gnd_net_),
            .in3(N__48215),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50829),
            .ce(N__48851),
            .sr(N__50279));
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_15_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_15_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_15_LC_15_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_15_LC_15_11_2  (
            .in0(N__45347),
            .in1(N__45364),
            .in2(_gnd_net_),
            .in3(N__51390),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50829),
            .ce(N__48851),
            .sr(N__50279));
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_15_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_25_LC_15_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_25_LC_15_11_3  (
            .in0(N__51388),
            .in1(N__39577),
            .in2(_gnd_net_),
            .in3(N__44618),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50829),
            .ce(N__48851),
            .sr(N__50279));
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_15_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_15_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_20_LC_15_11_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_20_LC_15_11_6  (
            .in0(N__44806),
            .in1(N__39559),
            .in2(_gnd_net_),
            .in3(N__51391),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50829),
            .ce(N__48851),
            .sr(N__50279));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_12_1  (
            .in0(N__39561),
            .in1(N__44805),
            .in2(_gnd_net_),
            .in3(N__51318),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38252),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_15_13_2  (
            .in0(N__51415),
            .in1(N__47855),
            .in2(_gnd_net_),
            .in3(N__39476),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_15_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_15_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__38253),
            .in2(_gnd_net_),
            .in3(N__38296),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_341_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38376),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNI419P_LC_15_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNI419P_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNI419P_LC_15_14_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNI419P_LC_15_14_1  (
            .in0(N__38178),
            .in1(N__49130),
            .in2(_gnd_net_),
            .in3(N__38679),
            .lcout(\current_shift_inst.timer_s1.N_340_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38084),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.start_timer_s1_LC_15_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_15_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_15_15_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_15_15_4  (
            .in0(_gnd_net_),
            .in1(N__38185),
            .in2(_gnd_net_),
            .in3(N__38153),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50792),
            .ce(),
            .sr(N__50312));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_15_5  (
            .in0(N__38519),
            .in1(N__38048),
            .in2(_gnd_net_),
            .in3(N__38029),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_15_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_15_15_7  (
            .in0(N__38520),
            .in1(N__37961),
            .in2(_gnd_net_),
            .in3(N__37933),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_16_2  (
            .in0(N__38518),
            .in1(N__38602),
            .in2(_gnd_net_),
            .in3(N__38569),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_16_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_16_3 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_15_16_3  (
            .in0(N__38279),
            .in1(N__38250),
            .in2(_gnd_net_),
            .in3(N__38303),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_342_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_16_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_15_16_5  (
            .in0(N__38521),
            .in1(N__38377),
            .in2(_gnd_net_),
            .in3(N__38351),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_17_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_17_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_15_17_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_15_17_3  (
            .in0(N__38251),
            .in1(N__38304),
            .in2(_gnd_net_),
            .in3(N__38280),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50777),
            .ce(),
            .sr(N__50328));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_15_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_15_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_15_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38222),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50777),
            .ce(),
            .sr(N__50328));
    defparam \current_shift_inst.timer_s1.running_LC_15_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_15_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_15_17_7 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_15_17_7  (
            .in0(N__38186),
            .in1(N__49119),
            .in2(_gnd_net_),
            .in3(N__38678),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50777),
            .ce(),
            .sr(N__50328));
    defparam \current_shift_inst.stop_timer_s1_er_LC_15_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_er_LC_15_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_er_LC_15_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.stop_timer_s1_er_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38187),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50772),
            .ce(N__38160),
            .sr(N__50336));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_15_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_15_19_2 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_15_19_2  (
            .in0(N__41627),
            .in1(N__41692),
            .in2(N__41794),
            .in3(N__42654),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_15_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_15_19_3 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_15_19_3  (
            .in0(N__40248),
            .in1(N__42374),
            .in2(N__38136),
            .in3(N__46891),
            .lcout(\current_shift_inst.PI_CTRL.N_286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNI8ENL_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNI8ENL_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNI8ENL_LC_15_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNI8ENL_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__49120),
            .in2(_gnd_net_),
            .in3(N__38674),
            .lcout(\current_shift_inst.timer_s1.N_339_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_15_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_15_20_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_15_20_0  (
            .in0(N__46556),
            .in1(N__43403),
            .in2(N__43232),
            .in3(N__43462),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_15_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_15_20_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_15_20_5  (
            .in0(N__42893),
            .in1(N__46234),
            .in2(N__42301),
            .in3(N__42835),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_15_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_15_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_15_20_6  (
            .in0(N__46825),
            .in1(N__43801),
            .in2(N__38640),
            .in3(N__38622),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_15_20_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_15_20_7  (
            .in0(N__38637),
            .in1(N__38628),
            .in2(N__38631),
            .in3(N__40422),
            .lcout(\current_shift_inst.PI_CTRL.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_15_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_15_21_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_15_21_1  (
            .in0(N__43979),
            .in1(N__43166),
            .in2(N__43922),
            .in3(N__43096),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_15_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_15_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_15_21_6  (
            .in0(_gnd_net_),
            .in1(N__42958),
            .in2(_gnd_net_),
            .in3(N__42226),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_15_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_15_22_2 .LUT_INIT=16'b0011110000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_15_22_2  (
            .in0(N__46748),
            .in1(N__41777),
            .in2(N__41742),
            .in3(N__46374),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50763),
            .ce(),
            .sr(N__50362));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_15_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_15_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_15_22_3 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_15_22_3  (
            .in0(N__46372),
            .in1(N__46545),
            .in2(N__42684),
            .in3(N__46749),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50763),
            .ce(),
            .sr(N__50362));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_15_22_6 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_15_22_6  (
            .in0(N__46544),
            .in1(N__46373),
            .in2(N__46781),
            .in3(N__43425),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50763),
            .ce(),
            .sr(N__50362));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_15_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_15_23_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_15_23_1  (
            .in0(N__41646),
            .in1(N__46418),
            .in2(_gnd_net_),
            .in3(N__46751),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50760),
            .ce(),
            .sr(N__50367));
    defparam \phase_controller_inst1.start_timer_hc_LC_16_3_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_16_3_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_16_3_4 .LUT_INIT=16'b0111011101110000;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_16_3_4  (
            .in0(N__38834),
            .in1(N__40615),
            .in2(N__40554),
            .in3(N__38786),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50908),
            .ce(N__43625),
            .sr(N__50230));
    defparam \phase_controller_inst1.test22_LC_16_4_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.test22_LC_16_4_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.test22_LC_16_4_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \phase_controller_inst1.test22_LC_16_4_0  (
            .in0(N__43606),
            .in1(N__38726),
            .in2(_gnd_net_),
            .in3(N__38774),
            .lcout(test22_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50902),
            .ce(),
            .sr(N__50233));
    defparam \phase_controller_inst2.state_0_LC_16_4_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_16_4_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_16_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.state_0_LC_16_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38715),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50902),
            .ce(),
            .sr(N__50233));
    defparam \phase_controller_inst1.state_0_LC_16_4_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_16_4_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_16_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.state_0_LC_16_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38703),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50902),
            .ce(),
            .sr(N__50233));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_16_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_16_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_16_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_16_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40550),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50902),
            .ce(),
            .sr(N__50233));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_0_30_LC_16_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_0_30_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_0_30_LC_16_5_6 .LUT_INIT=16'b0101110111011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_0_30_LC_16_5_6  (
            .in0(N__40551),
            .in1(N__40511),
            .in2(N__40487),
            .in3(N__40463),
            .lcout(\phase_controller_inst1.stoper_hc.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_5_7 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_16_5_7  (
            .in0(N__40512),
            .in1(N__40552),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_16_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_16_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_16_6_0  (
            .in0(_gnd_net_),
            .in1(N__44016),
            .in2(N__38691),
            .in3(N__40570),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_16_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_16_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_16_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_16_6_1  (
            .in0(_gnd_net_),
            .in1(N__47931),
            .in2(N__39012),
            .in3(N__39023),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_16_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_16_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_16_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_16_6_2  (
            .in0(_gnd_net_),
            .in1(N__38991),
            .in2(N__44157),
            .in3(N__39002),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_16_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_16_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_16_6_3  (
            .in0(_gnd_net_),
            .in1(N__40752),
            .in2(N__38973),
            .in3(N__38984),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_16_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_16_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_16_6_4  (
            .in0(_gnd_net_),
            .in1(N__40710),
            .in2(N__38952),
            .in3(N__38963),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_16_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_16_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(N__38943),
            .in2(N__38919),
            .in3(N__38930),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_16_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_16_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_16_6_6  (
            .in0(_gnd_net_),
            .in1(N__38910),
            .in2(N__38886),
            .in3(N__38897),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_16_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_16_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_16_6_7  (
            .in0(_gnd_net_),
            .in1(N__44028),
            .in2(N__38865),
            .in3(N__38876),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_16_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_16_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_16_7_0  (
            .in0(N__39188),
            .in1(N__39177),
            .in2(N__47919),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_16_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_16_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_16_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_16_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(N__40716),
            .in2(N__39159),
            .in3(N__39170),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_16_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_16_7_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(N__47907),
            .in2(N__39138),
            .in3(N__39149),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_16_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_16_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(N__39117),
            .in2(N__40725),
            .in3(N__39128),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_16_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_16_7_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(N__39111),
            .in2(N__39090),
            .in3(N__39101),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_16_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_16_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(N__39306),
            .in2(N__39066),
            .in3(N__39077),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_16_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_16_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_16_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(N__39057),
            .in2(N__39033),
            .in3(N__39044),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_16_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_16_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_16_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(N__40824),
            .in2(N__40770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_16_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_16_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__39315),
            .in2(N__39198),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_16_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_16_8_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__39375),
            .in2(N__39279),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_16_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_16_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__40845),
            .in2(N__40908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_16_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_16_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__39267),
            .in2(N__39258),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_16_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_16_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__40650),
            .in2(N__40704),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_16_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_16_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__39243),
            .in2(N__39231),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_16_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_16_8_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__39216),
            .in2(N__39210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un4_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39201),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_9_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_16_9_0  (
            .in0(N__39354),
            .in1(N__47969),
            .in2(N__39336),
            .in3(N__39297),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_16_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_16_9_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_16_9_1  (
            .in0(N__39296),
            .in1(N__39353),
            .in2(N__47973),
            .in3(N__39335),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_16_9_3  (
            .in0(N__45425),
            .in1(N__45383),
            .in2(_gnd_net_),
            .in3(N__51280),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(elapsed_time_ns_1_RNI13CN9_0_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_14_LC_16_9_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_14_LC_16_9_4  (
            .in0(N__51281),
            .in1(_gnd_net_),
            .in2(N__39309),
            .in3(N__45426),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50864),
            .ce(N__48825),
            .sr(N__50257));
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_16_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_16_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_18_LC_16_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_18_LC_16_9_7  (
            .in0(N__45275),
            .in1(N__45252),
            .in2(_gnd_net_),
            .in3(N__51282),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50864),
            .ce(N__48825),
            .sr(N__50257));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_16_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_16_10_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_16_10_0  (
            .in0(N__45045),
            .in1(N__45183),
            .in2(N__44619),
            .in3(N__44982),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_16_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_16_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_16_10_1  (
            .in0(N__39360),
            .in1(N__39366),
            .in2(N__39288),
            .in3(N__44004),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_10_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_16_10_2  (
            .in0(N__42191),
            .in1(N__51317),
            .in2(_gnd_net_),
            .in3(N__44983),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_10_3 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_10_3  (
            .in0(N__39423),
            .in1(N__39414),
            .in2(N__48894),
            .in3(N__39396),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_16_10_4  (
            .in0(N__51287),
            .in1(N__48961),
            .in2(_gnd_net_),
            .in3(N__48936),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_16_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_16_10_5 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_16_10_5  (
            .in0(N__39422),
            .in1(N__39413),
            .in2(N__48893),
            .in3(N__39395),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_10_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_16_10_6  (
            .in0(N__51286),
            .in1(N__45493),
            .in2(_gnd_net_),
            .in3(N__45470),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_10_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_16_10_7  (
            .in0(N__39518),
            .in1(_gnd_net_),
            .in2(N__48214),
            .in3(N__51288),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_16_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_16_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_16_11_0  (
            .in0(N__51123),
            .in1(N__51763),
            .in2(N__48939),
            .in3(N__44671),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_16_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_16_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_16_11_2  (
            .in0(N__49473),
            .in1(N__45246),
            .in2(N__44808),
            .in3(N__45540),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_16_11_3  (
            .in0(N__45368),
            .in1(N__45346),
            .in2(_gnd_net_),
            .in3(N__51315),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_16_11_4  (
            .in0(N__51314),
            .in1(N__45274),
            .in2(_gnd_net_),
            .in3(N__45247),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_11_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_16_11_6  (
            .in0(N__51313),
            .in1(N__41476),
            .in2(N__45192),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_16_11_7  (
            .in0(N__39579),
            .in1(N__44617),
            .in2(_gnd_net_),
            .in3(N__51316),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_16_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_16_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_25_LC_16_12_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_25_LC_16_12_1  (
            .in0(N__39578),
            .in1(N__51321),
            .in2(_gnd_net_),
            .in3(N__44613),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50830),
            .ce(N__49244),
            .sr(N__50280));
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_16_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_16_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_20_LC_16_12_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_20_LC_16_12_3  (
            .in0(N__39560),
            .in1(N__51319),
            .in2(_gnd_net_),
            .in3(N__44807),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50830),
            .ce(N__49244),
            .sr(N__50280));
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_16_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_24_LC_16_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_24_LC_16_12_5  (
            .in0(N__39543),
            .in1(N__51320),
            .in2(_gnd_net_),
            .in3(N__44670),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50830),
            .ce(N__49244),
            .sr(N__50280));
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_16_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_16_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_7_LC_16_12_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_7_LC_16_12_7  (
            .in0(N__39519),
            .in1(N__51322),
            .in2(_gnd_net_),
            .in3(N__48216),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50830),
            .ce(N__49244),
            .sr(N__50280));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_13_0 .LUT_INIT=16'b0111000101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_16_13_0  (
            .in0(N__41373),
            .in1(N__41396),
            .in2(N__39489),
            .in3(N__39498),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_13_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_16_13_1  (
            .in0(N__39497),
            .in1(N__41372),
            .in2(N__41400),
            .in3(N__39485),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_16_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_16_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_21_LC_16_13_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_21_LC_16_13_3  (
            .in0(N__48962),
            .in1(N__48937),
            .in2(_gnd_net_),
            .in3(N__51518),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50818),
            .ce(N__49242),
            .sr(N__50289));
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_16_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_16_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_5_LC_16_13_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_5_LC_16_13_4  (
            .in0(N__51517),
            .in1(N__47820),
            .in2(_gnd_net_),
            .in3(N__40932),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50818),
            .ce(N__49242),
            .sr(N__50289));
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_16_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_16_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_6_LC_16_13_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_6_LC_16_13_5  (
            .in0(N__47856),
            .in1(N__39472),
            .in2(_gnd_net_),
            .in3(N__51519),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50818),
            .ce(N__49242),
            .sr(N__50289));
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_16_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_16_14_0  (
            .in0(N__49074),
            .in1(N__39445),
            .in2(_gnd_net_),
            .in3(N__39426),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_16_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_16_14_1  (
            .in0(N__49029),
            .in1(N__39772),
            .in2(_gnd_net_),
            .in3(N__39753),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_16_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_16_14_2  (
            .in0(N__49075),
            .in1(N__39748),
            .in2(_gnd_net_),
            .in3(N__39732),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_16_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_16_14_3  (
            .in0(N__49030),
            .in1(N__39727),
            .in2(_gnd_net_),
            .in3(N__39711),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_16_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_16_14_4  (
            .in0(N__49076),
            .in1(N__39700),
            .in2(_gnd_net_),
            .in3(N__39684),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_16_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_16_14_5  (
            .in0(N__49031),
            .in1(N__39673),
            .in2(_gnd_net_),
            .in3(N__39657),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_14_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_16_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_16_14_6  (
            .in0(N__49077),
            .in1(N__39652),
            .in2(_gnd_net_),
            .in3(N__39636),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_14_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_16_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_16_14_7  (
            .in0(N__49032),
            .in1(N__39631),
            .in2(_gnd_net_),
            .in3(N__39615),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__50809),
            .ce(N__40314),
            .sr(N__50297));
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_16_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_16_15_0  (
            .in0(N__49081),
            .in1(N__39604),
            .in2(_gnd_net_),
            .in3(N__39582),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_16_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_16_15_1  (
            .in0(N__49085),
            .in1(N__40015),
            .in2(_gnd_net_),
            .in3(N__39993),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_16_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_16_15_2  (
            .in0(N__49078),
            .in1(N__39988),
            .in2(_gnd_net_),
            .in3(N__39972),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_16_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_16_15_3  (
            .in0(N__49082),
            .in1(N__39967),
            .in2(_gnd_net_),
            .in3(N__39951),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_16_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_16_15_4  (
            .in0(N__49079),
            .in1(N__39943),
            .in2(_gnd_net_),
            .in3(N__39924),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_16_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_16_15_5  (
            .in0(N__49083),
            .in1(N__39913),
            .in2(_gnd_net_),
            .in3(N__39897),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_16_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_16_15_6  (
            .in0(N__49080),
            .in1(N__39886),
            .in2(_gnd_net_),
            .in3(N__39870),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_16_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_16_15_7  (
            .in0(N__49084),
            .in1(N__39865),
            .in2(_gnd_net_),
            .in3(N__39849),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__50801),
            .ce(N__40322),
            .sr(N__50304));
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_16_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_16_16_0  (
            .in0(N__49025),
            .in1(N__39841),
            .in2(_gnd_net_),
            .in3(N__39819),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_16_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_16_16_1  (
            .in0(N__49090),
            .in1(N__39802),
            .in2(_gnd_net_),
            .in3(N__40242),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_16_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_16_16_2  (
            .in0(N__49026),
            .in1(N__40237),
            .in2(_gnd_net_),
            .in3(N__40221),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_16_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_16_16_3  (
            .in0(N__49091),
            .in1(N__40216),
            .in2(_gnd_net_),
            .in3(N__40197),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_16_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_16_16_4  (
            .in0(N__49027),
            .in1(N__40189),
            .in2(_gnd_net_),
            .in3(N__40170),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_16_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_16_16_5  (
            .in0(N__49092),
            .in1(N__40162),
            .in2(_gnd_net_),
            .in3(N__40143),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_16_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_16_16_6  (
            .in0(N__49028),
            .in1(N__40132),
            .in2(_gnd_net_),
            .in3(N__40116),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_16_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_16_16_7  (
            .in0(N__49093),
            .in1(N__40105),
            .in2(_gnd_net_),
            .in3(N__40089),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__50793),
            .ce(N__40315),
            .sr(N__50313));
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_16_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_16_17_0  (
            .in0(N__49086),
            .in1(N__40081),
            .in2(_gnd_net_),
            .in3(N__40059),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_16_17_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__50783),
            .ce(N__40323),
            .sr(N__50320));
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_16_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_16_17_1  (
            .in0(N__49094),
            .in1(N__40045),
            .in2(_gnd_net_),
            .in3(N__40029),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__50783),
            .ce(N__40323),
            .sr(N__50320));
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_16_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_16_17_2  (
            .in0(N__49087),
            .in1(N__40405),
            .in2(_gnd_net_),
            .in3(N__40386),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__50783),
            .ce(N__40323),
            .sr(N__50320));
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_16_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_16_17_3  (
            .in0(N__49095),
            .in1(N__40381),
            .in2(_gnd_net_),
            .in3(N__40365),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__50783),
            .ce(N__40323),
            .sr(N__50320));
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_16_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_16_17_4  (
            .in0(N__49088),
            .in1(N__40361),
            .in2(_gnd_net_),
            .in3(N__40347),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__50783),
            .ce(N__40323),
            .sr(N__50320));
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_16_17_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_16_17_5  (
            .in0(N__40337),
            .in1(N__49089),
            .in2(_gnd_net_),
            .in3(N__40344),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50783),
            .ce(N__40323),
            .sr(N__50320));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_16_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_16_18_0 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_16_18_0  (
            .in0(N__41324),
            .in1(N__40280),
            .in2(N__40266),
            .in3(N__41346),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_16_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_16_18_1 .LUT_INIT=16'b1111011100110001;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_16_18_1  (
            .in0(N__41345),
            .in1(N__41323),
            .in2(N__40284),
            .in3(N__40265),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_16_18_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_16_18_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_16_18_5  (
            .in0(N__47894),
            .in1(N__40736),
            .in2(_gnd_net_),
            .in3(N__51501),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(elapsed_time_ns_1_RNIV0CN9_0_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_12_LC_16_18_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_12_LC_16_18_6  (
            .in0(N__51502),
            .in1(_gnd_net_),
            .in2(N__40251),
            .in3(N__47895),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50778),
            .ce(N__49239),
            .sr(N__50329));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_16_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_16_19_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_16_19_5  (
            .in0(N__42570),
            .in1(N__42456),
            .in2(_gnd_net_),
            .in3(N__46943),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_16_20_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_16_20_2  (
            .in0(N__42458),
            .in1(N__46936),
            .in2(N__46892),
            .in3(N__42373),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_16_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_16_20_3 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_16_20_3  (
            .in0(N__42659),
            .in1(N__41614),
            .in2(N__40428),
            .in3(N__42561),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_16_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_16_20_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_16_20_4  (
            .in0(N__40416),
            .in1(N__43855),
            .in2(N__40425),
            .in3(N__43286),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_16_20_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_16_20_6  (
            .in0(N__43512),
            .in1(N__42717),
            .in2(N__43348),
            .in3(N__42776),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_16_21_1 .LUT_INIT=16'b1100111011001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_16_21_1  (
            .in0(N__46560),
            .in1(N__43035),
            .in2(N__46764),
            .in3(N__46401),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50769),
            .ce(),
            .sr(N__50351));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_16_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_16_21_2 .LUT_INIT=16'b1011101110101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_16_21_2  (
            .in0(N__42855),
            .in1(N__46713),
            .in2(N__46421),
            .in3(N__46565),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50769),
            .ce(),
            .sr(N__50351));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_16_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_16_21_3 .LUT_INIT=16'b1100111011001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_16_21_3  (
            .in0(N__46561),
            .in1(N__42924),
            .in2(N__46765),
            .in3(N__46402),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50769),
            .ce(),
            .sr(N__50351));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_16_21_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_16_21_4  (
            .in0(N__46394),
            .in1(N__46563),
            .in2(N__43488),
            .in3(N__46711),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50769),
            .ce(),
            .sr(N__50351));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_16_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_16_21_6 .LUT_INIT=16'b1011101110101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_16_21_6  (
            .in0(N__42252),
            .in1(N__46712),
            .in2(N__46420),
            .in3(N__46564),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50769),
            .ce(),
            .sr(N__50351));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_16_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_16_21_7 .LUT_INIT=16'b1100010011000101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_16_21_7  (
            .in0(N__46562),
            .in1(N__42327),
            .in2(N__46766),
            .in3(N__46403),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50769),
            .ce(),
            .sr(N__50351));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_16_22_0 .LUT_INIT=16'b1111001011100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_16_22_0  (
            .in0(N__46539),
            .in1(N__46778),
            .in2(N__43185),
            .in3(N__46417),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50767),
            .ce(),
            .sr(N__50357));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_16_22_1 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_16_22_1  (
            .in0(N__46776),
            .in1(N__46542),
            .in2(N__46424),
            .in3(N__43305),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50767),
            .ce(),
            .sr(N__50357));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_16_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_16_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_16_22_2 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_16_22_2  (
            .in0(N__46538),
            .in1(N__46416),
            .in2(N__42798),
            .in3(N__46779),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50767),
            .ce(),
            .sr(N__50357));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_22_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_16_22_3 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_16_22_3  (
            .in0(N__46777),
            .in1(N__46543),
            .in2(N__46425),
            .in3(N__43251),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50767),
            .ce(),
            .sr(N__50357));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_16_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_16_22_5 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_16_22_5  (
            .in0(N__46775),
            .in1(N__46541),
            .in2(N__46423),
            .in3(N__43371),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50767),
            .ce(),
            .sr(N__50357));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_16_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_16_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_16_22_7 .LUT_INIT=16'b1111111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_16_22_7  (
            .in0(N__46774),
            .in1(N__46540),
            .in2(N__46422),
            .in3(N__42741),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50767),
            .ce(),
            .sr(N__50357));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_16_23_0 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_16_23_0  (
            .in0(N__46388),
            .in1(N__46583),
            .in2(N__43824),
            .in3(N__46762),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50764),
            .ce(),
            .sr(N__50363));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_16_23_1 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_16_23_1  (
            .in0(N__46579),
            .in1(N__46390),
            .in2(N__46782),
            .in3(N__43062),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50764),
            .ce(),
            .sr(N__50363));
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_16_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_16_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_31_LC_16_23_3 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_31_LC_16_23_3  (
            .in0(N__46581),
            .in1(N__46392),
            .in2(N__46784),
            .in3(N__43743),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50764),
            .ce(),
            .sr(N__50363));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_16_23_4 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_16_23_4  (
            .in0(N__46389),
            .in1(N__46584),
            .in2(N__43758),
            .in3(N__46763),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50764),
            .ce(),
            .sr(N__50363));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_16_23_5 .LUT_INIT=16'b1111111000001010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_16_23_5  (
            .in0(N__46580),
            .in1(N__46391),
            .in2(N__46783),
            .in3(N__43881),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50764),
            .ce(),
            .sr(N__50363));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_16_23_6 .LUT_INIT=16'b1111000011101100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_16_23_6  (
            .in0(N__46387),
            .in1(N__46582),
            .in2(N__43131),
            .in3(N__46761),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50764),
            .ce(),
            .sr(N__50363));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_16_24_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_16_24_1 .LUT_INIT=16'b1111111000001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_16_24_1  (
            .in0(N__46393),
            .in1(N__46546),
            .in2(N__46785),
            .in3(N__43941),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50761),
            .ce(),
            .sr(N__50368));
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_LC_17_4_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_LC_17_4_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_er_LC_17_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_er_LC_17_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40517),
            .lcout(\phase_controller_inst1.stoper_hc.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50909),
            .ce(N__40437),
            .sr(N__50231));
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_17_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_17_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_17_5_0 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_17_5_0  (
            .in0(N__48711),
            .in1(N__40587),
            .in2(_gnd_net_),
            .in3(N__40574),
            .lcout(\phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50903),
            .ce(),
            .sr(N__50234));
    defparam \phase_controller_inst1.stoper_hc.running_LC_17_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_17_5_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_17_5_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_17_5_1  (
            .in0(N__40516),
            .in1(N__40486),
            .in2(_gnd_net_),
            .in3(N__40446),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50903),
            .ce(),
            .sr(N__50234));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_30_LC_17_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_30_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_30_LC_17_6_3 .LUT_INIT=16'b1101110101011101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNIR1181_30_LC_17_6_3  (
            .in0(N__40553),
            .in1(N__40518),
            .in2(N__40488),
            .in3(N__40464),
            .lcout(\phase_controller_inst1.stoper_hc.N_46 ),
            .ltout(\phase_controller_inst1.stoper_hc.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_sbtinv_LC_17_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_sbtinv_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_sbtinv_LC_17_6_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_sbtinv_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40440),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.N_46_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_6_6 .LUT_INIT=16'b0000100011001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_17_6_6  (
            .in0(N__40760),
            .in1(N__44169),
            .in2(N__40796),
            .in3(N__40818),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_6_7 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_17_6_7  (
            .in0(N__40817),
            .in1(N__40761),
            .in2(N__40797),
            .in3(N__44168),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_17_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_17_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_16_LC_17_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_16_LC_17_7_0  (
            .in0(N__45471),
            .in1(N__51440),
            .in2(_gnd_net_),
            .in3(N__45501),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50891),
            .ce(N__48852),
            .sr(N__50241));
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_4_LC_17_7_2  (
            .in0(N__47999),
            .in1(N__51441),
            .in2(_gnd_net_),
            .in3(N__48037),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50891),
            .ce(N__48852),
            .sr(N__50241));
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_17_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_17_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_12_LC_17_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_12_LC_17_7_3  (
            .in0(N__51437),
            .in1(N__47888),
            .in2(_gnd_net_),
            .in3(N__40746),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50891),
            .ce(N__48852),
            .sr(N__50241));
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_10_LC_17_7_4  (
            .in0(N__48308),
            .in1(N__51439),
            .in2(_gnd_net_),
            .in3(N__48284),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50891),
            .ce(N__48852),
            .sr(N__50241));
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_17_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_17_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_5_LC_17_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_5_LC_17_7_5  (
            .in0(N__51438),
            .in1(N__47818),
            .in2(_gnd_net_),
            .in3(N__40924),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50891),
            .ce(N__48852),
            .sr(N__50241));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_8_0 .LUT_INIT=16'b0000100010101110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_8_0  (
            .in0(N__44037),
            .in1(N__40941),
            .in2(N__40692),
            .in3(N__40669),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_17_8_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_17_8_1  (
            .in0(N__40940),
            .in1(N__40690),
            .in2(N__40671),
            .in3(N__44036),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_17_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_17_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_26_LC_17_8_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_26_LC_17_8_2  (
            .in0(N__51436),
            .in1(N__41483),
            .in2(_gnd_net_),
            .in3(N__45190),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50884),
            .ce(N__48812),
            .sr(N__50246));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_8_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_8_5  (
            .in0(N__40928),
            .in1(N__47817),
            .in2(_gnd_net_),
            .in3(N__51435),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_9_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_9_0  (
            .in0(N__40896),
            .in1(N__40887),
            .in2(N__47955),
            .in3(N__40866),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_17_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_22_LC_17_9_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_22_LC_17_9_2  (
            .in0(N__51762),
            .in1(N__51723),
            .in2(N__51460),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50874),
            .ce(N__48853),
            .sr(N__50250));
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_17_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_17_9_4 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_17_9_4  (
            .in0(N__40895),
            .in1(N__40886),
            .in2(N__47954),
            .in3(N__40865),
            .lcout(\phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_17_10_0  (
            .in0(N__41160),
            .in1(N__44929),
            .in2(_gnd_net_),
            .in3(N__40836),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_17_10_1  (
            .in0(N__41177),
            .in1(N__48109),
            .in2(_gnd_net_),
            .in3(N__40833),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_17_10_2  (
            .in0(N__41161),
            .in1(N__44324),
            .in2(_gnd_net_),
            .in3(N__40830),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_17_10_3  (
            .in0(N__41178),
            .in1(N__44300),
            .in2(_gnd_net_),
            .in3(N__40827),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_17_10_4  (
            .in0(N__41162),
            .in1(N__44276),
            .in2(_gnd_net_),
            .in3(N__40968),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_17_10_5  (
            .in0(N__41179),
            .in1(N__44252),
            .in2(_gnd_net_),
            .in3(N__40965),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_17_10_6  (
            .in0(N__41163),
            .in1(N__44228),
            .in2(_gnd_net_),
            .in3(N__40962),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_17_10_7  (
            .in0(N__41180),
            .in1(N__44570),
            .in2(_gnd_net_),
            .in3(N__40959),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__50865),
            .ce(N__41049),
            .sr(N__50258));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_17_11_0  (
            .in0(N__41159),
            .in1(N__44546),
            .in2(_gnd_net_),
            .in3(N__40956),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_17_11_1  (
            .in0(N__41167),
            .in1(N__44522),
            .in2(_gnd_net_),
            .in3(N__40953),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_17_11_2  (
            .in0(N__41156),
            .in1(N__44498),
            .in2(_gnd_net_),
            .in3(N__40950),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_17_11_3  (
            .in0(N__41164),
            .in1(N__44441),
            .in2(_gnd_net_),
            .in3(N__40947),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_17_11_4  (
            .in0(N__41157),
            .in1(N__44417),
            .in2(_gnd_net_),
            .in3(N__40944),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_17_11_5  (
            .in0(N__41165),
            .in1(N__44393),
            .in2(_gnd_net_),
            .in3(N__40995),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_17_11_6  (
            .in0(N__41158),
            .in1(N__44369),
            .in2(_gnd_net_),
            .in3(N__40992),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_17_11_7  (
            .in0(N__41166),
            .in1(N__44873),
            .in2(_gnd_net_),
            .in3(N__40989),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__50852),
            .ce(N__41048),
            .sr(N__50266));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_17_12_0  (
            .in0(N__41152),
            .in1(N__44849),
            .in2(_gnd_net_),
            .in3(N__40986),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_17_12_1  (
            .in0(N__41181),
            .in1(N__44825),
            .in2(_gnd_net_),
            .in3(N__40983),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_17_12_2  (
            .in0(N__41153),
            .in1(N__44768),
            .in2(_gnd_net_),
            .in3(N__40980),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_17_12_3  (
            .in0(N__41182),
            .in1(N__44744),
            .in2(_gnd_net_),
            .in3(N__40977),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_17_12_4  (
            .in0(N__41154),
            .in1(N__44720),
            .in2(_gnd_net_),
            .in3(N__40974),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_17_12_5  (
            .in0(N__41183),
            .in1(N__44696),
            .in2(_gnd_net_),
            .in3(N__40971),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_17_12_6  (
            .in0(N__41155),
            .in1(N__44636),
            .in2(_gnd_net_),
            .in3(N__41205),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_17_12_7  (
            .in0(N__41184),
            .in1(N__45209),
            .in2(_gnd_net_),
            .in3(N__41202),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__50842),
            .ce(N__41041),
            .sr(N__50272));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_17_13_0  (
            .in0(N__41137),
            .in1(N__45134),
            .in2(_gnd_net_),
            .in3(N__41199),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__50831),
            .ce(N__41040),
            .sr(N__50281));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_17_13_1  (
            .in0(N__41141),
            .in1(N__45110),
            .in2(_gnd_net_),
            .in3(N__41196),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__50831),
            .ce(N__41040),
            .sr(N__50281));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_17_13_2  (
            .in0(N__41138),
            .in1(N__45074),
            .in2(_gnd_net_),
            .in3(N__41193),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__50831),
            .ce(N__41040),
            .sr(N__50281));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_17_13_3  (
            .in0(N__41142),
            .in1(N__45002),
            .in2(_gnd_net_),
            .in3(N__41190),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__50831),
            .ce(N__41040),
            .sr(N__50281));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_17_13_4  (
            .in0(N__41139),
            .in1(N__45090),
            .in2(_gnd_net_),
            .in3(N__41187),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__50831),
            .ce(N__41040),
            .sr(N__50281));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_17_13_5  (
            .in0(N__45018),
            .in1(N__41140),
            .in2(_gnd_net_),
            .in3(N__41052),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50831),
            .ce(N__41040),
            .sr(N__50281));
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_17_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_17_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_c_inv_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__46980),
            .in2(N__41243),
            .in3(N__46995),
            .lcout(\phase_controller_inst2.stoper_hc.N_265_i ),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_14_1  (
            .in0(N__47155),
            .in1(N__45749),
            .in2(_gnd_net_),
            .in3(N__41247),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_14_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_14_2  (
            .in0(N__47144),
            .in1(N__45722),
            .in2(N__41244),
            .in3(N__41229),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_14_3  (
            .in0(N__47156),
            .in1(N__45692),
            .in2(_gnd_net_),
            .in3(N__41226),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_14_4  (
            .in0(N__47145),
            .in1(N__45668),
            .in2(_gnd_net_),
            .in3(N__41223),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_14_5  (
            .in0(N__47157),
            .in1(N__45617),
            .in2(_gnd_net_),
            .in3(N__41220),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_14_6  (
            .in0(N__47146),
            .in1(N__45581),
            .in2(_gnd_net_),
            .in3(N__41217),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_14_7  (
            .in0(N__47158),
            .in1(N__45995),
            .in2(_gnd_net_),
            .in3(N__41214),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7 ),
            .clk(N__50819),
            .ce(),
            .sr(N__50290));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_15_0  (
            .in0(N__47165),
            .in1(N__45968),
            .in2(_gnd_net_),
            .in3(N__41211),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9 ),
            .ltout(),
            .carryin(bfn_17_15_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_15_1  (
            .in0(N__47140),
            .in1(N__45947),
            .in2(_gnd_net_),
            .in3(N__41208),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_15_2  (
            .in0(N__47162),
            .in1(N__45923),
            .in2(_gnd_net_),
            .in3(N__41274),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_15_3  (
            .in0(N__47141),
            .in1(N__45887),
            .in2(_gnd_net_),
            .in3(N__41271),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_15_4  (
            .in0(N__47163),
            .in1(N__45860),
            .in2(_gnd_net_),
            .in3(N__41268),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_15_5  (
            .in0(N__47142),
            .in1(N__45824),
            .in2(_gnd_net_),
            .in3(N__41265),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_15_6  (
            .in0(N__47164),
            .in1(N__45779),
            .in2(_gnd_net_),
            .in3(N__41262),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_15_7  (
            .in0(N__47143),
            .in1(N__44913),
            .in2(_gnd_net_),
            .in3(N__41259),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15 ),
            .clk(N__50810),
            .ce(),
            .sr(N__50298));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_16_0  (
            .in0(N__47147),
            .in1(N__44893),
            .in2(_gnd_net_),
            .in3(N__41256),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17 ),
            .ltout(),
            .carryin(bfn_17_16_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_16_1  (
            .in0(N__47133),
            .in1(N__45294),
            .in2(_gnd_net_),
            .in3(N__41253),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_16_2  (
            .in0(N__47148),
            .in1(N__45311),
            .in2(_gnd_net_),
            .in3(N__41250),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_16_3  (
            .in0(N__47134),
            .in1(N__41390),
            .in2(_gnd_net_),
            .in3(N__41376),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_16_4  (
            .in0(N__47149),
            .in1(N__41371),
            .in2(_gnd_net_),
            .in3(N__41355),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_16_5  (
            .in0(N__47135),
            .in1(N__51013),
            .in2(_gnd_net_),
            .in3(N__41352),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_16_6  (
            .in0(N__47150),
            .in1(N__51043),
            .in2(_gnd_net_),
            .in3(N__41349),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_16_7  (
            .in0(N__47136),
            .in1(N__41344),
            .in2(_gnd_net_),
            .in3(N__41328),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23 ),
            .clk(N__50802),
            .ce(),
            .sr(N__50305));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_17_0  (
            .in0(N__47151),
            .in1(N__41325),
            .in2(_gnd_net_),
            .in3(N__41310),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25 ),
            .ltout(),
            .carryin(bfn_17_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_17_1  (
            .in0(N__47159),
            .in1(N__41499),
            .in2(_gnd_net_),
            .in3(N__41307),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_17_2  (
            .in0(N__47152),
            .in1(N__41516),
            .in2(_gnd_net_),
            .in3(N__41304),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_17_3  (
            .in0(N__47160),
            .in1(N__41291),
            .in2(_gnd_net_),
            .in3(N__41277),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_17_4  (
            .in0(N__47153),
            .in1(N__41540),
            .in2(_gnd_net_),
            .in3(N__41526),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_17_5  (
            .in0(N__47161),
            .in1(N__41415),
            .in2(_gnd_net_),
            .in3(N__41523),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29 ),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_17_6  (
            .in0(N__47154),
            .in1(N__41444),
            .in2(_gnd_net_),
            .in3(N__41520),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50794),
            .ce(),
            .sr(N__50314));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_18_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_17_18_0  (
            .in0(N__41498),
            .in1(N__49337),
            .in2(N__41517),
            .in3(N__41454),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_17_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_17_18_1 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_17_18_1  (
            .in0(N__41453),
            .in1(N__41515),
            .in2(N__49341),
            .in3(N__41497),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_17_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_26_LC_17_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_26_LC_17_18_2  (
            .in0(N__41484),
            .in1(N__45191),
            .in2(_gnd_net_),
            .in3(N__51622),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50784),
            .ce(N__49240),
            .sr(N__50321));
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_17_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_17_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_31_LC_17_18_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_31_LC_17_18_4  (
            .in0(N__49205),
            .in1(N__49154),
            .in2(_gnd_net_),
            .in3(N__51623),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50784),
            .ce(N__49240),
            .sr(N__50321));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_17_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_17_18_5 .LUT_INIT=16'b1101000011111101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_17_18_5  (
            .in0(N__41413),
            .in1(N__42170),
            .in2(N__41445),
            .in3(N__41423),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_18_6 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_17_18_6  (
            .in0(N__42171),
            .in1(N__41440),
            .in2(N__41427),
            .in3(N__41414),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_17_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_17_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_30_LC_17_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_30_LC_17_18_7  (
            .in0(N__51621),
            .in1(N__42198),
            .in2(_gnd_net_),
            .in3(N__44984),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50784),
            .ce(N__49240),
            .sr(N__50321));
    defparam \phase_controller_inst2.start_timer_hc_LC_17_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_17_19_2 .LUT_INIT=16'b0000111000001100;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_17_19_2  (
            .in0(N__41925),
            .in1(N__42005),
            .in2(N__42162),
            .in3(N__42128),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50779),
            .ce(N__43641),
            .sr(N__50330));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0_30_LC_17_19_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0_30_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0_30_LC_17_19_3 .LUT_INIT=16'b0111010111110101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0_30_LC_17_19_3  (
            .in0(N__42003),
            .in1(N__42089),
            .in2(N__42068),
            .in3(N__47174),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_30_LC_17_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_30_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_30_LC_17_19_4 .LUT_INIT=16'b1100010011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971_30_LC_17_19_4  (
            .in0(N__42090),
            .in1(N__42064),
            .in2(N__47178),
            .in3(N__42004),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIVQ971Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_17_19_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_17_19_7 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \phase_controller_inst2.state_3_LC_17_19_7  (
            .in0(N__41819),
            .in1(N__41961),
            .in2(N__41946),
            .in3(N__41924),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50779),
            .ce(N__43641),
            .sr(N__50330));
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_17_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__41790),
            .in2(N__41738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_17_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__41693),
            .in2(N__41664),
            .in3(N__41634),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_17_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__41613),
            .in2(N__41586),
            .in3(N__41556),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__42655),
            .in2(N__42618),
            .in3(N__42585),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__42582),
            .in2(N__42569),
            .in3(N__42507),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__46872),
            .in2(N__42504),
            .in3(N__42486),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__46932),
            .in2(N__42483),
            .in3(N__42465),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__42457),
            .in2(N__42420),
            .in3(N__42387),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__42369),
            .in2(N__42345),
            .in3(N__42321),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__42292),
            .in2(N__42273),
            .in3(N__42246),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__42222),
            .in2(N__43053),
            .in3(N__43029),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(N__46806),
            .in2(N__43026),
            .in3(N__43008),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__46219),
            .in2(N__43005),
            .in3(N__42987),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__42959),
            .in2(N__42942),
            .in3(N__42918),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__42892),
            .in2(N__42873),
            .in3(N__42849),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_17_21_7  (
            .in0(_gnd_net_),
            .in1(N__42825),
            .in2(N__46167),
            .in3(N__42789),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_17_22_0  (
            .in0(_gnd_net_),
            .in1(N__42762),
            .in2(N__47451),
            .in3(N__42735),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_17_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__42718),
            .in2(N__47406),
            .in3(N__42672),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(N__43513),
            .in2(N__47358),
            .in3(N__43476),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(N__43461),
            .in2(N__47328),
            .in3(N__43416),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(N__43395),
            .in2(N__47298),
            .in3(N__43365),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(N__43335),
            .in2(N__47271),
            .in3(N__43299),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_17_22_6  (
            .in0(_gnd_net_),
            .in1(N__43272),
            .in2(N__47241),
            .in3(N__43245),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_17_22_7  (
            .in0(_gnd_net_),
            .in1(N__43218),
            .in2(N__47211),
            .in3(N__43176),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_17_23_0  (
            .in0(_gnd_net_),
            .in1(N__43155),
            .in2(N__47748),
            .in3(N__43119),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_17_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__43092),
            .in2(N__47712),
            .in3(N__43056),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_17_23_2  (
            .in0(_gnd_net_),
            .in1(N__47682),
            .in2(N__43977),
            .in3(N__43935),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__43905),
            .in2(N__47652),
            .in3(N__43875),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_17_23_4  (
            .in0(_gnd_net_),
            .in1(N__43842),
            .in2(N__47625),
            .in3(N__43815),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_17_23_5  (
            .in0(_gnd_net_),
            .in1(N__43785),
            .in2(N__47514),
            .in3(N__43749),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_17_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_17_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_17_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_17_23_6  (
            .in0(N__46516),
            .in1(N__47499),
            .in2(N__43716),
            .in3(N__43746),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_17_24_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_17_24_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_17_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_17_24_2  (
            .in0(_gnd_net_),
            .in1(N__47607),
            .in2(_gnd_net_),
            .in3(N__43737),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_5_LC_17_30_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_5_LC_17_30_3 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_5_LC_17_30_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.state_5_LC_17_30_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(GNDG0),
            .lcout(\phase_controller_inst1.stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50752),
            .ce(N__43669),
            .sr(N__50384));
    defparam \phase_controller_inst1.test_LC_17_30_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.test_LC_17_30_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.test_LC_17_30_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \phase_controller_inst1.test_LC_17_30_5  (
            .in0(_gnd_net_),
            .in1(N__43700),
            .in2(_gnd_net_),
            .in3(N__43707),
            .lcout(test_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50752),
            .ce(N__43669),
            .sr(N__50384));
    defparam \phase_controller_inst2.stoper_tr.time_passed_er_LC_18_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_er_LC_18_5_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_er_LC_18_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_er_LC_18_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44127),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50910),
            .ce(N__44046),
            .sr(N__50232));
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_18_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_18_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_17_LC_18_6_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_17_LC_18_6_3  (
            .in0(N__45543),
            .in1(N__45561),
            .in2(_gnd_net_),
            .in3(N__51446),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50904),
            .ce(N__48867),
            .sr(N__50235));
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_18_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_18_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_3_LC_18_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_3_LC_18_6_6  (
            .in0(N__51445),
            .in1(N__48459),
            .in2(_gnd_net_),
            .in3(N__48429),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50904),
            .ce(N__48867),
            .sr(N__50235));
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_18_7_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_18_7_1  (
            .in0(N__44145),
            .in1(N__44074),
            .in2(_gnd_net_),
            .in3(N__44058),
            .lcout(\phase_controller_inst2.running ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50898),
            .ce(),
            .sr(N__50238));
    defparam \phase_controller_inst2.stoper_tr.time_passed_sbtinv_LC_18_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_sbtinv_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_sbtinv_LC_18_7_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_sbtinv_LC_18_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44057),
            .lcout(\phase_controller_inst2.stoper_tr.N_39_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_18_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_18_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_27_LC_18_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_27_LC_18_8_0  (
            .in0(N__51442),
            .in1(N__51693),
            .in2(_gnd_net_),
            .in3(N__51654),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50892),
            .ce(N__48824),
            .sr(N__50242));
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_18_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_18_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_8_LC_18_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_8_LC_18_8_4  (
            .in0(N__51443),
            .in1(N__48597),
            .in2(_gnd_net_),
            .in3(N__48567),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50892),
            .ce(N__48824),
            .sr(N__50242));
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_18_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_1_LC_18_8_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_1_LC_18_8_7  (
            .in0(N__49380),
            .in1(N__49421),
            .in2(_gnd_net_),
            .in3(N__51444),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50892),
            .ce(N__48824),
            .sr(N__50242));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_18_9_1  (
            .in0(N__45345),
            .in1(N__45415),
            .in2(N__44479),
            .in3(N__45462),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_9_5 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_18_9_5  (
            .in0(N__51431),
            .in1(N__44345),
            .in2(N__44480),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(elapsed_time_ns_1_RNI02CN9_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_18_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_13_LC_18_9_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_13_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(N__44475),
            .in2(N__44334),
            .in3(N__51432),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50885),
            .ce(N__49251),
            .sr(N__50247));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__44323),
            .in2(N__44936),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__44299),
            .in2(N__48116),
            .in3(N__44331),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(N__44275),
            .in2(N__44328),
            .in3(N__44307),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__44251),
            .in2(N__44304),
            .in3(N__44283),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_18_10_4  (
            .in0(_gnd_net_),
            .in1(N__44227),
            .in2(N__44280),
            .in3(N__44259),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__44569),
            .in2(N__44256),
            .in3(N__44235),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__44545),
            .in2(N__44232),
            .in3(N__44211),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(N__44521),
            .in2(N__44574),
            .in3(N__44553),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__50875),
            .ce(N__48089),
            .sr(N__50251));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__44497),
            .in2(N__44550),
            .in3(N__44529),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__44440),
            .in2(N__44526),
            .in3(N__44505),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__44416),
            .in2(N__44502),
            .in3(N__44448),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__44392),
            .in2(N__44445),
            .in3(N__44424),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__44368),
            .in2(N__44421),
            .in3(N__44400),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__44872),
            .in2(N__44397),
            .in3(N__44376),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__44848),
            .in2(N__44373),
            .in3(N__44352),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__44824),
            .in2(N__44877),
            .in3(N__44856),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__50866),
            .ce(N__48088),
            .sr(N__50259));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__44767),
            .in2(N__44853),
            .in3(N__44832),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__44743),
            .in2(N__44829),
            .in3(N__44775),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__44719),
            .in2(N__44772),
            .in3(N__44751),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(N__44695),
            .in2(N__44748),
            .in3(N__44727),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(N__44635),
            .in2(N__44724),
            .in3(N__44703),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(N__45208),
            .in2(N__44700),
            .in3(N__44643),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__45133),
            .in2(N__44640),
            .in3(N__44577),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(N__45109),
            .in2(N__45213),
            .in3(N__45141),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__50853),
            .ce(N__48087),
            .sr(N__50267));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__45073),
            .in2(N__45138),
            .in3(N__45117),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__50843),
            .ce(N__48074),
            .sr(N__50273));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__45001),
            .in2(N__45114),
            .in3(N__45093),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__50843),
            .ce(N__48074),
            .sr(N__50273));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__45089),
            .in2(N__45078),
            .in3(N__45021),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__50843),
            .ce(N__48074),
            .sr(N__50273));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__45017),
            .in2(N__45006),
            .in3(N__44946),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__50843),
            .ce(N__48074),
            .sr(N__50273));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44943),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50843),
            .ce(N__48074),
            .sr(N__50273));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_13_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44940),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50843),
            .ce(N__48074),
            .sr(N__50273));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_14_0 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_14_0  (
            .in0(N__44911),
            .in1(N__44894),
            .in2(N__45513),
            .in3(N__45435),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_14_1 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_14_1  (
            .in0(N__45434),
            .in1(N__44912),
            .in2(N__44898),
            .in3(N__45509),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_14_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_14_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_14_2  (
            .in0(N__45541),
            .in1(N__45557),
            .in2(_gnd_net_),
            .in3(N__51600),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(elapsed_time_ns_1_RNI46CN9_0_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_17_LC_18_14_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_17_LC_18_14_3  (
            .in0(N__51603),
            .in1(_gnd_net_),
            .in2(N__45546),
            .in3(N__45542),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50832),
            .ce(N__49245),
            .sr(N__50282));
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_16_LC_18_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_16_LC_18_14_5  (
            .in0(N__51602),
            .in1(N__45500),
            .in2(_gnd_net_),
            .in3(N__45466),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50832),
            .ce(N__49245),
            .sr(N__50282));
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_18_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_18_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_14_LC_18_14_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_14_LC_18_14_6  (
            .in0(N__45424),
            .in1(N__45393),
            .in2(_gnd_net_),
            .in3(N__51604),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50832),
            .ce(N__49245),
            .sr(N__50282));
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_18_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_18_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_15_LC_18_14_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_15_LC_18_14_7  (
            .in0(N__51601),
            .in1(N__45372),
            .in2(_gnd_net_),
            .in3(N__45348),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50832),
            .ce(N__49245),
            .sr(N__50282));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_15_0 .LUT_INIT=16'b0100000011110100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_18_15_0  (
            .in0(N__45293),
            .in1(N__45222),
            .in2(N__49440),
            .in3(N__45310),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_18_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_18_15_1 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_18_15_1  (
            .in0(N__45221),
            .in1(N__49439),
            .in2(N__45312),
            .in3(N__45292),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_18_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_18_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_18_LC_18_15_2 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_18_LC_18_15_2  (
            .in0(N__45279),
            .in1(N__45251),
            .in2(N__51624),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50820),
            .ce(N__49243),
            .sr(N__50291));
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_18_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_18_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_4_LC_18_15_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_4_LC_18_15_7  (
            .in0(N__48036),
            .in1(N__51612),
            .in2(_gnd_net_),
            .in3(N__48003),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50820),
            .ce(N__49243),
            .sr(N__50291));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_18_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_18_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(N__49350),
            .in2(N__45765),
            .in3(N__46976),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_1 ),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_18_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_18_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(N__48471),
            .in2(N__45735),
            .in3(N__45753),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_18_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_18_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(N__45708),
            .in2(N__48399),
            .in3(N__45726),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_18_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_18_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_18_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_18_16_3  (
            .in0(_gnd_net_),
            .in1(N__45702),
            .in2(N__45678),
            .in3(N__45696),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_18_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_18_16_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_18_16_4  (
            .in0(N__45669),
            .in1(N__45654),
            .in2(N__45642),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_18_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_18_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__45603),
            .in2(N__45633),
            .in3(N__45618),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_18_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_18_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(N__45567),
            .in2(N__45597),
            .in3(N__45582),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_18_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_18_16_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_18_16_7  (
            .in0(N__45996),
            .in1(N__48537),
            .in2(N__45981),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_8 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_7 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_18_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_18_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__45954),
            .in2(N__48327),
            .in3(N__45972),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_9 ),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_18_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_18_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__45933),
            .in2(N__48246),
            .in3(N__45948),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_18_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_18_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__49263),
            .in2(N__45909),
            .in3(N__45927),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_18_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_18_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__45900),
            .in2(N__45873),
            .in3(N__45888),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_18_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_18_17_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_18_17_4  (
            .in0(N__45861),
            .in1(N__45831),
            .in2(N__45846),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_18_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_18_17_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_18_17_5  (
            .in0(N__45825),
            .in1(N__45810),
            .in2(N__45801),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_18_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_18_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__45789),
            .in2(N__46158),
            .in3(N__45780),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_time_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_18_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_18_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__46149),
            .in2(N__46137),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_15 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_18_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_18_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__46122),
            .in2(N__46113),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_18_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_18_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__46098),
            .in2(N__46083),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_18_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_18_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__48231),
            .in2(N__50985),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_18_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_18_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__46065),
            .in2(N__46056),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_18_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_18_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__46044),
            .in2(N__46038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_18_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_18_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__46029),
            .in2(N__46017),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_18_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_18_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__47199),
            .in2(N__47193),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un4_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un4_running_cry_0_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_LUT4_0_LC_18_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_LUT4_0_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_LUT4_0_LC_18_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_LUT4_0_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47181),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_0_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_19_4 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_18_19_4  (
            .in0(N__47107),
            .in1(N__46994),
            .in2(_gnd_net_),
            .in3(N__46975),
            .lcout(\phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50785),
            .ce(),
            .sr(N__50322));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_18_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_18_20_0 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_18_20_0  (
            .in0(N__46719),
            .in1(N__46596),
            .in2(N__46419),
            .in3(N__46956),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50780),
            .ce(),
            .sr(N__50331));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_18_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_18_20_3 .LUT_INIT=16'b1111000001010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_18_20_3  (
            .in0(N__46595),
            .in1(N__46383),
            .in2(N__46908),
            .in3(N__46720),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50780),
            .ce(),
            .sr(N__50331));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_18_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_18_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_18_21_1 .LUT_INIT=16'b1111000011101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_18_21_1  (
            .in0(N__46593),
            .in1(N__46384),
            .in2(N__46848),
            .in3(N__46768),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50773),
            .ce(),
            .sr(N__50337));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_18_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_18_21_4 .LUT_INIT=16'b1111010011100100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_18_21_4  (
            .in0(N__46767),
            .in1(N__46594),
            .in2(N__46434),
            .in3(N__46385),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50773),
            .ce(),
            .sr(N__50337));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_18_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_18_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_18_22_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_18_22_0  (
            .in0(_gnd_net_),
            .in1(N__46203),
            .in2(N__46185),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_18_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_18_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_18_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_18_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_18_22_1  (
            .in0(_gnd_net_),
            .in1(N__47487),
            .in2(N__47469),
            .in3(N__47442),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_18_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_18_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_18_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_18_22_2  (
            .in0(_gnd_net_),
            .in1(N__47439),
            .in2(N__47424),
            .in3(N__47397),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_18_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_18_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_18_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(N__47394),
            .in2(N__47376),
            .in3(N__47349),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_18_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_18_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_18_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_18_22_4  (
            .in0(_gnd_net_),
            .in1(N__47346),
            .in2(N__47608),
            .in3(N__47316),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_18_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_18_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_18_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_18_22_5  (
            .in0(_gnd_net_),
            .in1(N__47313),
            .in2(N__47610),
            .in3(N__47289),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_18_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_18_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_18_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_18_22_6  (
            .in0(_gnd_net_),
            .in1(N__47286),
            .in2(N__47609),
            .in3(N__47262),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_18_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_18_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_18_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_18_22_7  (
            .in0(_gnd_net_),
            .in1(N__47590),
            .in2(N__47259),
            .in3(N__47232),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_18_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_18_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_18_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__47594),
            .in2(N__47229),
            .in3(N__47202),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_18_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_18_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_18_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_18_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_18_23_1  (
            .in0(_gnd_net_),
            .in1(N__47766),
            .in2(N__47611),
            .in3(N__47736),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_18_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_18_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_18_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_18_23_2  (
            .in0(_gnd_net_),
            .in1(N__47598),
            .in2(N__47733),
            .in3(N__47703),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_18_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_18_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_18_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_18_23_3  (
            .in0(_gnd_net_),
            .in1(N__47700),
            .in2(N__47612),
            .in3(N__47676),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_18_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_18_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_18_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__47602),
            .in2(N__47673),
            .in3(N__47643),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_18_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_18_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_18_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_18_23_5  (
            .in0(_gnd_net_),
            .in1(N__47640),
            .in2(N__47613),
            .in3(N__47616),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_18_23_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_18_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_18_23_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__47606),
            .in2(N__47535),
            .in3(N__47505),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_18_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_18_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_18_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_18_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47502),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_6.C_ON=1'b0;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_clock_output_0_THRU_LUT4_0_LC_18_30_6 (
            .in0(N__50919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_clock_output_0_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_20_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_20_6_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_2_LC_20_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_2_LC_20_6_6  (
            .in0(N__48501),
            .in1(N__48525),
            .in2(_gnd_net_),
            .in3(N__51620),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50912),
            .ce(N__48861),
            .sr(N__50236));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_20_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_20_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_20_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_20_7_4  (
            .in0(N__51616),
            .in1(N__48307),
            .in2(_gnd_net_),
            .in3(N__48283),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_20_7_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_20_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_20_7_5  (
            .in0(N__48382),
            .in1(N__48338),
            .in2(_gnd_net_),
            .in3(N__51617),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(elapsed_time_ns_1_RNIL73T9_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_20_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_20_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_9_LC_20_7_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_9_LC_20_7_6  (
            .in0(N__51618),
            .in1(_gnd_net_),
            .in2(N__47922),
            .in3(N__48383),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50911),
            .ce(N__48875),
            .sr(N__50239));
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_20_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_20_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_11_LC_20_8_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_11_LC_20_8_5  (
            .in0(N__49318),
            .in1(N__49301),
            .in2(_gnd_net_),
            .in3(N__51619),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50906),
            .ce(N__48860),
            .sr(N__50243));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_20_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_20_9_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_20_9_0  (
            .in0(N__48454),
            .in1(N__48431),
            .in2(_gnd_net_),
            .in3(N__51430),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_20_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_20_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_20_9_1  (
            .in0(N__49296),
            .in1(N__48282),
            .in2(N__48384),
            .in3(N__47887),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_20_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_20_9_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_20_9_2  (
            .in0(N__47854),
            .in1(N__47819),
            .in2(N__47784),
            .in3(N__48177),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_20_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_20_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_20_9_3  (
            .in0(N__49297),
            .in1(N__51433),
            .in2(_gnd_net_),
            .in3(N__49322),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_20_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_20_9_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_20_9_4  (
            .in0(_gnd_net_),
            .in1(N__48571),
            .in2(_gnd_net_),
            .in3(N__48213),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_20_9_5  (
            .in0(N__48430),
            .in1(N__48492),
            .in2(N__49425),
            .in3(N__48038),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_20_9_6  (
            .in0(_gnd_net_),
            .in1(N__48162),
            .in2(N__48129),
            .in3(N__51694),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_20_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_20_9_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_20_9_7  (
            .in0(N__48572),
            .in1(N__51434),
            .in2(_gnd_net_),
            .in3(N__48592),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_20_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_20_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_20_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_20_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48117),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50893),
            .ce(N__48093),
            .sr(N__50252));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_20_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_20_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_20_10_5  (
            .in0(N__48523),
            .in1(N__48493),
            .in2(_gnd_net_),
            .in3(N__51581),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_20_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_20_10_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_20_10_7  (
            .in0(N__47992),
            .in1(N__48039),
            .in2(_gnd_net_),
            .in3(N__51580),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_20_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_20_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_19_LC_20_11_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_19_LC_20_11_1  (
            .in0(N__49476),
            .in1(N__49497),
            .in2(_gnd_net_),
            .in3(N__51595),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50886),
            .ce(N__48868),
            .sr(N__50260));
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_20_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_20_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_23_LC_20_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_23_LC_20_11_3  (
            .in0(N__51087),
            .in1(N__51127),
            .in2(_gnd_net_),
            .in3(N__51596),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50886),
            .ce(N__48868),
            .sr(N__50260));
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_20_12_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_20_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_8_LC_20_12_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_8_LC_20_12_4  (
            .in0(N__51593),
            .in1(N__48593),
            .in2(_gnd_net_),
            .in3(N__48573),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50876),
            .ce(N__49250),
            .sr(N__50268));
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_20_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_20_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_2_LC_20_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_2_LC_20_12_5  (
            .in0(N__48524),
            .in1(N__51594),
            .in2(_gnd_net_),
            .in3(N__48500),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50876),
            .ce(N__49250),
            .sr(N__50268));
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_20_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_20_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_3_LC_20_12_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_3_LC_20_12_6  (
            .in0(N__51592),
            .in1(N__48455),
            .in2(_gnd_net_),
            .in3(N__48432),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50876),
            .ce(N__49250),
            .sr(N__50268));
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_20_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_20_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_23_LC_20_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_23_LC_20_13_0  (
            .in0(N__51556),
            .in1(N__51082),
            .in2(_gnd_net_),
            .in3(N__51128),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50867),
            .ce(N__49249),
            .sr(N__50274));
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_20_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_20_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_22_LC_20_13_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_22_LC_20_13_2  (
            .in0(N__51716),
            .in1(N__51555),
            .in2(_gnd_net_),
            .in3(N__51765),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50867),
            .ce(N__49249),
            .sr(N__50274));
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_20_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_20_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_9_LC_20_13_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_9_LC_20_13_6  (
            .in0(N__51557),
            .in1(N__48381),
            .in2(_gnd_net_),
            .in3(N__48345),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50867),
            .ce(N__49249),
            .sr(N__50274));
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_20_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_20_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_10_LC_20_13_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_10_LC_20_13_7  (
            .in0(N__48312),
            .in1(N__48285),
            .in2(_gnd_net_),
            .in3(N__51558),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50867),
            .ce(N__49249),
            .sr(N__50274));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_20_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_20_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_20_14_0 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_20_14_0  (
            .in0(N__51065),
            .in1(N__51050),
            .in2(N__51027),
            .in3(N__50996),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_20_14_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_20_14_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_20_14_1 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_20_14_1  (
            .in0(N__49496),
            .in1(N__49474),
            .in2(N__51579),
            .in3(_gnd_net_),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_14_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_14_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_20_14_4  (
            .in0(N__49419),
            .in1(N__51522),
            .in2(_gnd_net_),
            .in3(N__49372),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_20_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_20_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_19_LC_20_15_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_19_LC_20_15_7  (
            .in0(N__49492),
            .in1(N__49475),
            .in2(_gnd_net_),
            .in3(N__51554),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50844),
            .ce(N__49247),
            .sr(N__50292));
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_20_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_20_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_1_LC_20_16_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_1_LC_20_16_2  (
            .in0(N__49420),
            .in1(N__51551),
            .in2(_gnd_net_),
            .in3(N__49373),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50833),
            .ce(N__49246),
            .sr(N__50299));
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_27_LC_20_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_27_LC_20_16_4  (
            .in0(N__51552),
            .in1(N__51696),
            .in2(_gnd_net_),
            .in3(N__51653),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50833),
            .ce(N__49246),
            .sr(N__50299));
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_20_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_20_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.target_time_11_LC_20_16_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_time_11_LC_20_16_7  (
            .in0(N__49323),
            .in1(N__49302),
            .in2(_gnd_net_),
            .in3(N__51553),
            .lcout(\phase_controller_inst2.stoper_hc.target_timeZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50833),
            .ce(N__49246),
            .sr(N__50299));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_20_18_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_20_18_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_20_18_2  (
            .in0(N__49153),
            .in1(N__49206),
            .in2(_gnd_net_),
            .in3(N__51521),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_20_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_20_19_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_20_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49131),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_21_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_21_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.target_time_21_LC_21_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_time_21_LC_21_10_7  (
            .in0(N__51515),
            .in1(N__48963),
            .in2(_gnd_net_),
            .in3(N__48938),
            .lcout(\phase_controller_inst1.stoper_hc.target_timeZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50899),
            .ce(N__48876),
            .sr(N__50261));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_21_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_21_11_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_21_11_3  (
            .in0(N__51715),
            .in1(N__51764),
            .in2(_gnd_net_),
            .in3(N__51503),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_21_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_21_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_21_12_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_21_12_3  (
            .in0(N__51504),
            .in1(N__51695),
            .in2(_gnd_net_),
            .in3(N__51646),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_13_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_21_13_4  (
            .in0(N__51559),
            .in1(N__51086),
            .in2(_gnd_net_),
            .in3(N__51129),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_14_3 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_21_14_3  (
            .in0(N__51066),
            .in1(N__51054),
            .in2(N__51026),
            .in3(N__50997),
            .lcout(\phase_controller_inst2.stoper_hc.un4_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_21_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_21_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_21_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_21_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50966),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50834),
            .ce(),
            .sr(N__50315));
    defparam CONSTANT_ONE_LUT4_LC_22_6_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_22_6_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_22_6_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_22_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // MAIN
