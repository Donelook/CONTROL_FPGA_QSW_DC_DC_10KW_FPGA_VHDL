-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Nov 15 2024 21:13:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "MAIN" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of MAIN
entity MAIN is
port (
    start_stop : in std_logic;
    s2_phy : out std_logic;
    s3_phy : out std_logic;
    il_min_comp2 : in std_logic;
    il_max_comp1 : in std_logic;
    error_pin : in std_logic;
    s1_phy : out std_logic;
    reset : in std_logic;
    il_min_comp1 : in std_logic;
    delay_tr_input : in std_logic;
    s4_phy : out std_logic;
    rgb_g : out std_logic;
    rgb_r : out std_logic;
    rgb_b : out std_logic;
    pwm_output : out std_logic;
    il_max_comp2 : in std_logic;
    delay_hc_input : in std_logic);
end MAIN;

-- Architecture of MAIN
-- View name is \INTERFACE\
architecture \INTERFACE\ of MAIN is

signal \N__50511\ : std_logic;
signal \N__50510\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50499\ : std_logic;
signal \N__50498\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50489\ : std_logic;
signal \N__50482\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50473\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50464\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50462\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50445\ : std_logic;
signal \N__50444\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50436\ : std_logic;
signal \N__50435\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50426\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50410\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50400\ : std_logic;
signal \N__50399\ : std_logic;
signal \N__50382\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50376\ : std_logic;
signal \N__50375\ : std_logic;
signal \N__50372\ : std_logic;
signal \N__50371\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50365\ : std_logic;
signal \N__50362\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50345\ : std_logic;
signal \N__50344\ : std_logic;
signal \N__50341\ : std_logic;
signal \N__50338\ : std_logic;
signal \N__50335\ : std_logic;
signal \N__50332\ : std_logic;
signal \N__50325\ : std_logic;
signal \N__50324\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50320\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50310\ : std_logic;
signal \N__50307\ : std_logic;
signal \N__50304\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50288\ : std_logic;
signal \N__50283\ : std_logic;
signal \N__50280\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50278\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50271\ : std_logic;
signal \N__50268\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50238\ : std_logic;
signal \N__50235\ : std_logic;
signal \N__50234\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50180\ : std_logic;
signal \N__50179\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50177\ : std_logic;
signal \N__50176\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50174\ : std_logic;
signal \N__50173\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50171\ : std_logic;
signal \N__50170\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50168\ : std_logic;
signal \N__50167\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50165\ : std_logic;
signal \N__50164\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50162\ : std_logic;
signal \N__50161\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50159\ : std_logic;
signal \N__50150\ : std_logic;
signal \N__50149\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50147\ : std_logic;
signal \N__50146\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50128\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50105\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50093\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50063\ : std_logic;
signal \N__50060\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50042\ : std_logic;
signal \N__50039\ : std_logic;
signal \N__50036\ : std_logic;
signal \N__50035\ : std_logic;
signal \N__50032\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50022\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50013\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50000\ : std_logic;
signal \N__49995\ : std_logic;
signal \N__49992\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49990\ : std_logic;
signal \N__49987\ : std_logic;
signal \N__49982\ : std_logic;
signal \N__49979\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49973\ : std_logic;
signal \N__49972\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49956\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49953\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49950\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49946\ : std_logic;
signal \N__49945\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49942\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49938\ : std_logic;
signal \N__49937\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49934\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49931\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49928\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49925\ : std_logic;
signal \N__49924\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49922\ : std_logic;
signal \N__49921\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49919\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49916\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49913\ : std_logic;
signal \N__49912\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49907\ : std_logic;
signal \N__49906\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49904\ : std_logic;
signal \N__49903\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49901\ : std_logic;
signal \N__49900\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49898\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49895\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49892\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49889\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49886\ : std_logic;
signal \N__49885\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49882\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49880\ : std_logic;
signal \N__49879\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49877\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49874\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49871\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49868\ : std_logic;
signal \N__49867\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49865\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49862\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49856\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49853\ : std_logic;
signal \N__49852\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49849\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49844\ : std_logic;
signal \N__49843\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49841\ : std_logic;
signal \N__49840\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49838\ : std_logic;
signal \N__49837\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49835\ : std_logic;
signal \N__49834\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49830\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49827\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49824\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49817\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49814\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49811\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49808\ : std_logic;
signal \N__49807\ : std_logic;
signal \N__49806\ : std_logic;
signal \N__49805\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49802\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49482\ : std_logic;
signal \N__49479\ : std_logic;
signal \N__49478\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49473\ : std_logic;
signal \N__49470\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49452\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49446\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49443\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49441\ : std_logic;
signal \N__49440\ : std_logic;
signal \N__49439\ : std_logic;
signal \N__49438\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49436\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49433\ : std_logic;
signal \N__49432\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49425\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49422\ : std_logic;
signal \N__49421\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49419\ : std_logic;
signal \N__49418\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49416\ : std_logic;
signal \N__49415\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49413\ : std_logic;
signal \N__49412\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49410\ : std_logic;
signal \N__49409\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49406\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49403\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49401\ : std_logic;
signal \N__49400\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49398\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49393\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49390\ : std_logic;
signal \N__49389\ : std_logic;
signal \N__49388\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49385\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49381\ : std_logic;
signal \N__49380\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49377\ : std_logic;
signal \N__49376\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49374\ : std_logic;
signal \N__49373\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49371\ : std_logic;
signal \N__49370\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49368\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49365\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49362\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49359\ : std_logic;
signal \N__49358\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49356\ : std_logic;
signal \N__49355\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49353\ : std_logic;
signal \N__49352\ : std_logic;
signal \N__49351\ : std_logic;
signal \N__49350\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49347\ : std_logic;
signal \N__49346\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49343\ : std_logic;
signal \N__49342\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49337\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49334\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49331\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49329\ : std_logic;
signal \N__49328\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49326\ : std_logic;
signal \N__49325\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49322\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49319\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49316\ : std_logic;
signal \N__49315\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49312\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49310\ : std_logic;
signal \N__49309\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49305\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49300\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49297\ : std_logic;
signal \N__49296\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49294\ : std_logic;
signal \N__49293\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49291\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48957\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48952\ : std_logic;
signal \N__48951\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48944\ : std_logic;
signal \N__48941\ : std_logic;
signal \N__48940\ : std_logic;
signal \N__48937\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48933\ : std_logic;
signal \N__48932\ : std_logic;
signal \N__48919\ : std_logic;
signal \N__48916\ : std_logic;
signal \N__48913\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48902\ : std_logic;
signal \N__48899\ : std_logic;
signal \N__48896\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48881\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48869\ : std_logic;
signal \N__48868\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48865\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48861\ : std_logic;
signal \N__48860\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48858\ : std_logic;
signal \N__48857\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48855\ : std_logic;
signal \N__48854\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48852\ : std_logic;
signal \N__48851\ : std_logic;
signal \N__48850\ : std_logic;
signal \N__48849\ : std_logic;
signal \N__48846\ : std_logic;
signal \N__48843\ : std_logic;
signal \N__48840\ : std_logic;
signal \N__48839\ : std_logic;
signal \N__48838\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48836\ : std_logic;
signal \N__48835\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48803\ : std_logic;
signal \N__48800\ : std_logic;
signal \N__48797\ : std_logic;
signal \N__48796\ : std_logic;
signal \N__48793\ : std_logic;
signal \N__48790\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48781\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48775\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48758\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48730\ : std_logic;
signal \N__48729\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48719\ : std_logic;
signal \N__48716\ : std_logic;
signal \N__48713\ : std_logic;
signal \N__48710\ : std_logic;
signal \N__48707\ : std_logic;
signal \N__48704\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48689\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48683\ : std_logic;
signal \N__48680\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48660\ : std_logic;
signal \N__48657\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48648\ : std_logic;
signal \N__48647\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48645\ : std_logic;
signal \N__48644\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48629\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48627\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48625\ : std_logic;
signal \N__48624\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48622\ : std_logic;
signal \N__48619\ : std_logic;
signal \N__48612\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48601\ : std_logic;
signal \N__48592\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48584\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48563\ : std_logic;
signal \N__48552\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48550\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48540\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48523\ : std_logic;
signal \N__48520\ : std_logic;
signal \N__48517\ : std_logic;
signal \N__48514\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48503\ : std_logic;
signal \N__48502\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48491\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48477\ : std_logic;
signal \N__48474\ : std_logic;
signal \N__48471\ : std_logic;
signal \N__48468\ : std_logic;
signal \N__48467\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48460\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48450\ : std_logic;
signal \N__48447\ : std_logic;
signal \N__48442\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48429\ : std_logic;
signal \N__48426\ : std_logic;
signal \N__48425\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48418\ : std_logic;
signal \N__48415\ : std_logic;
signal \N__48412\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48385\ : std_logic;
signal \N__48384\ : std_logic;
signal \N__48381\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48368\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48354\ : std_logic;
signal \N__48353\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48327\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48318\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48313\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48299\ : std_logic;
signal \N__48296\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48277\ : std_logic;
signal \N__48270\ : std_logic;
signal \N__48267\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48261\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48255\ : std_logic;
signal \N__48254\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48252\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48243\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48240\ : std_logic;
signal \N__48239\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48237\ : std_logic;
signal \N__48236\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48234\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48228\ : std_logic;
signal \N__48227\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48215\ : std_logic;
signal \N__48214\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48212\ : std_logic;
signal \N__48211\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48208\ : std_logic;
signal \N__48207\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48186\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48170\ : std_logic;
signal \N__48169\ : std_logic;
signal \N__48168\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48165\ : std_logic;
signal \N__48164\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48154\ : std_logic;
signal \N__48151\ : std_logic;
signal \N__48142\ : std_logic;
signal \N__48127\ : std_logic;
signal \N__48110\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48104\ : std_logic;
signal \N__48101\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48095\ : std_logic;
signal \N__48094\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48092\ : std_logic;
signal \N__48091\ : std_logic;
signal \N__48088\ : std_logic;
signal \N__48087\ : std_logic;
signal \N__48086\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48084\ : std_logic;
signal \N__48083\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48079\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48068\ : std_logic;
signal \N__48061\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48047\ : std_logic;
signal \N__48044\ : std_logic;
signal \N__48031\ : std_logic;
signal \N__48016\ : std_logic;
signal \N__48011\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48008\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__47998\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47969\ : std_logic;
signal \N__47956\ : std_logic;
signal \N__47947\ : std_logic;
signal \N__47940\ : std_logic;
signal \N__47919\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47911\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47901\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47862\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47839\ : std_logic;
signal \N__47838\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47827\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47819\ : std_logic;
signal \N__47818\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47816\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47809\ : std_logic;
signal \N__47808\ : std_logic;
signal \N__47807\ : std_logic;
signal \N__47802\ : std_logic;
signal \N__47801\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47799\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47796\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47792\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47769\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47757\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47751\ : std_logic;
signal \N__47750\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47740\ : std_logic;
signal \N__47739\ : std_logic;
signal \N__47736\ : std_logic;
signal \N__47733\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47722\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47693\ : std_logic;
signal \N__47690\ : std_logic;
signal \N__47689\ : std_logic;
signal \N__47686\ : std_logic;
signal \N__47685\ : std_logic;
signal \N__47682\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47678\ : std_logic;
signal \N__47677\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47670\ : std_logic;
signal \N__47669\ : std_logic;
signal \N__47666\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47661\ : std_logic;
signal \N__47658\ : std_logic;
signal \N__47657\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47642\ : std_logic;
signal \N__47641\ : std_logic;
signal \N__47638\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47624\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47619\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47617\ : std_logic;
signal \N__47616\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47614\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47611\ : std_logic;
signal \N__47610\ : std_logic;
signal \N__47607\ : std_logic;
signal \N__47604\ : std_logic;
signal \N__47597\ : std_logic;
signal \N__47594\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47590\ : std_logic;
signal \N__47589\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47587\ : std_logic;
signal \N__47586\ : std_logic;
signal \N__47585\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47527\ : std_logic;
signal \N__47524\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47473\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47455\ : std_logic;
signal \N__47452\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47429\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47418\ : std_logic;
signal \N__47407\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47395\ : std_logic;
signal \N__47392\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47358\ : std_logic;
signal \N__47355\ : std_logic;
signal \N__47348\ : std_logic;
signal \N__47335\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47294\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47273\ : std_logic;
signal \N__47272\ : std_logic;
signal \N__47269\ : std_logic;
signal \N__47266\ : std_logic;
signal \N__47263\ : std_logic;
signal \N__47260\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47233\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47226\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47205\ : std_logic;
signal \N__47202\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47195\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47189\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47181\ : std_logic;
signal \N__47178\ : std_logic;
signal \N__47175\ : std_logic;
signal \N__47174\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47162\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47160\ : std_logic;
signal \N__47159\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47157\ : std_logic;
signal \N__47156\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47154\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47127\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47121\ : std_logic;
signal \N__47120\ : std_logic;
signal \N__47117\ : std_logic;
signal \N__47114\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47109\ : std_logic;
signal \N__47106\ : std_logic;
signal \N__47103\ : std_logic;
signal \N__47100\ : std_logic;
signal \N__47097\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47089\ : std_logic;
signal \N__47084\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47074\ : std_logic;
signal \N__47071\ : std_logic;
signal \N__47070\ : std_logic;
signal \N__47069\ : std_logic;
signal \N__47064\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47060\ : std_logic;
signal \N__47059\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47047\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47044\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47040\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47035\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47032\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47029\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47026\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47023\ : std_logic;
signal \N__47022\ : std_logic;
signal \N__47021\ : std_logic;
signal \N__47020\ : std_logic;
signal \N__47017\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47000\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46991\ : std_logic;
signal \N__46988\ : std_logic;
signal \N__46979\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46970\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46966\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46964\ : std_logic;
signal \N__46961\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46958\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46955\ : std_logic;
signal \N__46944\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46941\ : std_logic;
signal \N__46940\ : std_logic;
signal \N__46937\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46934\ : std_logic;
signal \N__46933\ : std_logic;
signal \N__46922\ : std_logic;
signal \N__46921\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46919\ : std_logic;
signal \N__46918\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46916\ : std_logic;
signal \N__46915\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46913\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46903\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46889\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46880\ : std_logic;
signal \N__46879\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46874\ : std_logic;
signal \N__46867\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46853\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46850\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46831\ : std_logic;
signal \N__46830\ : std_logic;
signal \N__46827\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46815\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46805\ : std_logic;
signal \N__46798\ : std_logic;
signal \N__46795\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46775\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46749\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46733\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46724\ : std_logic;
signal \N__46723\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46712\ : std_logic;
signal \N__46703\ : std_logic;
signal \N__46696\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46681\ : std_logic;
signal \N__46676\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46653\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46639\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46629\ : std_logic;
signal \N__46626\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46604\ : std_logic;
signal \N__46601\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46595\ : std_logic;
signal \N__46590\ : std_logic;
signal \N__46587\ : std_logic;
signal \N__46584\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46577\ : std_logic;
signal \N__46576\ : std_logic;
signal \N__46573\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46554\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46550\ : std_logic;
signal \N__46547\ : std_logic;
signal \N__46544\ : std_logic;
signal \N__46539\ : std_logic;
signal \N__46536\ : std_logic;
signal \N__46533\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46529\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46499\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46490\ : std_logic;
signal \N__46487\ : std_logic;
signal \N__46484\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46469\ : std_logic;
signal \N__46464\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46460\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46455\ : std_logic;
signal \N__46452\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46440\ : std_logic;
signal \N__46439\ : std_logic;
signal \N__46436\ : std_logic;
signal \N__46433\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46418\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46412\ : std_logic;
signal \N__46411\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46409\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46406\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46359\ : std_logic;
signal \N__46354\ : std_logic;
signal \N__46351\ : std_logic;
signal \N__46348\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46338\ : std_logic;
signal \N__46335\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46319\ : std_logic;
signal \N__46316\ : std_logic;
signal \N__46315\ : std_logic;
signal \N__46310\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46304\ : std_logic;
signal \N__46299\ : std_logic;
signal \N__46296\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46292\ : std_logic;
signal \N__46289\ : std_logic;
signal \N__46286\ : std_logic;
signal \N__46285\ : std_logic;
signal \N__46280\ : std_logic;
signal \N__46277\ : std_logic;
signal \N__46274\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46265\ : std_logic;
signal \N__46260\ : std_logic;
signal \N__46259\ : std_logic;
signal \N__46256\ : std_logic;
signal \N__46253\ : std_logic;
signal \N__46250\ : std_logic;
signal \N__46245\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46238\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46225\ : std_logic;
signal \N__46222\ : std_logic;
signal \N__46217\ : std_logic;
signal \N__46214\ : std_logic;
signal \N__46209\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46196\ : std_logic;
signal \N__46193\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46177\ : std_logic;
signal \N__46170\ : std_logic;
signal \N__46167\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46161\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46157\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46140\ : std_logic;
signal \N__46139\ : std_logic;
signal \N__46136\ : std_logic;
signal \N__46133\ : std_logic;
signal \N__46132\ : std_logic;
signal \N__46127\ : std_logic;
signal \N__46124\ : std_logic;
signal \N__46121\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46113\ : std_logic;
signal \N__46110\ : std_logic;
signal \N__46107\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46103\ : std_logic;
signal \N__46100\ : std_logic;
signal \N__46097\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46085\ : std_logic;
signal \N__46082\ : std_logic;
signal \N__46079\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46073\ : std_logic;
signal \N__46070\ : std_logic;
signal \N__46067\ : std_logic;
signal \N__46062\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46040\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46029\ : std_logic;
signal \N__46026\ : std_logic;
signal \N__46025\ : std_logic;
signal \N__46022\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46002\ : std_logic;
signal \N__45999\ : std_logic;
signal \N__45998\ : std_logic;
signal \N__45997\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45986\ : std_logic;
signal \N__45981\ : std_logic;
signal \N__45978\ : std_logic;
signal \N__45975\ : std_logic;
signal \N__45972\ : std_logic;
signal \N__45971\ : std_logic;
signal \N__45968\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45964\ : std_logic;
signal \N__45961\ : std_logic;
signal \N__45958\ : std_logic;
signal \N__45955\ : std_logic;
signal \N__45952\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45939\ : std_logic;
signal \N__45938\ : std_logic;
signal \N__45935\ : std_logic;
signal \N__45932\ : std_logic;
signal \N__45929\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45925\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45917\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45890\ : std_logic;
signal \N__45887\ : std_logic;
signal \N__45884\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45849\ : std_logic;
signal \N__45846\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45827\ : std_logic;
signal \N__45824\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45815\ : std_logic;
signal \N__45812\ : std_logic;
signal \N__45809\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45803\ : std_logic;
signal \N__45800\ : std_logic;
signal \N__45797\ : std_logic;
signal \N__45794\ : std_logic;
signal \N__45789\ : std_logic;
signal \N__45786\ : std_logic;
signal \N__45785\ : std_logic;
signal \N__45782\ : std_logic;
signal \N__45779\ : std_logic;
signal \N__45774\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45770\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45746\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45740\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45732\ : std_logic;
signal \N__45731\ : std_logic;
signal \N__45726\ : std_logic;
signal \N__45725\ : std_logic;
signal \N__45722\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45716\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45707\ : std_logic;
signal \N__45704\ : std_logic;
signal \N__45701\ : std_logic;
signal \N__45698\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45685\ : std_logic;
signal \N__45682\ : std_logic;
signal \N__45679\ : std_logic;
signal \N__45672\ : std_logic;
signal \N__45669\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45665\ : std_logic;
signal \N__45662\ : std_logic;
signal \N__45659\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45652\ : std_logic;
signal \N__45649\ : std_logic;
signal \N__45646\ : std_logic;
signal \N__45643\ : std_logic;
signal \N__45640\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45623\ : std_logic;
signal \N__45620\ : std_logic;
signal \N__45619\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45603\ : std_logic;
signal \N__45600\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45593\ : std_logic;
signal \N__45590\ : std_logic;
signal \N__45587\ : std_logic;
signal \N__45584\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45564\ : std_logic;
signal \N__45563\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45559\ : std_logic;
signal \N__45556\ : std_logic;
signal \N__45551\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45545\ : std_logic;
signal \N__45544\ : std_logic;
signal \N__45541\ : std_logic;
signal \N__45536\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45515\ : std_logic;
signal \N__45514\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45508\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45493\ : std_logic;
signal \N__45490\ : std_logic;
signal \N__45487\ : std_logic;
signal \N__45484\ : std_logic;
signal \N__45481\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45468\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45430\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45401\ : std_logic;
signal \N__45396\ : std_logic;
signal \N__45393\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45387\ : std_logic;
signal \N__45384\ : std_logic;
signal \N__45383\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45352\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45343\ : std_logic;
signal \N__45342\ : std_logic;
signal \N__45337\ : std_logic;
signal \N__45334\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45321\ : std_logic;
signal \N__45318\ : std_logic;
signal \N__45315\ : std_logic;
signal \N__45312\ : std_logic;
signal \N__45309\ : std_logic;
signal \N__45306\ : std_logic;
signal \N__45305\ : std_logic;
signal \N__45302\ : std_logic;
signal \N__45299\ : std_logic;
signal \N__45296\ : std_logic;
signal \N__45295\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45281\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45272\ : std_logic;
signal \N__45267\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45260\ : std_logic;
signal \N__45257\ : std_logic;
signal \N__45252\ : std_logic;
signal \N__45249\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45225\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45219\ : std_logic;
signal \N__45216\ : std_logic;
signal \N__45213\ : std_logic;
signal \N__45212\ : std_logic;
signal \N__45209\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45199\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45190\ : std_logic;
signal \N__45187\ : std_logic;
signal \N__45184\ : std_logic;
signal \N__45181\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45172\ : std_logic;
signal \N__45167\ : std_logic;
signal \N__45164\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45153\ : std_logic;
signal \N__45150\ : std_logic;
signal \N__45147\ : std_logic;
signal \N__45146\ : std_logic;
signal \N__45143\ : std_logic;
signal \N__45140\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45133\ : std_logic;
signal \N__45130\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45124\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45111\ : std_logic;
signal \N__45108\ : std_logic;
signal \N__45105\ : std_logic;
signal \N__45102\ : std_logic;
signal \N__45099\ : std_logic;
signal \N__45096\ : std_logic;
signal \N__45095\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45056\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45038\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45015\ : std_logic;
signal \N__45014\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45003\ : std_logic;
signal \N__45000\ : std_logic;
signal \N__44997\ : std_logic;
signal \N__44994\ : std_logic;
signal \N__44991\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44980\ : std_logic;
signal \N__44973\ : std_logic;
signal \N__44972\ : std_logic;
signal \N__44969\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44958\ : std_logic;
signal \N__44955\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44947\ : std_logic;
signal \N__44944\ : std_logic;
signal \N__44941\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44927\ : std_logic;
signal \N__44922\ : std_logic;
signal \N__44919\ : std_logic;
signal \N__44916\ : std_logic;
signal \N__44915\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44908\ : std_logic;
signal \N__44905\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44892\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44886\ : std_logic;
signal \N__44883\ : std_logic;
signal \N__44880\ : std_logic;
signal \N__44877\ : std_logic;
signal \N__44874\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44869\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44867\ : std_logic;
signal \N__44866\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44864\ : std_logic;
signal \N__44863\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44852\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44827\ : std_logic;
signal \N__44826\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44824\ : std_logic;
signal \N__44823\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44821\ : std_logic;
signal \N__44820\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44818\ : std_logic;
signal \N__44815\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44797\ : std_logic;
signal \N__44792\ : std_logic;
signal \N__44787\ : std_logic;
signal \N__44778\ : std_logic;
signal \N__44769\ : std_logic;
signal \N__44762\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44752\ : std_logic;
signal \N__44749\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44739\ : std_logic;
signal \N__44736\ : std_logic;
signal \N__44733\ : std_logic;
signal \N__44730\ : std_logic;
signal \N__44729\ : std_logic;
signal \N__44726\ : std_logic;
signal \N__44723\ : std_logic;
signal \N__44720\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44713\ : std_logic;
signal \N__44710\ : std_logic;
signal \N__44707\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44686\ : std_logic;
signal \N__44683\ : std_logic;
signal \N__44680\ : std_logic;
signal \N__44677\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44655\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44612\ : std_logic;
signal \N__44611\ : std_logic;
signal \N__44608\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44599\ : std_logic;
signal \N__44596\ : std_logic;
signal \N__44589\ : std_logic;
signal \N__44588\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44584\ : std_logic;
signal \N__44581\ : std_logic;
signal \N__44578\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44574\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44566\ : std_logic;
signal \N__44563\ : std_logic;
signal \N__44560\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44546\ : std_logic;
signal \N__44545\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44537\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44531\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44525\ : std_logic;
signal \N__44522\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44513\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44507\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44493\ : std_logic;
signal \N__44490\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44478\ : std_logic;
signal \N__44477\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44470\ : std_logic;
signal \N__44465\ : std_logic;
signal \N__44460\ : std_logic;
signal \N__44459\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44452\ : std_logic;
signal \N__44447\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44441\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44430\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44424\ : std_logic;
signal \N__44421\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44417\ : std_logic;
signal \N__44416\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44404\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44398\ : std_logic;
signal \N__44395\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44382\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44376\ : std_logic;
signal \N__44375\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44364\ : std_logic;
signal \N__44363\ : std_logic;
signal \N__44358\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44354\ : std_logic;
signal \N__44351\ : std_logic;
signal \N__44348\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44325\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44321\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44317\ : std_logic;
signal \N__44314\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44288\ : std_logic;
signal \N__44285\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44277\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44267\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44258\ : std_logic;
signal \N__44255\ : std_logic;
signal \N__44252\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44246\ : std_logic;
signal \N__44243\ : std_logic;
signal \N__44240\ : std_logic;
signal \N__44237\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44201\ : std_logic;
signal \N__44198\ : std_logic;
signal \N__44195\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44189\ : std_logic;
signal \N__44186\ : std_logic;
signal \N__44183\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44174\ : std_logic;
signal \N__44171\ : std_logic;
signal \N__44168\ : std_logic;
signal \N__44165\ : std_logic;
signal \N__44162\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44156\ : std_logic;
signal \N__44153\ : std_logic;
signal \N__44150\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44139\ : std_logic;
signal \N__44138\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44125\ : std_logic;
signal \N__44122\ : std_logic;
signal \N__44119\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44103\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44090\ : std_logic;
signal \N__44087\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44075\ : std_logic;
signal \N__44070\ : std_logic;
signal \N__44069\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44063\ : std_logic;
signal \N__44060\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44048\ : std_logic;
signal \N__44045\ : std_logic;
signal \N__44042\ : std_logic;
signal \N__44039\ : std_logic;
signal \N__44034\ : std_logic;
signal \N__44033\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44027\ : std_logic;
signal \N__44024\ : std_logic;
signal \N__44021\ : std_logic;
signal \N__44018\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__43998\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43983\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43976\ : std_logic;
signal \N__43973\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43967\ : std_logic;
signal \N__43964\ : std_logic;
signal \N__43961\ : std_logic;
signal \N__43958\ : std_logic;
signal \N__43953\ : std_logic;
signal \N__43950\ : std_logic;
signal \N__43947\ : std_logic;
signal \N__43946\ : std_logic;
signal \N__43943\ : std_logic;
signal \N__43940\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43934\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43916\ : std_logic;
signal \N__43913\ : std_logic;
signal \N__43910\ : std_logic;
signal \N__43909\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43883\ : std_logic;
signal \N__43880\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43876\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43870\ : std_logic;
signal \N__43867\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43838\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43824\ : std_logic;
signal \N__43823\ : std_logic;
signal \N__43820\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43809\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43805\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43779\ : std_logic;
signal \N__43776\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43763\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43757\ : std_logic;
signal \N__43754\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43742\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43736\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43730\ : std_logic;
signal \N__43727\ : std_logic;
signal \N__43724\ : std_logic;
signal \N__43719\ : std_logic;
signal \N__43716\ : std_logic;
signal \N__43715\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43706\ : std_logic;
signal \N__43703\ : std_logic;
signal \N__43700\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43691\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43682\ : std_logic;
signal \N__43679\ : std_logic;
signal \N__43676\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43668\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43654\ : std_logic;
signal \N__43649\ : std_logic;
signal \N__43646\ : std_logic;
signal \N__43643\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43634\ : std_logic;
signal \N__43631\ : std_logic;
signal \N__43628\ : std_logic;
signal \N__43625\ : std_logic;
signal \N__43622\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43604\ : std_logic;
signal \N__43599\ : std_logic;
signal \N__43596\ : std_logic;
signal \N__43593\ : std_logic;
signal \N__43592\ : std_logic;
signal \N__43589\ : std_logic;
signal \N__43586\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43565\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43536\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43510\ : std_logic;
signal \N__43507\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43494\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43485\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43480\ : std_logic;
signal \N__43477\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43470\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43459\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43449\ : std_logic;
signal \N__43448\ : std_logic;
signal \N__43445\ : std_logic;
signal \N__43442\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43429\ : std_logic;
signal \N__43426\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43407\ : std_logic;
signal \N__43404\ : std_logic;
signal \N__43401\ : std_logic;
signal \N__43398\ : std_logic;
signal \N__43395\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43386\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43372\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43368\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43349\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43343\ : std_logic;
signal \N__43340\ : std_logic;
signal \N__43337\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43327\ : std_logic;
signal \N__43324\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43314\ : std_logic;
signal \N__43311\ : std_logic;
signal \N__43308\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43302\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43298\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43289\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43283\ : std_logic;
signal \N__43280\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43266\ : std_logic;
signal \N__43263\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43256\ : std_logic;
signal \N__43253\ : std_logic;
signal \N__43250\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43240\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43233\ : std_logic;
signal \N__43230\ : std_logic;
signal \N__43227\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43191\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43163\ : std_logic;
signal \N__43160\ : std_logic;
signal \N__43157\ : std_logic;
signal \N__43154\ : std_logic;
signal \N__43151\ : std_logic;
signal \N__43150\ : std_logic;
signal \N__43147\ : std_logic;
signal \N__43144\ : std_logic;
signal \N__43141\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43132\ : std_logic;
signal \N__43129\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43103\ : std_logic;
signal \N__43102\ : std_logic;
signal \N__43099\ : std_logic;
signal \N__43096\ : std_logic;
signal \N__43093\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43084\ : std_logic;
signal \N__43081\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43061\ : std_logic;
signal \N__43058\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43052\ : std_logic;
signal \N__43049\ : std_logic;
signal \N__43048\ : std_logic;
signal \N__43043\ : std_logic;
signal \N__43040\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43036\ : std_logic;
signal \N__43033\ : std_logic;
signal \N__43030\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43013\ : std_logic;
signal \N__43010\ : std_logic;
signal \N__43007\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43001\ : std_logic;
signal \N__42998\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42987\ : std_logic;
signal \N__42984\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42959\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42953\ : std_logic;
signal \N__42950\ : std_logic;
signal \N__42947\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42908\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42902\ : std_logic;
signal \N__42897\ : std_logic;
signal \N__42896\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42866\ : std_logic;
signal \N__42863\ : std_logic;
signal \N__42860\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42853\ : std_logic;
signal \N__42850\ : std_logic;
signal \N__42845\ : std_logic;
signal \N__42844\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42838\ : std_logic;
signal \N__42835\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42818\ : std_logic;
signal \N__42817\ : std_logic;
signal \N__42814\ : std_logic;
signal \N__42811\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42799\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42791\ : std_logic;
signal \N__42786\ : std_logic;
signal \N__42783\ : std_logic;
signal \N__42780\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42757\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42745\ : std_logic;
signal \N__42742\ : std_logic;
signal \N__42739\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42731\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42723\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42714\ : std_logic;
signal \N__42713\ : std_logic;
signal \N__42710\ : std_logic;
signal \N__42707\ : std_logic;
signal \N__42704\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42688\ : std_logic;
signal \N__42687\ : std_logic;
signal \N__42684\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42676\ : std_logic;
signal \N__42669\ : std_logic;
signal \N__42666\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42660\ : std_logic;
signal \N__42657\ : std_logic;
signal \N__42656\ : std_logic;
signal \N__42653\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42647\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42631\ : std_logic;
signal \N__42628\ : std_logic;
signal \N__42621\ : std_logic;
signal \N__42618\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42602\ : std_logic;
signal \N__42599\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42589\ : std_logic;
signal \N__42586\ : std_logic;
signal \N__42583\ : std_logic;
signal \N__42580\ : std_logic;
signal \N__42573\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42564\ : std_logic;
signal \N__42561\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42552\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42525\ : std_logic;
signal \N__42522\ : std_logic;
signal \N__42519\ : std_logic;
signal \N__42516\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42512\ : std_logic;
signal \N__42509\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42499\ : std_logic;
signal \N__42492\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42485\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42479\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42473\ : std_logic;
signal \N__42470\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42462\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42457\ : std_logic;
signal \N__42454\ : std_logic;
signal \N__42451\ : std_logic;
signal \N__42448\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42442\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42418\ : std_logic;
signal \N__42415\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42406\ : std_logic;
signal \N__42401\ : std_logic;
signal \N__42398\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42389\ : std_logic;
signal \N__42388\ : std_logic;
signal \N__42385\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42379\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42362\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42352\ : std_logic;
signal \N__42349\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42337\ : std_logic;
signal \N__42334\ : std_logic;
signal \N__42331\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42314\ : std_logic;
signal \N__42311\ : std_logic;
signal \N__42310\ : std_logic;
signal \N__42307\ : std_logic;
signal \N__42304\ : std_logic;
signal \N__42301\ : std_logic;
signal \N__42298\ : std_logic;
signal \N__42295\ : std_logic;
signal \N__42292\ : std_logic;
signal \N__42289\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42275\ : std_logic;
signal \N__42272\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42245\ : std_logic;
signal \N__42242\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42222\ : std_logic;
signal \N__42219\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42211\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42193\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42152\ : std_logic;
signal \N__42149\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42137\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42133\ : std_logic;
signal \N__42130\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42124\ : std_logic;
signal \N__42121\ : std_logic;
signal \N__42118\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42089\ : std_logic;
signal \N__42086\ : std_logic;
signal \N__42085\ : std_logic;
signal \N__42082\ : std_logic;
signal \N__42079\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42073\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42053\ : std_logic;
signal \N__42050\ : std_logic;
signal \N__42047\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42040\ : std_logic;
signal \N__42037\ : std_logic;
signal \N__42034\ : std_logic;
signal \N__42031\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42002\ : std_logic;
signal \N__41999\ : std_logic;
signal \N__41996\ : std_logic;
signal \N__41995\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41986\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41972\ : std_logic;
signal \N__41969\ : std_logic;
signal \N__41966\ : std_logic;
signal \N__41965\ : std_logic;
signal \N__41960\ : std_logic;
signal \N__41957\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41936\ : std_logic;
signal \N__41935\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41879\ : std_logic;
signal \N__41876\ : std_logic;
signal \N__41873\ : std_logic;
signal \N__41870\ : std_logic;
signal \N__41867\ : std_logic;
signal \N__41864\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41837\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41828\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41824\ : std_logic;
signal \N__41821\ : std_logic;
signal \N__41818\ : std_logic;
signal \N__41815\ : std_logic;
signal \N__41812\ : std_logic;
signal \N__41809\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41799\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41793\ : std_logic;
signal \N__41790\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41784\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41774\ : std_logic;
signal \N__41771\ : std_logic;
signal \N__41768\ : std_logic;
signal \N__41767\ : std_logic;
signal \N__41762\ : std_logic;
signal \N__41759\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41737\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41727\ : std_logic;
signal \N__41724\ : std_logic;
signal \N__41721\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41716\ : std_logic;
signal \N__41713\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41696\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41687\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41677\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41673\ : std_logic;
signal \N__41670\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41651\ : std_logic;
signal \N__41648\ : std_logic;
signal \N__41645\ : std_logic;
signal \N__41640\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41634\ : std_logic;
signal \N__41631\ : std_logic;
signal \N__41630\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41624\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41620\ : std_logic;
signal \N__41617\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41604\ : std_logic;
signal \N__41601\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41597\ : std_logic;
signal \N__41594\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41570\ : std_logic;
signal \N__41567\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41559\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41550\ : std_logic;
signal \N__41547\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41533\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41525\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41519\ : std_logic;
signal \N__41514\ : std_logic;
signal \N__41513\ : std_logic;
signal \N__41510\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41496\ : std_logic;
signal \N__41493\ : std_logic;
signal \N__41490\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41474\ : std_logic;
signal \N__41471\ : std_logic;
signal \N__41468\ : std_logic;
signal \N__41465\ : std_logic;
signal \N__41462\ : std_logic;
signal \N__41461\ : std_logic;
signal \N__41456\ : std_logic;
signal \N__41453\ : std_logic;
signal \N__41450\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41432\ : std_logic;
signal \N__41431\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41418\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41408\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41395\ : std_logic;
signal \N__41392\ : std_logic;
signal \N__41389\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41374\ : std_logic;
signal \N__41371\ : std_logic;
signal \N__41368\ : std_logic;
signal \N__41367\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41359\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41353\ : std_logic;
signal \N__41350\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41341\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41332\ : std_logic;
signal \N__41329\ : std_logic;
signal \N__41326\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41308\ : std_logic;
signal \N__41305\ : std_logic;
signal \N__41302\ : std_logic;
signal \N__41299\ : std_logic;
signal \N__41294\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41279\ : std_logic;
signal \N__41278\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41276\ : std_logic;
signal \N__41275\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41273\ : std_logic;
signal \N__41272\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41270\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41264\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41254\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41252\ : std_logic;
signal \N__41251\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41249\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41246\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41243\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41226\ : std_logic;
signal \N__41223\ : std_logic;
signal \N__41216\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41214\ : std_logic;
signal \N__41213\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41211\ : std_logic;
signal \N__41208\ : std_logic;
signal \N__41199\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41181\ : std_logic;
signal \N__41178\ : std_logic;
signal \N__41175\ : std_logic;
signal \N__41172\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41144\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41124\ : std_logic;
signal \N__41121\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41091\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41085\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41077\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41069\ : std_logic;
signal \N__41066\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41057\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41042\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41024\ : std_logic;
signal \N__41023\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41001\ : std_logic;
signal \N__40998\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40996\ : std_logic;
signal \N__40993\ : std_logic;
signal \N__40988\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40976\ : std_logic;
signal \N__40971\ : std_logic;
signal \N__40968\ : std_logic;
signal \N__40965\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40960\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40951\ : std_logic;
signal \N__40948\ : std_logic;
signal \N__40947\ : std_logic;
signal \N__40940\ : std_logic;
signal \N__40937\ : std_logic;
signal \N__40934\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40921\ : std_logic;
signal \N__40918\ : std_logic;
signal \N__40915\ : std_logic;
signal \N__40912\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40890\ : std_logic;
signal \N__40887\ : std_logic;
signal \N__40884\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40866\ : std_logic;
signal \N__40863\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40846\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40835\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40817\ : std_logic;
signal \N__40814\ : std_logic;
signal \N__40811\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40802\ : std_logic;
signal \N__40799\ : std_logic;
signal \N__40796\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40787\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40761\ : std_logic;
signal \N__40758\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40746\ : std_logic;
signal \N__40743\ : std_logic;
signal \N__40740\ : std_logic;
signal \N__40737\ : std_logic;
signal \N__40734\ : std_logic;
signal \N__40733\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40727\ : std_logic;
signal \N__40724\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40713\ : std_logic;
signal \N__40710\ : std_logic;
signal \N__40709\ : std_logic;
signal \N__40704\ : std_logic;
signal \N__40703\ : std_logic;
signal \N__40700\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40694\ : std_logic;
signal \N__40689\ : std_logic;
signal \N__40686\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40682\ : std_logic;
signal \N__40679\ : std_logic;
signal \N__40676\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40667\ : std_logic;
signal \N__40664\ : std_logic;
signal \N__40661\ : std_logic;
signal \N__40656\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40652\ : std_logic;
signal \N__40649\ : std_logic;
signal \N__40646\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40637\ : std_logic;
signal \N__40634\ : std_logic;
signal \N__40631\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40622\ : std_logic;
signal \N__40619\ : std_logic;
signal \N__40616\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40607\ : std_logic;
signal \N__40604\ : std_logic;
signal \N__40601\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40592\ : std_logic;
signal \N__40589\ : std_logic;
signal \N__40586\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40577\ : std_logic;
signal \N__40574\ : std_logic;
signal \N__40571\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40562\ : std_logic;
signal \N__40559\ : std_logic;
signal \N__40556\ : std_logic;
signal \N__40553\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40549\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40525\ : std_logic;
signal \N__40518\ : std_logic;
signal \N__40515\ : std_logic;
signal \N__40512\ : std_logic;
signal \N__40509\ : std_logic;
signal \N__40506\ : std_logic;
signal \N__40503\ : std_logic;
signal \N__40500\ : std_logic;
signal \N__40497\ : std_logic;
signal \N__40494\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40478\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40469\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40454\ : std_logic;
signal \N__40451\ : std_logic;
signal \N__40448\ : std_logic;
signal \N__40445\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40436\ : std_logic;
signal \N__40433\ : std_logic;
signal \N__40430\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40418\ : std_logic;
signal \N__40415\ : std_logic;
signal \N__40414\ : std_logic;
signal \N__40411\ : std_logic;
signal \N__40408\ : std_logic;
signal \N__40405\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40394\ : std_logic;
signal \N__40391\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40325\ : std_logic;
signal \N__40324\ : std_logic;
signal \N__40321\ : std_logic;
signal \N__40318\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40309\ : std_logic;
signal \N__40306\ : std_logic;
signal \N__40303\ : std_logic;
signal \N__40298\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40249\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40237\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40217\ : std_logic;
signal \N__40214\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40207\ : std_logic;
signal \N__40204\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40166\ : std_logic;
signal \N__40163\ : std_logic;
signal \N__40160\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40142\ : std_logic;
signal \N__40139\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40095\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40081\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40075\ : std_logic;
signal \N__40072\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40050\ : std_logic;
signal \N__40047\ : std_logic;
signal \N__40044\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40031\ : std_logic;
signal \N__40028\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39984\ : std_logic;
signal \N__39981\ : std_logic;
signal \N__39978\ : std_logic;
signal \N__39975\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39969\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39876\ : std_logic;
signal \N__39873\ : std_logic;
signal \N__39870\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39861\ : std_logic;
signal \N__39858\ : std_logic;
signal \N__39855\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39846\ : std_logic;
signal \N__39843\ : std_logic;
signal \N__39840\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39831\ : std_logic;
signal \N__39828\ : std_logic;
signal \N__39825\ : std_logic;
signal \N__39822\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39777\ : std_logic;
signal \N__39774\ : std_logic;
signal \N__39771\ : std_logic;
signal \N__39768\ : std_logic;
signal \N__39765\ : std_logic;
signal \N__39762\ : std_logic;
signal \N__39759\ : std_logic;
signal \N__39756\ : std_logic;
signal \N__39753\ : std_logic;
signal \N__39750\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39741\ : std_logic;
signal \N__39738\ : std_logic;
signal \N__39735\ : std_logic;
signal \N__39732\ : std_logic;
signal \N__39729\ : std_logic;
signal \N__39726\ : std_logic;
signal \N__39723\ : std_logic;
signal \N__39720\ : std_logic;
signal \N__39717\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39708\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39694\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39685\ : std_logic;
signal \N__39682\ : std_logic;
signal \N__39679\ : std_logic;
signal \N__39676\ : std_logic;
signal \N__39673\ : std_logic;
signal \N__39670\ : std_logic;
signal \N__39667\ : std_logic;
signal \N__39664\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39648\ : std_logic;
signal \N__39645\ : std_logic;
signal \N__39642\ : std_logic;
signal \N__39639\ : std_logic;
signal \N__39636\ : std_logic;
signal \N__39633\ : std_logic;
signal \N__39626\ : std_logic;
signal \N__39623\ : std_logic;
signal \N__39620\ : std_logic;
signal \N__39615\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39600\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39592\ : std_logic;
signal \N__39589\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39581\ : std_logic;
signal \N__39578\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39562\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39550\ : std_logic;
signal \N__39543\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39534\ : std_logic;
signal \N__39533\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39525\ : std_logic;
signal \N__39522\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39507\ : std_logic;
signal \N__39504\ : std_logic;
signal \N__39501\ : std_logic;
signal \N__39498\ : std_logic;
signal \N__39495\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39461\ : std_logic;
signal \N__39460\ : std_logic;
signal \N__39457\ : std_logic;
signal \N__39454\ : std_logic;
signal \N__39451\ : std_logic;
signal \N__39450\ : std_logic;
signal \N__39447\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39423\ : std_logic;
signal \N__39420\ : std_logic;
signal \N__39417\ : std_logic;
signal \N__39414\ : std_logic;
signal \N__39411\ : std_logic;
signal \N__39408\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39399\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39371\ : std_logic;
signal \N__39370\ : std_logic;
signal \N__39365\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39352\ : std_logic;
signal \N__39349\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39343\ : std_logic;
signal \N__39338\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39321\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39310\ : std_logic;
signal \N__39307\ : std_logic;
signal \N__39304\ : std_logic;
signal \N__39301\ : std_logic;
signal \N__39298\ : std_logic;
signal \N__39295\ : std_logic;
signal \N__39292\ : std_logic;
signal \N__39289\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39279\ : std_logic;
signal \N__39276\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39268\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39264\ : std_logic;
signal \N__39261\ : std_logic;
signal \N__39258\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39252\ : std_logic;
signal \N__39247\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39234\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39228\ : std_logic;
signal \N__39225\ : std_logic;
signal \N__39222\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39216\ : std_logic;
signal \N__39213\ : std_logic;
signal \N__39210\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39201\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39192\ : std_logic;
signal \N__39189\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39135\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39129\ : std_logic;
signal \N__39126\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39111\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39090\ : std_logic;
signal \N__39087\ : std_logic;
signal \N__39084\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39078\ : std_logic;
signal \N__39075\ : std_logic;
signal \N__39072\ : std_logic;
signal \N__39069\ : std_logic;
signal \N__39066\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39062\ : std_logic;
signal \N__39061\ : std_logic;
signal \N__39060\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39052\ : std_logic;
signal \N__39047\ : std_logic;
signal \N__39044\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39035\ : std_logic;
signal \N__39030\ : std_logic;
signal \N__39027\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39020\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38984\ : std_logic;
signal \N__38981\ : std_logic;
signal \N__38980\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38910\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38901\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38895\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38889\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38883\ : std_logic;
signal \N__38880\ : std_logic;
signal \N__38877\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38871\ : std_logic;
signal \N__38868\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38861\ : std_logic;
signal \N__38860\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38858\ : std_logic;
signal \N__38857\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38854\ : std_logic;
signal \N__38853\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38850\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38828\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38824\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38816\ : std_logic;
signal \N__38815\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38811\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38804\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38800\ : std_logic;
signal \N__38793\ : std_logic;
signal \N__38778\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38762\ : std_logic;
signal \N__38761\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38758\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38755\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38749\ : std_logic;
signal \N__38748\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38746\ : std_logic;
signal \N__38743\ : std_logic;
signal \N__38740\ : std_logic;
signal \N__38737\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38728\ : std_logic;
signal \N__38725\ : std_logic;
signal \N__38724\ : std_logic;
signal \N__38721\ : std_logic;
signal \N__38718\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38710\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38708\ : std_logic;
signal \N__38707\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38689\ : std_logic;
signal \N__38686\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38681\ : std_logic;
signal \N__38680\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38678\ : std_logic;
signal \N__38677\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38672\ : std_logic;
signal \N__38671\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38630\ : std_logic;
signal \N__38627\ : std_logic;
signal \N__38622\ : std_logic;
signal \N__38619\ : std_logic;
signal \N__38602\ : std_logic;
signal \N__38599\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38572\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38556\ : std_logic;
signal \N__38553\ : std_logic;
signal \N__38548\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38531\ : std_logic;
signal \N__38528\ : std_logic;
signal \N__38525\ : std_logic;
signal \N__38516\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38495\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38492\ : std_logic;
signal \N__38491\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38489\ : std_logic;
signal \N__38486\ : std_logic;
signal \N__38485\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38471\ : std_logic;
signal \N__38468\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38462\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38459\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38456\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38449\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38432\ : std_logic;
signal \N__38431\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38428\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38393\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38365\ : std_logic;
signal \N__38358\ : std_logic;
signal \N__38349\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38335\ : std_logic;
signal \N__38332\ : std_logic;
signal \N__38327\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38321\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38310\ : std_logic;
signal \N__38307\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38280\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38271\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38265\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38249\ : std_logic;
signal \N__38244\ : std_logic;
signal \N__38241\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38235\ : std_logic;
signal \N__38226\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38205\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38199\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38187\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38181\ : std_logic;
signal \N__38178\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38160\ : std_logic;
signal \N__38157\ : std_logic;
signal \N__38154\ : std_logic;
signal \N__38151\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38145\ : std_logic;
signal \N__38142\ : std_logic;
signal \N__38139\ : std_logic;
signal \N__38136\ : std_logic;
signal \N__38133\ : std_logic;
signal \N__38130\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38058\ : std_logic;
signal \N__38055\ : std_logic;
signal \N__38052\ : std_logic;
signal \N__38049\ : std_logic;
signal \N__38046\ : std_logic;
signal \N__38043\ : std_logic;
signal \N__38040\ : std_logic;
signal \N__38037\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37929\ : std_logic;
signal \N__37926\ : std_logic;
signal \N__37923\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37900\ : std_logic;
signal \N__37897\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37886\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37857\ : std_logic;
signal \N__37854\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37842\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37830\ : std_logic;
signal \N__37829\ : std_logic;
signal \N__37826\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37818\ : std_logic;
signal \N__37815\ : std_logic;
signal \N__37812\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37800\ : std_logic;
signal \N__37797\ : std_logic;
signal \N__37794\ : std_logic;
signal \N__37791\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37773\ : std_logic;
signal \N__37770\ : std_logic;
signal \N__37767\ : std_logic;
signal \N__37764\ : std_logic;
signal \N__37761\ : std_logic;
signal \N__37758\ : std_logic;
signal \N__37757\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37753\ : std_logic;
signal \N__37748\ : std_logic;
signal \N__37745\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37737\ : std_logic;
signal \N__37736\ : std_logic;
signal \N__37733\ : std_logic;
signal \N__37732\ : std_logic;
signal \N__37727\ : std_logic;
signal \N__37724\ : std_logic;
signal \N__37721\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37704\ : std_logic;
signal \N__37703\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37692\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37680\ : std_logic;
signal \N__37679\ : std_logic;
signal \N__37676\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37638\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37634\ : std_logic;
signal \N__37631\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37626\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37624\ : std_logic;
signal \N__37623\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37621\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37619\ : std_logic;
signal \N__37616\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37612\ : std_logic;
signal \N__37611\ : std_logic;
signal \N__37610\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37608\ : std_logic;
signal \N__37607\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37601\ : std_logic;
signal \N__37598\ : std_logic;
signal \N__37597\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37591\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37588\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37586\ : std_logic;
signal \N__37585\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37568\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37558\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37556\ : std_logic;
signal \N__37555\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37543\ : std_logic;
signal \N__37534\ : std_logic;
signal \N__37531\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37520\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37510\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37508\ : std_logic;
signal \N__37507\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37496\ : std_logic;
signal \N__37487\ : std_logic;
signal \N__37478\ : std_logic;
signal \N__37469\ : std_logic;
signal \N__37460\ : std_logic;
signal \N__37457\ : std_logic;
signal \N__37454\ : std_logic;
signal \N__37451\ : std_logic;
signal \N__37448\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37442\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37430\ : std_logic;
signal \N__37427\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37409\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37397\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37337\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37328\ : std_logic;
signal \N__37327\ : std_logic;
signal \N__37324\ : std_logic;
signal \N__37319\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37313\ : std_logic;
signal \N__37310\ : std_logic;
signal \N__37307\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37298\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37289\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37262\ : std_logic;
signal \N__37259\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37249\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37241\ : std_logic;
signal \N__37238\ : std_logic;
signal \N__37235\ : std_logic;
signal \N__37232\ : std_logic;
signal \N__37229\ : std_logic;
signal \N__37226\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37220\ : std_logic;
signal \N__37217\ : std_logic;
signal \N__37214\ : std_logic;
signal \N__37211\ : std_logic;
signal \N__37208\ : std_logic;
signal \N__37205\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37199\ : std_logic;
signal \N__37198\ : std_logic;
signal \N__37195\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37184\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37178\ : std_logic;
signal \N__37177\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37163\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37151\ : std_logic;
signal \N__37146\ : std_logic;
signal \N__37143\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37134\ : std_logic;
signal \N__37131\ : std_logic;
signal \N__37130\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37115\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37101\ : std_logic;
signal \N__37098\ : std_logic;
signal \N__37095\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37080\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37067\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37052\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37044\ : std_logic;
signal \N__37041\ : std_logic;
signal \N__37040\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37034\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37026\ : std_logic;
signal \N__37023\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37012\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37010\ : std_logic;
signal \N__37007\ : std_logic;
signal \N__37004\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36980\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36953\ : std_logic;
signal \N__36950\ : std_logic;
signal \N__36945\ : std_logic;
signal \N__36942\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36936\ : std_logic;
signal \N__36933\ : std_logic;
signal \N__36930\ : std_logic;
signal \N__36927\ : std_logic;
signal \N__36924\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36915\ : std_logic;
signal \N__36912\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36910\ : std_logic;
signal \N__36907\ : std_logic;
signal \N__36902\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36893\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36875\ : std_logic;
signal \N__36872\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36864\ : std_logic;
signal \N__36861\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36852\ : std_logic;
signal \N__36849\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36813\ : std_logic;
signal \N__36810\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36794\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36788\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36782\ : std_logic;
signal \N__36779\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36773\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36763\ : std_logic;
signal \N__36762\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36733\ : std_logic;
signal \N__36728\ : std_logic;
signal \N__36723\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36720\ : std_logic;
signal \N__36719\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36712\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36705\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36702\ : std_logic;
signal \N__36701\ : std_logic;
signal \N__36700\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36692\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36687\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36681\ : std_logic;
signal \N__36680\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36674\ : std_logic;
signal \N__36673\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36671\ : std_logic;
signal \N__36670\ : std_logic;
signal \N__36667\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36659\ : std_logic;
signal \N__36652\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36649\ : std_logic;
signal \N__36646\ : std_logic;
signal \N__36645\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36633\ : std_logic;
signal \N__36632\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36630\ : std_logic;
signal \N__36625\ : std_logic;
signal \N__36620\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36610\ : std_logic;
signal \N__36607\ : std_logic;
signal \N__36604\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36602\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36597\ : std_logic;
signal \N__36594\ : std_logic;
signal \N__36591\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36562\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36559\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36556\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36550\ : std_logic;
signal \N__36547\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36544\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36542\ : std_logic;
signal \N__36539\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36518\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36506\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36498\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36479\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36470\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36467\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36464\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36457\ : std_logic;
signal \N__36454\ : std_logic;
signal \N__36451\ : std_logic;
signal \N__36446\ : std_logic;
signal \N__36439\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36418\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36416\ : std_logic;
signal \N__36415\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36413\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36410\ : std_logic;
signal \N__36409\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36407\ : std_logic;
signal \N__36406\ : std_logic;
signal \N__36401\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36371\ : std_logic;
signal \N__36368\ : std_logic;
signal \N__36365\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36341\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36284\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36264\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36231\ : std_logic;
signal \N__36230\ : std_logic;
signal \N__36227\ : std_logic;
signal \N__36224\ : std_logic;
signal \N__36223\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36217\ : std_logic;
signal \N__36214\ : std_logic;
signal \N__36209\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36197\ : std_logic;
signal \N__36196\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36184\ : std_logic;
signal \N__36177\ : std_logic;
signal \N__36174\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36156\ : std_logic;
signal \N__36153\ : std_logic;
signal \N__36150\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36138\ : std_logic;
signal \N__36135\ : std_logic;
signal \N__36132\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36111\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36102\ : std_logic;
signal \N__36099\ : std_logic;
signal \N__36096\ : std_logic;
signal \N__36093\ : std_logic;
signal \N__36090\ : std_logic;
signal \N__36087\ : std_logic;
signal \N__36084\ : std_logic;
signal \N__36081\ : std_logic;
signal \N__36078\ : std_logic;
signal \N__36075\ : std_logic;
signal \N__36072\ : std_logic;
signal \N__36069\ : std_logic;
signal \N__36066\ : std_logic;
signal \N__36063\ : std_logic;
signal \N__36060\ : std_logic;
signal \N__36057\ : std_logic;
signal \N__36054\ : std_logic;
signal \N__36051\ : std_logic;
signal \N__36048\ : std_logic;
signal \N__36045\ : std_logic;
signal \N__36042\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36027\ : std_logic;
signal \N__36024\ : std_logic;
signal \N__36021\ : std_logic;
signal \N__36018\ : std_logic;
signal \N__36015\ : std_logic;
signal \N__36012\ : std_logic;
signal \N__36009\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35994\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35976\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35970\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35946\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35940\ : std_logic;
signal \N__35937\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35931\ : std_logic;
signal \N__35928\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35913\ : std_logic;
signal \N__35910\ : std_logic;
signal \N__35907\ : std_logic;
signal \N__35904\ : std_logic;
signal \N__35901\ : std_logic;
signal \N__35898\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35883\ : std_logic;
signal \N__35880\ : std_logic;
signal \N__35877\ : std_logic;
signal \N__35874\ : std_logic;
signal \N__35871\ : std_logic;
signal \N__35868\ : std_logic;
signal \N__35865\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35859\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35850\ : std_logic;
signal \N__35847\ : std_logic;
signal \N__35844\ : std_logic;
signal \N__35841\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35817\ : std_logic;
signal \N__35814\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35805\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35793\ : std_logic;
signal \N__35790\ : std_logic;
signal \N__35787\ : std_logic;
signal \N__35784\ : std_logic;
signal \N__35781\ : std_logic;
signal \N__35778\ : std_logic;
signal \N__35775\ : std_logic;
signal \N__35772\ : std_logic;
signal \N__35769\ : std_logic;
signal \N__35766\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35760\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35730\ : std_logic;
signal \N__35727\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35721\ : std_logic;
signal \N__35718\ : std_logic;
signal \N__35717\ : std_logic;
signal \N__35714\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35706\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35702\ : std_logic;
signal \N__35699\ : std_logic;
signal \N__35696\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35679\ : std_logic;
signal \N__35678\ : std_logic;
signal \N__35675\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35669\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35660\ : std_logic;
signal \N__35657\ : std_logic;
signal \N__35656\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35643\ : std_logic;
signal \N__35638\ : std_logic;
signal \N__35635\ : std_logic;
signal \N__35632\ : std_logic;
signal \N__35629\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35621\ : std_logic;
signal \N__35620\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35606\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35582\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35565\ : std_logic;
signal \N__35562\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35539\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35528\ : std_logic;
signal \N__35523\ : std_logic;
signal \N__35520\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35507\ : std_logic;
signal \N__35506\ : std_logic;
signal \N__35503\ : std_logic;
signal \N__35500\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35478\ : std_logic;
signal \N__35477\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35412\ : std_logic;
signal \N__35409\ : std_logic;
signal \N__35406\ : std_logic;
signal \N__35403\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35390\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35379\ : std_logic;
signal \N__35376\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35372\ : std_logic;
signal \N__35371\ : std_logic;
signal \N__35366\ : std_logic;
signal \N__35363\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35355\ : std_logic;
signal \N__35352\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35342\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35333\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35318\ : std_logic;
signal \N__35315\ : std_logic;
signal \N__35312\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35285\ : std_logic;
signal \N__35282\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35262\ : std_logic;
signal \N__35259\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35223\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35210\ : std_logic;
signal \N__35207\ : std_logic;
signal \N__35204\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35196\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35180\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35169\ : std_logic;
signal \N__35166\ : std_logic;
signal \N__35165\ : std_logic;
signal \N__35162\ : std_logic;
signal \N__35159\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35150\ : std_logic;
signal \N__35147\ : std_logic;
signal \N__35144\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35135\ : std_logic;
signal \N__35132\ : std_logic;
signal \N__35129\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35120\ : std_logic;
signal \N__35117\ : std_logic;
signal \N__35114\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35105\ : std_logic;
signal \N__35102\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35094\ : std_logic;
signal \N__35091\ : std_logic;
signal \N__35088\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35085\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35071\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35042\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35036\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35027\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35021\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34986\ : std_logic;
signal \N__34983\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34977\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34961\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34946\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34942\ : std_logic;
signal \N__34939\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34933\ : std_logic;
signal \N__34926\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34916\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34899\ : std_logic;
signal \N__34896\ : std_logic;
signal \N__34893\ : std_logic;
signal \N__34888\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34849\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34839\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34836\ : std_logic;
signal \N__34833\ : std_logic;
signal \N__34828\ : std_logic;
signal \N__34825\ : std_logic;
signal \N__34822\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34814\ : std_logic;
signal \N__34813\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34807\ : std_logic;
signal \N__34804\ : std_logic;
signal \N__34801\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34778\ : std_logic;
signal \N__34777\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34759\ : std_logic;
signal \N__34756\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34727\ : std_logic;
signal \N__34726\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34668\ : std_logic;
signal \N__34665\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34653\ : std_logic;
signal \N__34650\ : std_logic;
signal \N__34647\ : std_logic;
signal \N__34644\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34623\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34614\ : std_logic;
signal \N__34611\ : std_logic;
signal \N__34608\ : std_logic;
signal \N__34605\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34596\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34587\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34554\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34548\ : std_logic;
signal \N__34545\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34539\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34509\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34447\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34439\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34431\ : std_logic;
signal \N__34430\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34424\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34415\ : std_logic;
signal \N__34412\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34401\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34395\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34377\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34342\ : std_logic;
signal \N__34339\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34329\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34323\ : std_logic;
signal \N__34320\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34284\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34278\ : std_logic;
signal \N__34275\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34251\ : std_logic;
signal \N__34250\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34243\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34223\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34212\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34208\ : std_logic;
signal \N__34203\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34188\ : std_logic;
signal \N__34185\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34179\ : std_logic;
signal \N__34176\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34161\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34135\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34127\ : std_logic;
signal \N__34124\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34104\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34098\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34082\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34044\ : std_logic;
signal \N__34041\ : std_logic;
signal \N__34038\ : std_logic;
signal \N__34035\ : std_logic;
signal \N__34032\ : std_logic;
signal \N__34029\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33996\ : std_logic;
signal \N__33993\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33981\ : std_logic;
signal \N__33978\ : std_logic;
signal \N__33975\ : std_logic;
signal \N__33972\ : std_logic;
signal \N__33969\ : std_logic;
signal \N__33966\ : std_logic;
signal \N__33963\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33912\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33906\ : std_logic;
signal \N__33903\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33897\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33876\ : std_logic;
signal \N__33875\ : std_logic;
signal \N__33872\ : std_logic;
signal \N__33869\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33856\ : std_logic;
signal \N__33853\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33845\ : std_logic;
signal \N__33840\ : std_logic;
signal \N__33837\ : std_logic;
signal \N__33834\ : std_logic;
signal \N__33833\ : std_logic;
signal \N__33830\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33828\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33806\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33778\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33768\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33759\ : std_logic;
signal \N__33756\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33749\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33708\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33699\ : std_logic;
signal \N__33698\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33695\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33692\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33689\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33686\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33680\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33671\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33668\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33643\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33628\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33543\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33516\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33507\ : std_logic;
signal \N__33504\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33484\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33474\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33451\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33423\ : std_logic;
signal \N__33420\ : std_logic;
signal \N__33417\ : std_logic;
signal \N__33414\ : std_logic;
signal \N__33411\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33357\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33347\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33341\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33338\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33335\ : std_logic;
signal \N__33334\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33332\ : std_logic;
signal \N__33331\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33293\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33263\ : std_logic;
signal \N__33260\ : std_logic;
signal \N__33257\ : std_logic;
signal \N__33254\ : std_logic;
signal \N__33251\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33239\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33155\ : std_logic;
signal \N__33152\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33143\ : std_logic;
signal \N__33140\ : std_logic;
signal \N__33137\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33119\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33107\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33068\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33026\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33013\ : std_logic;
signal \N__33008\ : std_logic;
signal \N__33005\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32998\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32981\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32966\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32947\ : std_logic;
signal \N__32940\ : std_logic;
signal \N__32937\ : std_logic;
signal \N__32934\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32911\ : std_logic;
signal \N__32906\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32888\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32854\ : std_logic;
signal \N__32851\ : std_logic;
signal \N__32848\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32828\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32808\ : std_logic;
signal \N__32805\ : std_logic;
signal \N__32802\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32798\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32785\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32772\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32738\ : std_logic;
signal \N__32737\ : std_logic;
signal \N__32734\ : std_logic;
signal \N__32729\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32691\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32684\ : std_logic;
signal \N__32683\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32677\ : std_logic;
signal \N__32674\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32663\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32639\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32615\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32605\ : std_logic;
signal \N__32604\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32579\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32572\ : std_logic;
signal \N__32569\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32559\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32555\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32545\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32534\ : std_logic;
signal \N__32533\ : std_logic;
signal \N__32528\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32487\ : std_logic;
signal \N__32486\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32461\ : std_logic;
signal \N__32458\ : std_logic;
signal \N__32453\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32387\ : std_logic;
signal \N__32384\ : std_logic;
signal \N__32381\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32358\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32346\ : std_logic;
signal \N__32343\ : std_logic;
signal \N__32340\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32334\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32325\ : std_logic;
signal \N__32322\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32295\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32283\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32274\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32256\ : std_logic;
signal \N__32253\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32220\ : std_logic;
signal \N__32217\ : std_logic;
signal \N__32214\ : std_logic;
signal \N__32211\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32205\ : std_logic;
signal \N__32202\ : std_logic;
signal \N__32199\ : std_logic;
signal \N__32196\ : std_logic;
signal \N__32193\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32175\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32166\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32154\ : std_logic;
signal \N__32151\ : std_logic;
signal \N__32148\ : std_logic;
signal \N__32145\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32121\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32115\ : std_logic;
signal \N__32112\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32106\ : std_logic;
signal \N__32103\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32037\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32005\ : std_logic;
signal \N__32002\ : std_logic;
signal \N__31997\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31984\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31958\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31946\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31930\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31919\ : std_logic;
signal \N__31918\ : std_logic;
signal \N__31915\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31886\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31877\ : std_logic;
signal \N__31874\ : std_logic;
signal \N__31871\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31862\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31856\ : std_logic;
signal \N__31853\ : std_logic;
signal \N__31850\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31841\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31835\ : std_logic;
signal \N__31832\ : std_logic;
signal \N__31829\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31817\ : std_logic;
signal \N__31816\ : std_logic;
signal \N__31811\ : std_logic;
signal \N__31808\ : std_logic;
signal \N__31805\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31796\ : std_logic;
signal \N__31793\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31784\ : std_logic;
signal \N__31781\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31772\ : std_logic;
signal \N__31771\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31718\ : std_logic;
signal \N__31715\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31709\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31670\ : std_logic;
signal \N__31667\ : std_logic;
signal \N__31664\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31655\ : std_logic;
signal \N__31652\ : std_logic;
signal \N__31649\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31640\ : std_logic;
signal \N__31637\ : std_logic;
signal \N__31634\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31625\ : std_logic;
signal \N__31622\ : std_logic;
signal \N__31619\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31610\ : std_logic;
signal \N__31607\ : std_logic;
signal \N__31604\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31592\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31577\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31571\ : std_logic;
signal \N__31568\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31559\ : std_logic;
signal \N__31556\ : std_logic;
signal \N__31553\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31535\ : std_logic;
signal \N__31532\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31505\ : std_logic;
signal \N__31502\ : std_logic;
signal \N__31499\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31490\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31484\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31476\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31469\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31454\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31424\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31415\ : std_logic;
signal \N__31414\ : std_logic;
signal \N__31411\ : std_logic;
signal \N__31408\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31402\ : std_logic;
signal \N__31397\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31391\ : std_logic;
signal \N__31388\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31380\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31307\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31300\ : std_logic;
signal \N__31297\ : std_logic;
signal \N__31294\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31272\ : std_logic;
signal \N__31269\ : std_logic;
signal \N__31266\ : std_logic;
signal \N__31265\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31254\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31250\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31245\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31238\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31236\ : std_logic;
signal \N__31235\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31233\ : std_logic;
signal \N__31232\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31230\ : std_logic;
signal \N__31229\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31223\ : std_logic;
signal \N__31220\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31217\ : std_logic;
signal \N__31216\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31213\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31211\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31205\ : std_logic;
signal \N__31202\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31199\ : std_logic;
signal \N__31196\ : std_logic;
signal \N__31193\ : std_logic;
signal \N__31190\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31178\ : std_logic;
signal \N__31169\ : std_logic;
signal \N__31166\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31142\ : std_logic;
signal \N__31133\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31122\ : std_logic;
signal \N__31121\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31118\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31106\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31100\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31058\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31031\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31004\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30997\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30988\ : std_logic;
signal \N__30985\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30971\ : std_logic;
signal \N__30970\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30964\ : std_logic;
signal \N__30961\ : std_logic;
signal \N__30960\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30938\ : std_logic;
signal \N__30935\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30916\ : std_logic;
signal \N__30913\ : std_logic;
signal \N__30910\ : std_logic;
signal \N__30907\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30901\ : std_logic;
signal \N__30894\ : std_logic;
signal \N__30893\ : std_logic;
signal \N__30890\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30876\ : std_logic;
signal \N__30873\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30858\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30836\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30824\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30782\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30773\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30766\ : std_logic;
signal \N__30763\ : std_logic;
signal \N__30760\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30733\ : std_logic;
signal \N__30730\ : std_logic;
signal \N__30727\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30650\ : std_logic;
signal \N__30647\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30632\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30622\ : std_logic;
signal \N__30619\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30611\ : std_logic;
signal \N__30606\ : std_logic;
signal \N__30605\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30582\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30566\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30540\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30486\ : std_logic;
signal \N__30483\ : std_logic;
signal \N__30480\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30468\ : std_logic;
signal \N__30465\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30456\ : std_logic;
signal \N__30453\ : std_logic;
signal \N__30450\ : std_logic;
signal \N__30447\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30432\ : std_logic;
signal \N__30429\ : std_logic;
signal \N__30426\ : std_logic;
signal \N__30423\ : std_logic;
signal \N__30420\ : std_logic;
signal \N__30417\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30399\ : std_logic;
signal \N__30396\ : std_logic;
signal \N__30393\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30369\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30339\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30321\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30309\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30298\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30279\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30272\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30268\ : std_logic;
signal \N__30265\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30253\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30241\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30227\ : std_logic;
signal \N__30224\ : std_logic;
signal \N__30223\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30184\ : std_logic;
signal \N__30181\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30161\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30155\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30126\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30097\ : std_logic;
signal \N__30094\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30080\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30076\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30048\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30039\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30024\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29964\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29948\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29939\ : std_logic;
signal \N__29938\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29922\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29917\ : std_logic;
signal \N__29914\ : std_logic;
signal \N__29911\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29901\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29861\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29844\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29834\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29786\ : std_logic;
signal \N__29785\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29779\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29762\ : std_logic;
signal \N__29759\ : std_logic;
signal \N__29758\ : std_logic;
signal \N__29755\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29711\ : std_logic;
signal \N__29708\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29688\ : std_logic;
signal \N__29685\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29679\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29669\ : std_logic;
signal \N__29666\ : std_logic;
signal \N__29663\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29654\ : std_logic;
signal \N__29651\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29645\ : std_logic;
signal \N__29642\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29624\ : std_logic;
signal \N__29621\ : std_logic;
signal \N__29618\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29585\ : std_logic;
signal \N__29582\ : std_logic;
signal \N__29579\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29564\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29558\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29531\ : std_logic;
signal \N__29528\ : std_logic;
signal \N__29525\ : std_logic;
signal \N__29522\ : std_logic;
signal \N__29519\ : std_logic;
signal \N__29516\ : std_logic;
signal \N__29513\ : std_logic;
signal \N__29510\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29492\ : std_logic;
signal \N__29489\ : std_logic;
signal \N__29486\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29468\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29462\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29456\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29444\ : std_logic;
signal \N__29441\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29435\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29429\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29411\ : std_logic;
signal \N__29408\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29375\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29361\ : std_logic;
signal \N__29358\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29351\ : std_logic;
signal \N__29348\ : std_logic;
signal \N__29345\ : std_logic;
signal \N__29342\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29312\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29303\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29291\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29264\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29243\ : std_logic;
signal \N__29240\ : std_logic;
signal \N__29237\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29231\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29213\ : std_logic;
signal \N__29210\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29193\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29150\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29120\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29082\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29073\ : std_logic;
signal \N__29072\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29063\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29040\ : std_logic;
signal \N__29039\ : std_logic;
signal \N__29036\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29018\ : std_logic;
signal \N__29013\ : std_logic;
signal \N__29010\ : std_logic;
signal \N__29009\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28997\ : std_logic;
signal \N__28994\ : std_logic;
signal \N__28991\ : std_logic;
signal \N__28988\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28970\ : std_logic;
signal \N__28967\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28936\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28906\ : std_logic;
signal \N__28903\ : std_logic;
signal \N__28900\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28894\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28878\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28842\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28840\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28828\ : std_logic;
signal \N__28825\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28811\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28792\ : std_logic;
signal \N__28789\ : std_logic;
signal \N__28786\ : std_logic;
signal \N__28783\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28768\ : std_logic;
signal \N__28765\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28745\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28730\ : std_logic;
signal \N__28727\ : std_logic;
signal \N__28724\ : std_logic;
signal \N__28721\ : std_logic;
signal \N__28718\ : std_logic;
signal \N__28715\ : std_logic;
signal \N__28712\ : std_logic;
signal \N__28709\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28703\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28688\ : std_logic;
signal \N__28685\ : std_logic;
signal \N__28682\ : std_logic;
signal \N__28679\ : std_logic;
signal \N__28676\ : std_logic;
signal \N__28673\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28652\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28610\ : std_logic;
signal \N__28609\ : std_logic;
signal \N__28606\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28571\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28558\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28549\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28541\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28528\ : std_logic;
signal \N__28525\ : std_logic;
signal \N__28520\ : std_logic;
signal \N__28517\ : std_logic;
signal \N__28514\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28508\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28504\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28495\ : std_logic;
signal \N__28492\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28478\ : std_logic;
signal \N__28477\ : std_logic;
signal \N__28474\ : std_logic;
signal \N__28471\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28445\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28430\ : std_logic;
signal \N__28427\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28402\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28393\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28387\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28381\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28343\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28339\ : std_logic;
signal \N__28336\ : std_logic;
signal \N__28333\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28323\ : std_logic;
signal \N__28320\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28280\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28265\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28259\ : std_logic;
signal \N__28256\ : std_logic;
signal \N__28253\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28244\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28235\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28220\ : std_logic;
signal \N__28217\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28210\ : std_logic;
signal \N__28207\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28193\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28173\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28167\ : std_logic;
signal \N__28164\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28145\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28133\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28103\ : std_logic;
signal \N__28102\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28075\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28066\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28048\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28016\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__28001\ : std_logic;
signal \N__28000\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27982\ : std_logic;
signal \N__27979\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27961\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27947\ : std_logic;
signal \N__27946\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27938\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27929\ : std_logic;
signal \N__27926\ : std_logic;
signal \N__27923\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27893\ : std_logic;
signal \N__27890\ : std_logic;
signal \N__27887\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27879\ : std_logic;
signal \N__27876\ : std_logic;
signal \N__27875\ : std_logic;
signal \N__27872\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27833\ : std_logic;
signal \N__27830\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27815\ : std_logic;
signal \N__27812\ : std_logic;
signal \N__27809\ : std_logic;
signal \N__27806\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27761\ : std_logic;
signal \N__27758\ : std_logic;
signal \N__27755\ : std_logic;
signal \N__27752\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27744\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27734\ : std_logic;
signal \N__27729\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27725\ : std_logic;
signal \N__27722\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27716\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27693\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27689\ : std_logic;
signal \N__27686\ : std_logic;
signal \N__27683\ : std_logic;
signal \N__27680\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27668\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27651\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27644\ : std_logic;
signal \N__27641\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27633\ : std_logic;
signal \N__27630\ : std_logic;
signal \N__27629\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27604\ : std_logic;
signal \N__27601\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27586\ : std_logic;
signal \N__27583\ : std_logic;
signal \N__27580\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27521\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27511\ : std_logic;
signal \N__27508\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27500\ : std_logic;
signal \N__27499\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27476\ : std_logic;
signal \N__27475\ : std_logic;
signal \N__27472\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27463\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27449\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27425\ : std_logic;
signal \N__27424\ : std_logic;
signal \N__27421\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27404\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27392\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27225\ : std_logic;
signal \N__27222\ : std_logic;
signal \N__27219\ : std_logic;
signal \N__27216\ : std_logic;
signal \N__27213\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27201\ : std_logic;
signal \N__27198\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27192\ : std_logic;
signal \N__27189\ : std_logic;
signal \N__27186\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27180\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27173\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27158\ : std_logic;
signal \N__27153\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27104\ : std_logic;
signal \N__27101\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27093\ : std_logic;
signal \N__27090\ : std_logic;
signal \N__27089\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27085\ : std_logic;
signal \N__27082\ : std_logic;
signal \N__27079\ : std_logic;
signal \N__27074\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27062\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27059\ : std_logic;
signal \N__27056\ : std_logic;
signal \N__27053\ : std_logic;
signal \N__27050\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27029\ : std_logic;
signal \N__27026\ : std_logic;
signal \N__27023\ : std_logic;
signal \N__27020\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27005\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27002\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26980\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26963\ : std_logic;
signal \N__26960\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26952\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26922\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26918\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26913\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26908\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26900\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26800\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26794\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26774\ : std_logic;
signal \N__26771\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26750\ : std_logic;
signal \N__26747\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26741\ : std_logic;
signal \N__26740\ : std_logic;
signal \N__26737\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26708\ : std_logic;
signal \N__26705\ : std_logic;
signal \N__26702\ : std_logic;
signal \N__26699\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26678\ : std_logic;
signal \N__26677\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26661\ : std_logic;
signal \N__26654\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26605\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26588\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26584\ : std_logic;
signal \N__26579\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26575\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26546\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26540\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26534\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26526\ : std_logic;
signal \N__26523\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26507\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26462\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26439\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26433\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26429\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26386\ : std_logic;
signal \N__26383\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26368\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26318\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26306\ : std_logic;
signal \N__26303\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26291\ : std_logic;
signal \N__26290\ : std_logic;
signal \N__26287\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26244\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26240\ : std_logic;
signal \N__26237\ : std_logic;
signal \N__26234\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26225\ : std_logic;
signal \N__26222\ : std_logic;
signal \N__26219\ : std_logic;
signal \N__26214\ : std_logic;
signal \N__26211\ : std_logic;
signal \N__26210\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26109\ : std_logic;
signal \N__26106\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26065\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26055\ : std_logic;
signal \N__26052\ : std_logic;
signal \N__26049\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26045\ : std_logic;
signal \N__26042\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26033\ : std_logic;
signal \N__26030\ : std_logic;
signal \N__26025\ : std_logic;
signal \N__26022\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26018\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26014\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25994\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25980\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25956\ : std_logic;
signal \N__25953\ : std_logic;
signal \N__25950\ : std_logic;
signal \N__25947\ : std_logic;
signal \N__25944\ : std_logic;
signal \N__25941\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25928\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25916\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25794\ : std_logic;
signal \N__25791\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25764\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25757\ : std_logic;
signal \N__25754\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25739\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25731\ : std_logic;
signal \N__25728\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25692\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25679\ : std_logic;
signal \N__25676\ : std_logic;
signal \N__25671\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25625\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25610\ : std_logic;
signal \N__25607\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25596\ : std_logic;
signal \N__25593\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25551\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25476\ : std_logic;
signal \N__25473\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25452\ : std_logic;
signal \N__25449\ : std_logic;
signal \N__25446\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25383\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25368\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25323\ : std_logic;
signal \N__25320\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25308\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25242\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25233\ : std_logic;
signal \N__25230\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25161\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25141\ : std_logic;
signal \N__25138\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25120\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25114\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25111\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25107\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25098\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25095\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25034\ : std_logic;
signal \N__25025\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24987\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24981\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24951\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24945\ : std_logic;
signal \N__24942\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24863\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24835\ : std_logic;
signal \N__24832\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24810\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24721\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24706\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24576\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24561\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24531\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24519\ : std_logic;
signal \N__24516\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24444\ : std_logic;
signal \N__24441\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24423\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24390\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24366\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24267\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24207\ : std_logic;
signal \N__24204\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24171\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23970\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23936\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23916\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23897\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23817\ : std_logic;
signal \N__23814\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23796\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23765\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23702\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23679\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23619\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23594\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23585\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23556\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23549\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23526\ : std_logic;
signal \N__23525\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23491\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23445\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23427\ : std_logic;
signal \N__23426\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23423\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23243\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23240\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23237\ : std_logic;
signal \N__23234\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23207\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23114\ : std_logic;
signal \N__23111\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23076\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22881\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22757\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22722\ : std_logic;
signal \N__22719\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22448\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22241\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22170\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22136\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22029\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22023\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21909\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21789\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21627\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21618\ : std_logic;
signal \N__21615\ : std_logic;
signal \N__21612\ : std_logic;
signal \N__21609\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21492\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21396\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21136\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21058\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20902\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20841\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20826\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20769\ : std_logic;
signal \N__20766\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20751\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20715\ : std_logic;
signal \N__20712\ : std_logic;
signal \N__20709\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20700\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20613\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20585\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20543\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20448\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20315\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20121\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19970\ : std_logic;
signal \N__19967\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19773\ : std_logic;
signal \N__19770\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19764\ : std_logic;
signal \N__19761\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19581\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19482\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19476\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19395\ : std_logic;
signal \N__19392\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19241\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19235\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19107\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18999\ : std_logic;
signal delay_tr_input_ibuf_gb_io_gb_input : std_logic;
signal delay_hc_input_ibuf_gb_io_gb_input : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_9\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_17\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_25\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\ : std_logic;
signal un7_start_stop : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.un1_integrator\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_44\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_77\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_43_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_91\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_98_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_158\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_96_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_160\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_94\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_97\ : std_logic;
signal pwm_duty_input_1 : std_logic;
signal pwm_duty_input_2 : std_logic;
signal pwm_duty_input_0 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_1Z0Z_0\ : std_logic;
signal \pwm_generator_inst.N_7_cascade_\ : std_logic;
signal pwm_duty_input_9 : std_logic;
signal pwm_duty_input_6 : std_logic;
signal pwm_duty_input_7 : std_logic;
signal pwm_duty_input_8 : std_logic;
signal pwm_duty_input_3 : std_logic;
signal pwm_duty_input_4 : std_logic;
signal \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\ : std_logic;
signal pwm_duty_input_5 : std_logic;
signal \pwm_generator_inst.O_0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_0\ : std_logic;
signal \bfn_2_24_0_\ : std_logic;
signal \pwm_generator_inst.O_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_1\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_0\ : std_logic;
signal \pwm_generator_inst.O_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_1\ : std_logic;
signal \pwm_generator_inst.O_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_3\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_2\ : std_logic;
signal \pwm_generator_inst.O_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_3\ : std_logic;
signal \pwm_generator_inst.O_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_4\ : std_logic;
signal \pwm_generator_inst.O_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_5\ : std_logic;
signal \pwm_generator_inst.O_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_7\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_7\ : std_logic;
signal \pwm_generator_inst.O_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_8\ : std_logic;
signal \bfn_2_25_0_\ : std_logic;
signal \pwm_generator_inst.O_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15\ : std_logic;
signal \bfn_2_26_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18\ : std_logic;
signal \N_88_i_i\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_1\ : std_logic;
signal \bfn_3_17_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto3\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.un7_enablelto4\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_9\ : std_logic;
signal \bfn_3_18_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\ : std_logic;
signal \bfn_3_19_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\ : std_logic;
signal \bfn_3_20_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\ : std_logic;
signal \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_27\ : std_logic;
signal \bfn_3_24_0_\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7\ : std_logic;
signal \bfn_3_25_0_\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_16\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_6\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_15\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_5\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_18\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_8\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_17\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_47\ : std_logic;
signal \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.N_46\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.integratorZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_26\ : std_logic;
signal \pwm_generator_inst.un3_threshold\ : std_logic;
signal \bfn_4_22_0_\ : std_logic;
signal \pwm_generator_inst.O_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0\ : std_logic;
signal \pwm_generator_inst.O_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1\ : std_logic;
signal \pwm_generator_inst.O_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_3\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_4\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_5\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\ : std_logic;
signal \bfn_4_23_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15\ : std_logic;
signal \bfn_4_24_0_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_2\ : std_logic;
signal \pwm_generator_inst.O_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_10\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_0\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_14\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_4\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\ : std_logic;
signal \pwm_generator_inst.un19_threshold_axb_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_30\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_axbZ0Z_4\ : std_logic;
signal \bfn_5_23_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_17\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_18\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_2\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_19\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_3\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_20\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_4\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_21\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_6\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_5\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_22\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_7\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_6\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_7\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_23\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_8\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\ : std_logic;
signal \bfn_5_24_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_1_24\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_9\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_8\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_10\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_9\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_11\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_10\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_12\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_11\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_12\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_14\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_13\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_14\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15\ : std_logic;
signal \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\ : std_logic;
signal \bfn_5_25_0_\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\ : std_logic;
signal \elapsed_time_ns_1_RNI2COBB_0_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIJI91B_0_7\ : std_logic;
signal \elapsed_time_ns_1_RNIU7OBB_0_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_7\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_15\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_23\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_166_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.running_i\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.runningZ0\ : std_logic;
signal \delay_measurement_inst.stop_timer_trZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_trZ0\ : std_logic;
signal delay_tr_input_c_g : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\ : std_logic;
signal \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\ : std_logic;
signal \bfn_7_26_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_0\ : std_logic;
signal \pwm_generator_inst.counter_cry_1\ : std_logic;
signal \pwm_generator_inst.counter_cry_2\ : std_logic;
signal \pwm_generator_inst.counter_cry_3\ : std_logic;
signal \pwm_generator_inst.counter_cry_4\ : std_logic;
signal \pwm_generator_inst.counter_cry_5\ : std_logic;
signal \pwm_generator_inst.counter_cry_6\ : std_logic;
signal \pwm_generator_inst.counter_cry_7\ : std_logic;
signal \bfn_7_27_0_\ : std_logic;
signal \pwm_generator_inst.counter_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt18\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22\ : std_logic;
signal \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt24\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25\ : std_logic;
signal \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNI1CPBB_0_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\ : std_logic;
signal \bfn_8_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.N_165_i\ : std_logic;
signal \pwm_generator_inst.N_16\ : std_logic;
signal \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\ : std_logic;
signal \pwm_generator_inst.N_17\ : std_logic;
signal \pwm_generator_inst.threshold_0\ : std_logic;
signal \pwm_generator_inst.counter_i_0\ : std_logic;
signal \bfn_8_24_0_\ : std_logic;
signal \pwm_generator_inst.threshold_1\ : std_logic;
signal \pwm_generator_inst.counter_i_1\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_0\ : std_logic;
signal \pwm_generator_inst.threshold_2\ : std_logic;
signal \pwm_generator_inst.counter_i_2\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_1\ : std_logic;
signal \pwm_generator_inst.threshold_3\ : std_logic;
signal \pwm_generator_inst.counter_i_3\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_2\ : std_logic;
signal \pwm_generator_inst.threshold_4\ : std_logic;
signal \pwm_generator_inst.counter_i_4\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_3\ : std_logic;
signal \pwm_generator_inst.threshold_5\ : std_logic;
signal \pwm_generator_inst.counter_i_5\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_4\ : std_logic;
signal \pwm_generator_inst.threshold_6\ : std_logic;
signal \pwm_generator_inst.counter_i_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_5\ : std_logic;
signal \pwm_generator_inst.threshold_7\ : std_logic;
signal \pwm_generator_inst.counter_i_7\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_6\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_7\ : std_logic;
signal \pwm_generator_inst.threshold_8\ : std_logic;
signal \pwm_generator_inst.counter_i_8\ : std_logic;
signal \bfn_8_25_0_\ : std_logic;
signal \pwm_generator_inst.threshold_9\ : std_logic;
signal \pwm_generator_inst.counter_i_9\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_8\ : std_logic;
signal \pwm_generator_inst.un14_counter_cry_9\ : std_logic;
signal pwm_output_c : std_logic;
signal \pwm_generator_inst.counterZ0Z_8\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_9\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_7\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_0\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_4\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_1\ : std_logic;
signal \pwm_generator_inst.un1_counterlto2_0_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_3\ : std_logic;
signal \pwm_generator_inst.un1_counterlto9_2\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_6\ : std_logic;
signal \pwm_generator_inst.un1_counterlt9_cascade_\ : std_logic;
signal \pwm_generator_inst.counterZ0Z_5\ : std_logic;
signal \pwm_generator_inst.un1_counter_0\ : std_logic;
signal clk_12mhz : std_logic;
signal \GB_BUFFER_clk_12mhz_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI2DPBB_0_24\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNIV8OBB_0_12\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\ : std_logic;
signal \elapsed_time_ns_1_RNIED91B_0_2\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\ : std_logic;
signal \elapsed_time_ns_1_RNIIH91B_0_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\ : std_logic;
signal \elapsed_time_ns_1_RNIGF91B_0_4\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\ : std_logic;
signal \elapsed_time_ns_1_RNI0CQBB_0_31\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\ : std_logic;
signal \elapsed_time_ns_1_RNI5GPBB_0_27\ : std_logic;
signal \elapsed_time_ns_1_RNIV9PBB_0_21\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNI6GOBB_0_19\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axb_0\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_6\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_8\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_14\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_16\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_22\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_24\ : std_logic;
signal \bfn_9_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_28\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_cry_30\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_termZ0Z_31\ : std_logic;
signal \current_shift_inst.PI_CTRL.un8_enablelto31\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \elapsed_time_ns_1_RNI0AOBB_0_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\ : std_logic;
signal \elapsed_time_ns_1_RNIHG91B_0_5\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\ : std_logic;
signal \elapsed_time_ns_1_RNILK91B_0_9\ : std_logic;
signal \elapsed_time_ns_1_RNIT6OBB_0_10\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_1\ : std_logic;
signal \bfn_10_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_9\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_16\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\ : std_logic;
signal \elapsed_time_ns_1_RNI4FPBB_0_26\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt30\ : std_logic;
signal \elapsed_time_ns_1_RNIVAQBB_0_30\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.prop_term_1_0\ : std_logic;
signal \elapsed_time_ns_1_RNI7IPBB_0_29\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_16\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_tr.runningZ0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\ : std_logic;
signal \elapsed_time_ns_1_RNIFE91B_0_3\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\ : std_logic;
signal \elapsed_time_ns_1_RNI5FOBB_0_18\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\ : std_logic;
signal \elapsed_time_ns_1_RNIKJ91B_0_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\ : std_logic;
signal \elapsed_time_ns_1_RNI1BOBB_0_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\ : std_logic;
signal \current_shift_inst.N_1263_i\ : std_logic;
signal \current_shift_inst.control_input_1\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\ : std_logic;
signal \current_shift_inst.control_input_cry_0\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\ : std_logic;
signal \current_shift_inst.control_input_cry_1\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\ : std_logic;
signal \current_shift_inst.control_input_cry_2\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\ : std_logic;
signal \current_shift_inst.control_input_cry_3\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\ : std_logic;
signal \current_shift_inst.control_input_cry_4\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\ : std_logic;
signal \current_shift_inst.control_input_cry_5\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\ : std_logic;
signal \current_shift_inst.control_input_cry_6\ : std_logic;
signal \current_shift_inst.control_input_cry_7\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\ : std_logic;
signal \current_shift_inst.control_input_cry_8\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\ : std_logic;
signal \current_shift_inst.control_input_cry_9\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\ : std_logic;
signal \current_shift_inst.control_input_cry_10\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\ : std_logic;
signal \current_shift_inst.control_input_cry_11\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\ : std_logic;
signal \current_shift_inst.control_input_cry_12\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\ : std_logic;
signal \current_shift_inst.control_input_cry_13\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\ : std_logic;
signal \current_shift_inst.control_input_cry_14\ : std_logic;
signal \current_shift_inst.control_input_cry_15\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\ : std_logic;
signal \current_shift_inst.control_input_cry_16\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\ : std_logic;
signal \current_shift_inst.control_input_cry_17\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\ : std_logic;
signal \current_shift_inst.control_input_cry_18\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\ : std_logic;
signal \current_shift_inst.control_input_cry_19\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\ : std_logic;
signal \current_shift_inst.control_input_cry_20\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\ : std_logic;
signal \current_shift_inst.control_input_cry_21\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\ : std_logic;
signal \current_shift_inst.control_input_cry_22\ : std_logic;
signal \current_shift_inst.control_input_cry_23\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\ : std_logic;
signal \bfn_11_16_0_\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\ : std_logic;
signal \current_shift_inst.control_input_cry_24\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\ : std_logic;
signal \current_shift_inst.control_input_cry_25\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\ : std_logic;
signal \current_shift_inst.control_input_cry_26\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\ : std_logic;
signal \current_shift_inst.control_input_cry_27\ : std_logic;
signal \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\ : std_logic;
signal \current_shift_inst.control_input_cry_28\ : std_logic;
signal \current_shift_inst.control_input_cry_29\ : std_logic;
signal \current_shift_inst.control_input_31\ : std_logic;
signal \current_shift_inst.control_input_axb_26\ : std_logic;
signal \current_shift_inst.control_input_axb_29\ : std_logic;
signal \current_shift_inst.control_input_axb_17\ : std_logic;
signal s4_phy_c : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\ : std_logic;
signal \elapsed_time_ns_1_RNIDC91B_0_1\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst1.stoper_tr.start_latchedZ0\ : std_logic;
signal \elapsed_time_ns_1_RNI3DOBB_0_16\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\ : std_logic;
signal il_max_comp2_c : std_logic;
signal il_min_comp2_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst2.N_54_0\ : std_logic;
signal \phase_controller_inst2.tr_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\ : std_logic;
signal \elapsed_time_ns_1_RNI6HPBB_0_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un1_start_g\ : std_logic;
signal \current_shift_inst.control_input_axb_2\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un4_running_lt28\ : std_logic;
signal \current_shift_inst.control_input_axb_6\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU8PBB_0_20\ : std_logic;
signal \current_shift_inst.control_input_axb_9\ : std_logic;
signal \current_shift_inst.control_input_axb_12\ : std_logic;
signal \current_shift_inst.control_input_axb_13\ : std_logic;
signal \current_shift_inst.control_input_axb_11\ : std_logic;
signal \current_shift_inst.control_input_axb_15\ : std_logic;
signal \current_shift_inst.control_input_axb_14\ : std_logic;
signal \current_shift_inst.control_input_axb_16\ : std_logic;
signal \current_shift_inst.control_input_axb_18\ : std_logic;
signal \current_shift_inst.control_input_axb_19\ : std_logic;
signal \current_shift_inst.control_input_axb_20\ : std_logic;
signal \current_shift_inst.control_input_axb_10\ : std_logic;
signal \current_shift_inst.control_input_axb_23\ : std_logic;
signal \current_shift_inst.control_input_axb_24\ : std_logic;
signal \current_shift_inst.control_input_axb_25\ : std_logic;
signal \current_shift_inst.control_input_axb_27\ : std_logic;
signal delay_hc_input_c_g : std_logic;
signal s3_phy_c : std_logic;
signal \GB_BUFFER_red_c_g_THRU_CO\ : std_logic;
signal \phase_controller_inst1.state_ns_0_0_1\ : std_logic;
signal \phase_controller_inst1.tr_time_passed\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst1.start_flagZ0\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst1.N_54_0\ : std_logic;
signal \phase_controller_inst1.hc_time_passed\ : std_logic;
signal il_max_comp1_c : std_logic;
signal \phase_controller_inst2.state_ns_0_0_1\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stateZ0Z_2\ : std_logic;
signal \phase_controller_inst2.N_61\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_16\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28\ : std_logic;
signal \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI7ADN9_0_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV2EN9_0_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\ : std_logic;
signal \elapsed_time_ns_1_RNI04EN9_0_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s1\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_16\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s1\ : std_logic;
signal \bfn_13_19_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s1\ : std_logic;
signal s2_phy_c : std_logic;
signal state_3 : std_logic;
signal s1_phy_c : std_logic;
signal \current_shift_inst.start_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.stop_timer_sZ0Z1\ : std_logic;
signal \current_shift_inst.timer_s1.N_161_i\ : std_logic;
signal il_min_comp1_c : std_logic;
signal \phase_controller_inst1.N_61\ : std_logic;
signal \phase_controller_inst1.stateZ0Z_1\ : std_logic;
signal start_stop_c : std_logic;
signal \phase_controller_inst2.stateZ0Z_4\ : std_logic;
signal \phase_controller_inst2.start_flagZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\ : std_logic;
signal \phase_controller_inst2.stoper_tr.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.runningZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_trZ0\ : std_logic;
signal \phase_controller_inst2.stoper_tr.un2_start_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\ : std_logic;
signal \bfn_14_13_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_3_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_5\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_4_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_5_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_6_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_7_s0\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_9\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_8_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_9_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_10_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_12\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_11_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_13\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_12_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_14\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_13_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_15\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_14_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_15_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_16\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_16_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_18\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_17_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_19\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_18_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_19_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_21\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_20_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_22\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_21_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_23\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_22_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_23_s0\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_24_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_26\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_25_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_27\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_26_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_28\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_27_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_29\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_28_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_30\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_29_s0\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_31\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_30_s0\ : std_logic;
signal \current_shift_inst.control_input_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_19\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_25\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_25\ : std_logic;
signal \current_shift_inst.control_input_axb_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_24\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_24\ : std_logic;
signal \current_shift_inst.control_input_axb_21\ : std_logic;
signal \current_shift_inst.un38_control_input_5_0\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\ : std_logic;
signal \delay_measurement_inst.delay_tr_timer.delay_tr3\ : std_logic;
signal \elapsed_time_ns_1_RNI4EOBB_0_17\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_fast_31\ : std_logic;
signal \current_shift_inst.timer_s1.runningZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst1.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt16\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \elapsed_time_ns_1_RNIH33T9_0_5\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\ : std_logic;
signal \elapsed_time_ns_1_RNI68CN9_0_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\ : std_logic;
signal \elapsed_time_ns_1_RNIE03T9_0_2\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \elapsed_time_ns_1_RNIG23T9_0_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_4\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_4\ : std_logic;
signal \current_shift_inst.control_input_axb_1\ : std_logic;
signal \elapsed_time_ns_1_RNIK63T9_0_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_8\ : std_logic;
signal \current_shift_inst.control_input_axb_5\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_3\ : std_logic;
signal \current_shift_inst.control_input_axb_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_7\ : std_logic;
signal \current_shift_inst.control_input_axb_4\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_10\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_10\ : std_logic;
signal \current_shift_inst.control_input_axb_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_11\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_11\ : std_logic;
signal \current_shift_inst.control_input_axb_8\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s0_6\ : std_logic;
signal \current_shift_inst.un38_control_input_0_s1_6\ : std_logic;
signal \current_shift_inst.control_input_axb_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_31\ : std_logic;
signal \bfn_15_21_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7\ : std_logic;
signal \bfn_15_22_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15\ : std_logic;
signal \bfn_15_23_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23\ : std_logic;
signal \bfn_15_24_0_\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\ : std_logic;
signal \phase_controller_inst2.hc_time_passed\ : std_logic;
signal \phase_controller_inst2.stoper_hc.runningZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un2_start_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latchedZ0\ : std_logic;
signal \phase_controller_inst2.start_timer_hcZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_1\ : std_logic;
signal \bfn_16_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_9\ : std_logic;
signal \bfn_16_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_time_i_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt18\ : std_logic;
signal \bfn_16_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\ : std_logic;
signal \bfn_16_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_16_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_3\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\ : std_logic;
signal \bfn_16_20_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\ : std_logic;
signal \bfn_16_21_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\ : std_logic;
signal \bfn_16_22_0_\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_22\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_18\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\ : std_logic;
signal \elapsed_time_ns_1_RNI25DN9_0_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\ : std_logic;
signal \bfn_17_8_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\ : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\ : std_logic;
signal \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\ : std_logic;
signal \elapsed_time_ns_1_RNITUBN9_0_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\ : std_logic;
signal \elapsed_time_ns_1_RNIUVBN9_0_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\ : std_logic;
signal \elapsed_time_ns_1_RNI03DN9_0_22\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\ : std_logic;
signal \elapsed_time_ns_1_RNI47DN9_0_26\ : std_logic;
signal \elapsed_time_ns_1_RNI14DN9_0_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\ : std_logic;
signal \elapsed_time_ns_1_RNIF13T9_0_3\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_0_s0_sf\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\ : std_logic;
signal \elapsed_time_ns_1_RNIL73T9_0_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\ : std_logic;
signal \elapsed_time_ns_1_RNIV0CN9_0_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_5\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\ : std_logic;
signal \bfn_17_15_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_3\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_1\ : std_logic;
signal \current_shift_inst.un4_control_input1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_2\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_3\ : std_logic;
signal \current_shift_inst.un4_control_input1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_4\ : std_logic;
signal \current_shift_inst.un4_control_input1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_7\ : std_logic;
signal \current_shift_inst.un4_control_input1_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_6\ : std_logic;
signal \current_shift_inst.un4_control_input1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_8\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_9\ : std_logic;
signal \current_shift_inst.un4_control_input1_10\ : std_logic;
signal \bfn_17_16_0_\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_10\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_11\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_12\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_14\ : std_logic;
signal \current_shift_inst.un4_control_input1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_15\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_18\ : std_logic;
signal \bfn_17_17_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_17\ : std_logic;
signal \current_shift_inst.un4_control_input1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_18\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_22\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_21\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_23\ : std_logic;
signal \current_shift_inst.un4_control_input1_24\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_22\ : std_logic;
signal \current_shift_inst.un4_control_input1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_23\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_24\ : std_logic;
signal \bfn_17_18_0_\ : std_logic;
signal \current_shift_inst.un4_control_input1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_25\ : std_logic;
signal \current_shift_inst.un4_control_input1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_26\ : std_logic;
signal \current_shift_inst.un4_control_input1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_27\ : std_logic;
signal \current_shift_inst.un4_control_input1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_cry_28\ : std_logic;
signal \current_shift_inst.un4_control_input1_31\ : std_logic;
signal \current_shift_inst.un4_control_input1_31_THRU_CO\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_4\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_3\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_6\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_5\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_13\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_12\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_7\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_6\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_9\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_8\ : std_logic;
signal \current_shift_inst.un4_control_input1_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNISV131_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_20\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_17\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_16\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_26\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_25\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_19\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_18\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_16\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_15\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_25\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_24\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_29\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_28\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_26\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_28\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_27\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_20\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_30\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_29\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_15\ : std_logic;
signal \current_shift_inst.un4_control_input1_15\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_12\ : std_logic;
signal \current_shift_inst.un4_control_input1_12\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\ : std_logic;
signal \bfn_17_23_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_0\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_2\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_3\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_2\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_4\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_3\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_5\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_4\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_5\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_7\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_6\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_7\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_8\ : std_logic;
signal \bfn_17_24_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_9\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_8\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_10\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_9\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_11\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_10\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_12\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_11\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_13\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_12\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_13\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_15\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_14\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_15\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_16\ : std_logic;
signal \bfn_17_25_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_17\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_16\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_18\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_17\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_19\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_18\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_20\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_19\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_21\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_20\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_21\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_23\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_22\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_23\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_24\ : std_logic;
signal \bfn_17_26_0_\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_25\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_24\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_26\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_25\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_27\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_26\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_28\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_27\ : std_logic;
signal \current_shift_inst.timer_s1.running_i\ : std_logic;
signal \current_shift_inst.timer_s1.counter_cry_28\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.timer_s1.N_162_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\ : std_logic;
signal \elapsed_time_ns_1_RNIU0DN9_0_20\ : std_logic;
signal \elapsed_time_ns_1_RNI46CN9_0_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\ : std_logic;
signal \elapsed_time_ns_1_RNI13CN9_0_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\ : std_logic;
signal \elapsed_time_ns_1_RNI35CN9_0_16\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\ : std_logic;
signal \elapsed_time_ns_1_RNI02CN9_0_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\ : std_logic;
signal \elapsed_time_ns_1_RNI24CN9_0_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\ : std_logic;
signal \elapsed_time_ns_1_RNIDV2T9_0_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\ : std_logic;
signal \elapsed_time_ns_1_RNI36DN9_0_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt26\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_lt20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\ : std_logic;
signal \elapsed_time_ns_1_RNIV1DN9_0_21\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\ : std_logic;
signal \elapsed_time_ns_1_RNII43T9_0_6\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\ : std_logic;
signal \elapsed_time_ns_1_RNIJ53T9_0_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\ : std_logic;
signal \bfn_18_11_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_2\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_3\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_4\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_5\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_6\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_7\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_8\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_9\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_10\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_11\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_12\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_13\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_15\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_16\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_17\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_18\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_19\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_20\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_21\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_22\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_23\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_24\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_25\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_26\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counter_cry_28\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\ : std_logic;
signal \current_shift_inst.un38_control_input_axb_31_s0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\ : std_logic;
signal \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_1\ : std_logic;
signal \current_shift_inst.timer_s1.counterZ0Z_1\ : std_logic;
signal \current_shift_inst.timer_s1.N_161_i_g\ : std_logic;
signal \current_shift_inst.un4_control_input_1_axb_1\ : std_logic;
signal \current_shift_inst.un38_control_input_5_1\ : std_logic;
signal \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31_rep1\ : std_logic;
signal \current_shift_inst.un4_control_input1_2\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_2\ : std_logic;
signal \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_13\ : std_logic;
signal \current_shift_inst.un4_control_input1_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_11\ : std_logic;
signal \current_shift_inst.un4_control_input1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_21\ : std_logic;
signal \current_shift_inst.un4_control_input1_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_31\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_s1_14\ : std_logic;
signal \current_shift_inst.un38_control_input_5_2\ : std_logic;
signal \current_shift_inst.un4_control_input1_14\ : std_logic;
signal \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\ : std_logic;
signal \elapsed_time_ns_1_RNI57CN9_0_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\ : std_logic;
signal \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\ : std_logic;
signal \phase_controller_inst2.stoper_hc.un1_start_g\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.delay_hc3\ : std_logic;
signal \elapsed_time_ns_1_RNI58DN9_0_27\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_164_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.N_163_i\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.running_i\ : std_logic;
signal \delay_measurement_inst.stop_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.start_timer_hcZ0\ : std_logic;
signal \delay_measurement_inst.delay_hc_timer.runningZ0\ : std_logic;
signal clk_100mhz_0 : std_logic;
signal red_c_g : std_logic;
signal \pwm_generator_inst.un2_threshold_1_25\ : std_logic;
signal \pwm_generator_inst.un2_threshold_2_1_15\ : std_logic;
signal \N_19_1\ : std_logic;
signal \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal reset_wire : std_logic;
signal start_stop_wire : std_logic;
signal il_max_comp2_wire : std_logic;
signal pwm_output_wire : std_logic;
signal il_max_comp1_wire : std_logic;
signal s2_phy_wire : std_logic;
signal il_min_comp2_wire : std_logic;
signal s1_phy_wire : std_logic;
signal s4_phy_wire : std_logic;
signal il_min_comp1_wire : std_logic;
signal s3_phy_wire : std_logic;
signal delay_hc_input_wire : std_logic;
signal delay_tr_input_wire : std_logic;
signal rgb_b_wire : std_logic;
signal rgb_g_wire : std_logic;
signal rgb_r_wire : std_logic;
signal \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ : std_logic_vector(15 downto 0);
signal \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\ : std_logic_vector(31 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ : std_logic_vector(15 downto 0);
signal \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\ : std_logic_vector(31 downto 0);

begin
    reset_wire <= reset;
    start_stop_wire <= start_stop;
    il_max_comp2_wire <= il_max_comp2;
    pwm_output <= pwm_output_wire;
    il_max_comp1_wire <= il_max_comp1;
    s2_phy <= s2_phy_wire;
    il_min_comp2_wire <= il_min_comp2;
    s1_phy <= s1_phy_wire;
    s4_phy <= s4_phy_wire;
    il_min_comp1_wire <= il_min_comp1;
    s3_phy <= s3_phy_wire;
    delay_hc_input_wire <= delay_hc_input;
    delay_tr_input_wire <= delay_tr_input;
    rgb_b <= rgb_b_wire;
    rgb_g <= rgb_g_wire;
    rgb_r <= rgb_r_wire;
    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\ <= \N__29838\&\N__29861\&\N__29499\&\N__29532\&\N__29565\&\N__29598\&\N__29624\&\N__29654\&\N__29685\&\N__29711\&\N__29270\&\N__29304\&\N__29334\&\N__29358\&\N__29391\&\N__29415\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38708\&'0'&\N__38707\;
    \current_shift_inst.PI_CTRL.integrator_1_0_2_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_1\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.integrator_1_0_2_0\ <= \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\ <= '0'&\N__48866\&\N__48859\&\N__48864\&\N__48858\&\N__48865\&\N__48857\&\N__48867\&\N__48854\&\N__48860\&\N__48853\&\N__48861\&\N__48855\&\N__48862\&\N__48856\&\N__48863\;
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38861\&\N__38858\&'0'&'0'&'0'&\N__38856\&\N__38860\&\N__38857\&\N__38859\;
    \pwm_generator_inst.un2_threshold_2_1_16\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_2_1_15\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.un2_threshold_2_14\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.un2_threshold_2_13\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.un2_threshold_2_12\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un2_threshold_2_11\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.un2_threshold_2_10\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.un2_threshold_2_9\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.un2_threshold_2_8\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.un2_threshold_2_7\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.un2_threshold_2_6\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.un2_threshold_2_5\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.un2_threshold_2_4\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.un2_threshold_2_3\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.un2_threshold_2_2\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.un2_threshold_2_1\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.un2_threshold_2_0\ <= \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\(0);
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\ <= '0'&\N__48835\&\N__48838\&\N__48836\&\N__48839\&\N__48837\&\N__20634\&\N__20565\&\N__20588\&\N__20613\&\N__20504\&\N__20526\&\N__20544\&\N__20232\&\N__20247\&\N__20211\;
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38676\&\N__38673\&'0'&'0'&'0'&\N__38671\&\N__38675\&\N__38672\&\N__38674\;
    \pwm_generator_inst.un2_threshold_1_25\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(25);
    \pwm_generator_inst.un2_threshold_1_24\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(24);
    \pwm_generator_inst.un2_threshold_1_23\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(23);
    \pwm_generator_inst.un2_threshold_1_22\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(22);
    \pwm_generator_inst.un2_threshold_1_21\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(21);
    \pwm_generator_inst.un2_threshold_1_20\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(20);
    \pwm_generator_inst.un2_threshold_1_19\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(19);
    \pwm_generator_inst.un2_threshold_1_18\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(18);
    \pwm_generator_inst.un2_threshold_1_17\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(17);
    \pwm_generator_inst.un2_threshold_1_16\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(16);
    \pwm_generator_inst.un2_threshold_1_15\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(15);
    \pwm_generator_inst.O_14\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(14);
    \pwm_generator_inst.O_13\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(13);
    \pwm_generator_inst.O_12\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(12);
    \pwm_generator_inst.un3_threshold\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(11);
    \pwm_generator_inst.O_10\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(10);
    \pwm_generator_inst.O_9\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(9);
    \pwm_generator_inst.O_8\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(8);
    \pwm_generator_inst.O_7\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(7);
    \pwm_generator_inst.O_6\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(6);
    \pwm_generator_inst.O_5\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(5);
    \pwm_generator_inst.O_4\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(4);
    \pwm_generator_inst.O_3\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(3);
    \pwm_generator_inst.O_2\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(2);
    \pwm_generator_inst.O_1\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(1);
    \pwm_generator_inst.O_0\ <= \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\(0);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\ <= '0'&\N__29445\&\N__29469\&\N__29010\&\N__29043\&\N__29076\&\N__29106\&\N__29139\&\N__29169\&\N__29193\&\N__29214\&\N__29243\&\N__28665\&\N__28695\&\N__28733\&\N__30807\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__38757\&'0'&\N__38756\;
    \current_shift_inst.PI_CTRL.integrator_1_0_1_19\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(19);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_18\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(18);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_17\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(17);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_16\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(16);
    \current_shift_inst.PI_CTRL.integrator_1_0_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(15);
    \current_shift_inst.PI_CTRL.integrator_1_15\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(14);
    \current_shift_inst.PI_CTRL.integrator_1_14\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(13);
    \current_shift_inst.PI_CTRL.integrator_1_13\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(12);
    \current_shift_inst.PI_CTRL.integrator_1_12\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(11);
    \current_shift_inst.PI_CTRL.integrator_1_11\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(10);
    \current_shift_inst.PI_CTRL.integrator_1_10\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(9);
    \current_shift_inst.PI_CTRL.integrator_1_9\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(8);
    \current_shift_inst.PI_CTRL.integrator_1_8\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(7);
    \current_shift_inst.PI_CTRL.integrator_1_7\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(6);
    \current_shift_inst.PI_CTRL.integrator_1_6\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(5);
    \current_shift_inst.PI_CTRL.integrator_1_5\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(4);
    \current_shift_inst.PI_CTRL.integrator_1_4\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(3);
    \current_shift_inst.PI_CTRL.integrator_1_3\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(2);
    \current_shift_inst.PI_CTRL.integrator_1_2\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(1);
    \current_shift_inst.PI_CTRL.un1_integrator\ <= \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\(0);

    \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__27351\,
            RESETB => \N__33516\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => clk_100mhz_0
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38709\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38706\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38862\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38855\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_2_1_mulonly_0_25_0_O_wire\
        );

    \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38677\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38670\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_D_wire\,
            ADDSUBBOT => '0',
            A => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_A_wire\,
            C => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_C_wire\,
            B => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_B_wire\,
            OHOLDTOP => '0',
            O => \pwm_generator_inst.un2_threshold_1_mulonly_0_25_0_O_wire\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0\ : SB_MAC16
    generic map (
            A_REG => '0',
            TOP_8x8_MULT_REG => '0',
            TOPOUTPUT_SELECT => "11",
            TOPADDSUB_UPPERINPUT => '0',
            TOPADDSUB_LOWERINPUT => "00",
            TOPADDSUB_CARRYSELECT => "00",
            PIPELINE_16x16_MULT_REG2 => '0',
            PIPELINE_16x16_MULT_REG1 => '0',
            NEG_TRIGGER => '0',
            MODE_8x8 => '0',
            D_REG => '0',
            C_REG => '0',
            B_SIGNED => '1',
            B_REG => '0',
            BOT_8x8_MULT_REG => '0',
            BOTOUTPUT_SELECT => "11",
            BOTADDSUB_UPPERINPUT => '0',
            BOTADDSUB_LOWERINPUT => "00",
            BOTADDSUB_CARRYSELECT => "00",
            A_SIGNED => '1'
        )
    port map (
            ACCUMCO => OPEN,
            DHOLD => '0',
            AHOLD => \N__38758\,
            SIGNEXTOUT => OPEN,
            ORSTTOP => '0',
            ORSTBOT => '0',
            CI => '0',
            IRSTTOP => '0',
            ACCUMCI => '0',
            OLOADBOT => '0',
            CHOLD => '0',
            IRSTBOT => '0',
            OHOLDBOT => '0',
            SIGNEXTIN => '0',
            ADDSUBTOP => '0',
            OLOADTOP => '0',
            CE => 'H',
            BHOLD => \N__38755\,
            CLK => \GNDG0\,
            CO => OPEN,
            D => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_D_wire\,
            ADDSUBBOT => '0',
            A => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_A_wire\,
            C => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_C_wire\,
            B => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_B_wire\,
            OHOLDTOP => '0',
            O => \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0_O_wire\
        );

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__50509\,
            GLOBALBUFFEROUTPUT => red_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50511\,
            DIN => \N__50510\,
            DOUT => \N__50509\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50511\,
            PADOUT => \N__50510\,
            PADIN => \N__50509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start_stop_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50500\,
            DIN => \N__50499\,
            DOUT => \N__50498\,
            PACKAGEPIN => start_stop_wire
        );

    \start_stop_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50500\,
            PADOUT => \N__50499\,
            PADIN => \N__50498\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => start_stop_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50491\,
            DIN => \N__50490\,
            DOUT => \N__50489\,
            PACKAGEPIN => il_max_comp2_wire
        );

    \il_max_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50491\,
            PADOUT => \N__50490\,
            PADIN => \N__50489\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_output_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50482\,
            DIN => \N__50481\,
            DOUT => \N__50480\,
            PACKAGEPIN => pwm_output_wire
        );

    \pwm_output_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50482\,
            PADOUT => \N__50481\,
            PADIN => \N__50480\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__27201\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_max_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50473\,
            DIN => \N__50472\,
            DOUT => \N__50471\,
            PACKAGEPIN => il_max_comp1_wire
        );

    \il_max_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50473\,
            PADOUT => \N__50472\,
            PADIN => \N__50471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_max_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50464\,
            DIN => \N__50463\,
            DOUT => \N__50462\,
            PACKAGEPIN => s2_phy_wire
        );

    \s2_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50464\,
            PADOUT => \N__50463\,
            PADIN => \N__50462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34926\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50455\,
            DIN => \N__50454\,
            DOUT => \N__50453\,
            PACKAGEPIN => il_min_comp2_wire
        );

    \il_min_comp2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50455\,
            PADOUT => \N__50454\,
            PADIN => \N__50453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp2_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50446\,
            DIN => \N__50445\,
            DOUT => \N__50444\,
            PACKAGEPIN => s1_phy_wire
        );

    \s1_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50446\,
            PADOUT => \N__50445\,
            PADIN => \N__50444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__34869\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s4_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50437\,
            DIN => \N__50436\,
            DOUT => \N__50435\,
            PACKAGEPIN => s4_phy_wire
        );

    \s4_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50437\,
            PADOUT => \N__50436\,
            PADIN => \N__50435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__32355\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \il_min_comp1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50428\,
            DIN => \N__50427\,
            DOUT => \N__50426\,
            PACKAGEPIN => il_min_comp1_wire
        );

    \il_min_comp1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50428\,
            PADOUT => \N__50427\,
            PADIN => \N__50426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => il_min_comp1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_phy_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50419\,
            DIN => \N__50418\,
            DOUT => \N__50417\,
            PACKAGEPIN => s3_phy_wire
        );

    \s3_phy_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__50419\,
            PADOUT => \N__50418\,
            PADIN => \N__50417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33534\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_hc_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50410\,
            DIN => \N__50409\,
            DOUT => \N__50408\,
            PACKAGEPIN => delay_hc_input_wire
        );

    \delay_hc_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50410\,
            PADOUT => \N__50409\,
            PADIN => \N__50408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_hc_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \delay_tr_input_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__50401\,
            DIN => \N__50400\,
            DOUT => \N__50399\,
            PACKAGEPIN => delay_tr_input_wire
        );

    \delay_tr_input_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__50401\,
            PADOUT => \N__50400\,
            PADIN => \N__50399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => delay_tr_input_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__12029\ : InMux
    port map (
            O => \N__50382\,
            I => \N__50379\
        );

    \I__12028\ : LocalMux
    port map (
            O => \N__50379\,
            I => \N__50376\
        );

    \I__12027\ : Span4Mux_v
    port map (
            O => \N__50376\,
            I => \N__50372\
        );

    \I__12026\ : InMux
    port map (
            O => \N__50375\,
            I => \N__50368\
        );

    \I__12025\ : Span4Mux_h
    port map (
            O => \N__50372\,
            I => \N__50365\
        );

    \I__12024\ : InMux
    port map (
            O => \N__50371\,
            I => \N__50362\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__50368\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__12022\ : Odrv4
    port map (
            O => \N__50365\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__12021\ : LocalMux
    port map (
            O => \N__50362\,
            I => \elapsed_time_ns_1_RNI58DN9_0_27\
        );

    \I__12020\ : CascadeMux
    port map (
            O => \N__50355\,
            I => \N__50352\
        );

    \I__12019\ : InMux
    port map (
            O => \N__50352\,
            I => \N__50348\
        );

    \I__12018\ : InMux
    port map (
            O => \N__50351\,
            I => \N__50345\
        );

    \I__12017\ : LocalMux
    port map (
            O => \N__50348\,
            I => \N__50341\
        );

    \I__12016\ : LocalMux
    port map (
            O => \N__50345\,
            I => \N__50338\
        );

    \I__12015\ : InMux
    port map (
            O => \N__50344\,
            I => \N__50335\
        );

    \I__12014\ : Span4Mux_v
    port map (
            O => \N__50341\,
            I => \N__50332\
        );

    \I__12013\ : Odrv4
    port map (
            O => \N__50338\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__50335\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__12011\ : Odrv4
    port map (
            O => \N__50332\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\
        );

    \I__12010\ : InMux
    port map (
            O => \N__50325\,
            I => \N__50320\
        );

    \I__12009\ : InMux
    port map (
            O => \N__50324\,
            I => \N__50316\
        );

    \I__12008\ : InMux
    port map (
            O => \N__50323\,
            I => \N__50313\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__50320\,
            I => \N__50310\
        );

    \I__12006\ : InMux
    port map (
            O => \N__50319\,
            I => \N__50307\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__50316\,
            I => \N__50304\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__50313\,
            I => \N__50301\
        );

    \I__12003\ : Span4Mux_v
    port map (
            O => \N__50310\,
            I => \N__50296\
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50307\,
            I => \N__50296\
        );

    \I__12001\ : Span4Mux_h
    port map (
            O => \N__50304\,
            I => \N__50293\
        );

    \I__12000\ : Span4Mux_v
    port map (
            O => \N__50301\,
            I => \N__50288\
        );

    \I__11999\ : Span4Mux_h
    port map (
            O => \N__50296\,
            I => \N__50288\
        );

    \I__11998\ : Odrv4
    port map (
            O => \N__50293\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__11997\ : Odrv4
    port map (
            O => \N__50288\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\
        );

    \I__11996\ : CEMux
    port map (
            O => \N__50283\,
            I => \N__50280\
        );

    \I__11995\ : LocalMux
    port map (
            O => \N__50280\,
            I => \N__50274\
        );

    \I__11994\ : CEMux
    port map (
            O => \N__50279\,
            I => \N__50271\
        );

    \I__11993\ : CEMux
    port map (
            O => \N__50278\,
            I => \N__50268\
        );

    \I__11992\ : CEMux
    port map (
            O => \N__50277\,
            I => \N__50265\
        );

    \I__11991\ : Span4Mux_v
    port map (
            O => \N__50274\,
            I => \N__50260\
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__50271\,
            I => \N__50260\
        );

    \I__11989\ : LocalMux
    port map (
            O => \N__50268\,
            I => \N__50257\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__50265\,
            I => \N__50254\
        );

    \I__11987\ : Span4Mux_v
    port map (
            O => \N__50260\,
            I => \N__50251\
        );

    \I__11986\ : Span4Mux_h
    port map (
            O => \N__50257\,
            I => \N__50248\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__50254\,
            I => \N__50245\
        );

    \I__11984\ : Odrv4
    port map (
            O => \N__50251\,
            I => \delay_measurement_inst.delay_hc_timer.N_164_i\
        );

    \I__11983\ : Odrv4
    port map (
            O => \N__50248\,
            I => \delay_measurement_inst.delay_hc_timer.N_164_i\
        );

    \I__11982\ : Odrv4
    port map (
            O => \N__50245\,
            I => \delay_measurement_inst.delay_hc_timer.N_164_i\
        );

    \I__11981\ : CEMux
    port map (
            O => \N__50238\,
            I => \N__50235\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__50235\,
            I => \N__50230\
        );

    \I__11979\ : CEMux
    port map (
            O => \N__50234\,
            I => \N__50227\
        );

    \I__11978\ : CEMux
    port map (
            O => \N__50233\,
            I => \N__50223\
        );

    \I__11977\ : Span4Mux_v
    port map (
            O => \N__50230\,
            I => \N__50218\
        );

    \I__11976\ : LocalMux
    port map (
            O => \N__50227\,
            I => \N__50218\
        );

    \I__11975\ : CEMux
    port map (
            O => \N__50226\,
            I => \N__50215\
        );

    \I__11974\ : LocalMux
    port map (
            O => \N__50223\,
            I => \N__50211\
        );

    \I__11973\ : Span4Mux_h
    port map (
            O => \N__50218\,
            I => \N__50208\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__50215\,
            I => \N__50205\
        );

    \I__11971\ : CEMux
    port map (
            O => \N__50214\,
            I => \N__50202\
        );

    \I__11970\ : Span4Mux_h
    port map (
            O => \N__50211\,
            I => \N__50199\
        );

    \I__11969\ : Span4Mux_h
    port map (
            O => \N__50208\,
            I => \N__50196\
        );

    \I__11968\ : Span4Mux_h
    port map (
            O => \N__50205\,
            I => \N__50191\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__50202\,
            I => \N__50191\
        );

    \I__11966\ : Odrv4
    port map (
            O => \N__50199\,
            I => \delay_measurement_inst.delay_hc_timer.N_163_i\
        );

    \I__11965\ : Odrv4
    port map (
            O => \N__50196\,
            I => \delay_measurement_inst.delay_hc_timer.N_163_i\
        );

    \I__11964\ : Odrv4
    port map (
            O => \N__50191\,
            I => \delay_measurement_inst.delay_hc_timer.N_163_i\
        );

    \I__11963\ : InMux
    port map (
            O => \N__50184\,
            I => \N__50150\
        );

    \I__11962\ : InMux
    port map (
            O => \N__50183\,
            I => \N__50150\
        );

    \I__11961\ : InMux
    port map (
            O => \N__50182\,
            I => \N__50150\
        );

    \I__11960\ : InMux
    port map (
            O => \N__50181\,
            I => \N__50150\
        );

    \I__11959\ : InMux
    port map (
            O => \N__50180\,
            I => \N__50137\
        );

    \I__11958\ : InMux
    port map (
            O => \N__50179\,
            I => \N__50137\
        );

    \I__11957\ : InMux
    port map (
            O => \N__50178\,
            I => \N__50137\
        );

    \I__11956\ : InMux
    port map (
            O => \N__50177\,
            I => \N__50137\
        );

    \I__11955\ : InMux
    port map (
            O => \N__50176\,
            I => \N__50128\
        );

    \I__11954\ : InMux
    port map (
            O => \N__50175\,
            I => \N__50128\
        );

    \I__11953\ : InMux
    port map (
            O => \N__50174\,
            I => \N__50128\
        );

    \I__11952\ : InMux
    port map (
            O => \N__50173\,
            I => \N__50128\
        );

    \I__11951\ : InMux
    port map (
            O => \N__50172\,
            I => \N__50123\
        );

    \I__11950\ : InMux
    port map (
            O => \N__50171\,
            I => \N__50123\
        );

    \I__11949\ : InMux
    port map (
            O => \N__50170\,
            I => \N__50114\
        );

    \I__11948\ : InMux
    port map (
            O => \N__50169\,
            I => \N__50114\
        );

    \I__11947\ : InMux
    port map (
            O => \N__50168\,
            I => \N__50114\
        );

    \I__11946\ : InMux
    port map (
            O => \N__50167\,
            I => \N__50114\
        );

    \I__11945\ : InMux
    port map (
            O => \N__50166\,
            I => \N__50105\
        );

    \I__11944\ : InMux
    port map (
            O => \N__50165\,
            I => \N__50105\
        );

    \I__11943\ : InMux
    port map (
            O => \N__50164\,
            I => \N__50105\
        );

    \I__11942\ : InMux
    port map (
            O => \N__50163\,
            I => \N__50105\
        );

    \I__11941\ : InMux
    port map (
            O => \N__50162\,
            I => \N__50096\
        );

    \I__11940\ : InMux
    port map (
            O => \N__50161\,
            I => \N__50096\
        );

    \I__11939\ : InMux
    port map (
            O => \N__50160\,
            I => \N__50096\
        );

    \I__11938\ : InMux
    port map (
            O => \N__50159\,
            I => \N__50096\
        );

    \I__11937\ : LocalMux
    port map (
            O => \N__50150\,
            I => \N__50093\
        );

    \I__11936\ : InMux
    port map (
            O => \N__50149\,
            I => \N__50084\
        );

    \I__11935\ : InMux
    port map (
            O => \N__50148\,
            I => \N__50084\
        );

    \I__11934\ : InMux
    port map (
            O => \N__50147\,
            I => \N__50084\
        );

    \I__11933\ : InMux
    port map (
            O => \N__50146\,
            I => \N__50084\
        );

    \I__11932\ : LocalMux
    port map (
            O => \N__50137\,
            I => \N__50079\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__50128\,
            I => \N__50079\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__50123\,
            I => \N__50076\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__50114\,
            I => \N__50073\
        );

    \I__11928\ : LocalMux
    port map (
            O => \N__50105\,
            I => \N__50068\
        );

    \I__11927\ : LocalMux
    port map (
            O => \N__50096\,
            I => \N__50068\
        );

    \I__11926\ : Span4Mux_v
    port map (
            O => \N__50093\,
            I => \N__50063\
        );

    \I__11925\ : LocalMux
    port map (
            O => \N__50084\,
            I => \N__50063\
        );

    \I__11924\ : Span4Mux_h
    port map (
            O => \N__50079\,
            I => \N__50060\
        );

    \I__11923\ : Span4Mux_h
    port map (
            O => \N__50076\,
            I => \N__50055\
        );

    \I__11922\ : Span4Mux_h
    port map (
            O => \N__50073\,
            I => \N__50055\
        );

    \I__11921\ : Span4Mux_h
    port map (
            O => \N__50068\,
            I => \N__50052\
        );

    \I__11920\ : Odrv4
    port map (
            O => \N__50063\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11919\ : Odrv4
    port map (
            O => \N__50060\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11918\ : Odrv4
    port map (
            O => \N__50055\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11917\ : Odrv4
    port map (
            O => \N__50052\,
            I => \delay_measurement_inst.delay_hc_timer.running_i\
        );

    \I__11916\ : InMux
    port map (
            O => \N__50043\,
            I => \N__50039\
        );

    \I__11915\ : CascadeMux
    port map (
            O => \N__50042\,
            I => \N__50036\
        );

    \I__11914\ : LocalMux
    port map (
            O => \N__50039\,
            I => \N__50032\
        );

    \I__11913\ : InMux
    port map (
            O => \N__50036\,
            I => \N__50027\
        );

    \I__11912\ : InMux
    port map (
            O => \N__50035\,
            I => \N__50027\
        );

    \I__11911\ : Span4Mux_v
    port map (
            O => \N__50032\,
            I => \N__50022\
        );

    \I__11910\ : LocalMux
    port map (
            O => \N__50027\,
            I => \N__50022\
        );

    \I__11909\ : Span4Mux_h
    port map (
            O => \N__50022\,
            I => \N__50019\
        );

    \I__11908\ : Span4Mux_h
    port map (
            O => \N__50019\,
            I => \N__50016\
        );

    \I__11907\ : Span4Mux_v
    port map (
            O => \N__50016\,
            I => \N__50013\
        );

    \I__11906\ : Odrv4
    port map (
            O => \N__50013\,
            I => \delay_measurement_inst.stop_timer_hcZ0\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50010\,
            I => \N__50007\
        );

    \I__11904\ : LocalMux
    port map (
            O => \N__50007\,
            I => \N__50003\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50006\,
            I => \N__50000\
        );

    \I__11902\ : Span4Mux_v
    port map (
            O => \N__50003\,
            I => \N__49995\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__50000\,
            I => \N__49995\
        );

    \I__11900\ : Span4Mux_h
    port map (
            O => \N__49995\,
            I => \N__49992\
        );

    \I__11899\ : Span4Mux_h
    port map (
            O => \N__49992\,
            I => \N__49987\
        );

    \I__11898\ : InMux
    port map (
            O => \N__49991\,
            I => \N__49982\
        );

    \I__11897\ : InMux
    port map (
            O => \N__49990\,
            I => \N__49982\
        );

    \I__11896\ : Span4Mux_v
    port map (
            O => \N__49987\,
            I => \N__49979\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__49982\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__11894\ : Odrv4
    port map (
            O => \N__49979\,
            I => \delay_measurement_inst.start_timer_hcZ0\
        );

    \I__11893\ : InMux
    port map (
            O => \N__49974\,
            I => \N__49968\
        );

    \I__11892\ : InMux
    port map (
            O => \N__49973\,
            I => \N__49961\
        );

    \I__11891\ : InMux
    port map (
            O => \N__49972\,
            I => \N__49961\
        );

    \I__11890\ : InMux
    port map (
            O => \N__49971\,
            I => \N__49961\
        );

    \I__11889\ : LocalMux
    port map (
            O => \N__49968\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__11888\ : LocalMux
    port map (
            O => \N__49961\,
            I => \delay_measurement_inst.delay_hc_timer.runningZ0\
        );

    \I__11887\ : ClkMux
    port map (
            O => \N__49956\,
            I => \N__49482\
        );

    \I__11886\ : ClkMux
    port map (
            O => \N__49955\,
            I => \N__49482\
        );

    \I__11885\ : ClkMux
    port map (
            O => \N__49954\,
            I => \N__49482\
        );

    \I__11884\ : ClkMux
    port map (
            O => \N__49953\,
            I => \N__49482\
        );

    \I__11883\ : ClkMux
    port map (
            O => \N__49952\,
            I => \N__49482\
        );

    \I__11882\ : ClkMux
    port map (
            O => \N__49951\,
            I => \N__49482\
        );

    \I__11881\ : ClkMux
    port map (
            O => \N__49950\,
            I => \N__49482\
        );

    \I__11880\ : ClkMux
    port map (
            O => \N__49949\,
            I => \N__49482\
        );

    \I__11879\ : ClkMux
    port map (
            O => \N__49948\,
            I => \N__49482\
        );

    \I__11878\ : ClkMux
    port map (
            O => \N__49947\,
            I => \N__49482\
        );

    \I__11877\ : ClkMux
    port map (
            O => \N__49946\,
            I => \N__49482\
        );

    \I__11876\ : ClkMux
    port map (
            O => \N__49945\,
            I => \N__49482\
        );

    \I__11875\ : ClkMux
    port map (
            O => \N__49944\,
            I => \N__49482\
        );

    \I__11874\ : ClkMux
    port map (
            O => \N__49943\,
            I => \N__49482\
        );

    \I__11873\ : ClkMux
    port map (
            O => \N__49942\,
            I => \N__49482\
        );

    \I__11872\ : ClkMux
    port map (
            O => \N__49941\,
            I => \N__49482\
        );

    \I__11871\ : ClkMux
    port map (
            O => \N__49940\,
            I => \N__49482\
        );

    \I__11870\ : ClkMux
    port map (
            O => \N__49939\,
            I => \N__49482\
        );

    \I__11869\ : ClkMux
    port map (
            O => \N__49938\,
            I => \N__49482\
        );

    \I__11868\ : ClkMux
    port map (
            O => \N__49937\,
            I => \N__49482\
        );

    \I__11867\ : ClkMux
    port map (
            O => \N__49936\,
            I => \N__49482\
        );

    \I__11866\ : ClkMux
    port map (
            O => \N__49935\,
            I => \N__49482\
        );

    \I__11865\ : ClkMux
    port map (
            O => \N__49934\,
            I => \N__49482\
        );

    \I__11864\ : ClkMux
    port map (
            O => \N__49933\,
            I => \N__49482\
        );

    \I__11863\ : ClkMux
    port map (
            O => \N__49932\,
            I => \N__49482\
        );

    \I__11862\ : ClkMux
    port map (
            O => \N__49931\,
            I => \N__49482\
        );

    \I__11861\ : ClkMux
    port map (
            O => \N__49930\,
            I => \N__49482\
        );

    \I__11860\ : ClkMux
    port map (
            O => \N__49929\,
            I => \N__49482\
        );

    \I__11859\ : ClkMux
    port map (
            O => \N__49928\,
            I => \N__49482\
        );

    \I__11858\ : ClkMux
    port map (
            O => \N__49927\,
            I => \N__49482\
        );

    \I__11857\ : ClkMux
    port map (
            O => \N__49926\,
            I => \N__49482\
        );

    \I__11856\ : ClkMux
    port map (
            O => \N__49925\,
            I => \N__49482\
        );

    \I__11855\ : ClkMux
    port map (
            O => \N__49924\,
            I => \N__49482\
        );

    \I__11854\ : ClkMux
    port map (
            O => \N__49923\,
            I => \N__49482\
        );

    \I__11853\ : ClkMux
    port map (
            O => \N__49922\,
            I => \N__49482\
        );

    \I__11852\ : ClkMux
    port map (
            O => \N__49921\,
            I => \N__49482\
        );

    \I__11851\ : ClkMux
    port map (
            O => \N__49920\,
            I => \N__49482\
        );

    \I__11850\ : ClkMux
    port map (
            O => \N__49919\,
            I => \N__49482\
        );

    \I__11849\ : ClkMux
    port map (
            O => \N__49918\,
            I => \N__49482\
        );

    \I__11848\ : ClkMux
    port map (
            O => \N__49917\,
            I => \N__49482\
        );

    \I__11847\ : ClkMux
    port map (
            O => \N__49916\,
            I => \N__49482\
        );

    \I__11846\ : ClkMux
    port map (
            O => \N__49915\,
            I => \N__49482\
        );

    \I__11845\ : ClkMux
    port map (
            O => \N__49914\,
            I => \N__49482\
        );

    \I__11844\ : ClkMux
    port map (
            O => \N__49913\,
            I => \N__49482\
        );

    \I__11843\ : ClkMux
    port map (
            O => \N__49912\,
            I => \N__49482\
        );

    \I__11842\ : ClkMux
    port map (
            O => \N__49911\,
            I => \N__49482\
        );

    \I__11841\ : ClkMux
    port map (
            O => \N__49910\,
            I => \N__49482\
        );

    \I__11840\ : ClkMux
    port map (
            O => \N__49909\,
            I => \N__49482\
        );

    \I__11839\ : ClkMux
    port map (
            O => \N__49908\,
            I => \N__49482\
        );

    \I__11838\ : ClkMux
    port map (
            O => \N__49907\,
            I => \N__49482\
        );

    \I__11837\ : ClkMux
    port map (
            O => \N__49906\,
            I => \N__49482\
        );

    \I__11836\ : ClkMux
    port map (
            O => \N__49905\,
            I => \N__49482\
        );

    \I__11835\ : ClkMux
    port map (
            O => \N__49904\,
            I => \N__49482\
        );

    \I__11834\ : ClkMux
    port map (
            O => \N__49903\,
            I => \N__49482\
        );

    \I__11833\ : ClkMux
    port map (
            O => \N__49902\,
            I => \N__49482\
        );

    \I__11832\ : ClkMux
    port map (
            O => \N__49901\,
            I => \N__49482\
        );

    \I__11831\ : ClkMux
    port map (
            O => \N__49900\,
            I => \N__49482\
        );

    \I__11830\ : ClkMux
    port map (
            O => \N__49899\,
            I => \N__49482\
        );

    \I__11829\ : ClkMux
    port map (
            O => \N__49898\,
            I => \N__49482\
        );

    \I__11828\ : ClkMux
    port map (
            O => \N__49897\,
            I => \N__49482\
        );

    \I__11827\ : ClkMux
    port map (
            O => \N__49896\,
            I => \N__49482\
        );

    \I__11826\ : ClkMux
    port map (
            O => \N__49895\,
            I => \N__49482\
        );

    \I__11825\ : ClkMux
    port map (
            O => \N__49894\,
            I => \N__49482\
        );

    \I__11824\ : ClkMux
    port map (
            O => \N__49893\,
            I => \N__49482\
        );

    \I__11823\ : ClkMux
    port map (
            O => \N__49892\,
            I => \N__49482\
        );

    \I__11822\ : ClkMux
    port map (
            O => \N__49891\,
            I => \N__49482\
        );

    \I__11821\ : ClkMux
    port map (
            O => \N__49890\,
            I => \N__49482\
        );

    \I__11820\ : ClkMux
    port map (
            O => \N__49889\,
            I => \N__49482\
        );

    \I__11819\ : ClkMux
    port map (
            O => \N__49888\,
            I => \N__49482\
        );

    \I__11818\ : ClkMux
    port map (
            O => \N__49887\,
            I => \N__49482\
        );

    \I__11817\ : ClkMux
    port map (
            O => \N__49886\,
            I => \N__49482\
        );

    \I__11816\ : ClkMux
    port map (
            O => \N__49885\,
            I => \N__49482\
        );

    \I__11815\ : ClkMux
    port map (
            O => \N__49884\,
            I => \N__49482\
        );

    \I__11814\ : ClkMux
    port map (
            O => \N__49883\,
            I => \N__49482\
        );

    \I__11813\ : ClkMux
    port map (
            O => \N__49882\,
            I => \N__49482\
        );

    \I__11812\ : ClkMux
    port map (
            O => \N__49881\,
            I => \N__49482\
        );

    \I__11811\ : ClkMux
    port map (
            O => \N__49880\,
            I => \N__49482\
        );

    \I__11810\ : ClkMux
    port map (
            O => \N__49879\,
            I => \N__49482\
        );

    \I__11809\ : ClkMux
    port map (
            O => \N__49878\,
            I => \N__49482\
        );

    \I__11808\ : ClkMux
    port map (
            O => \N__49877\,
            I => \N__49482\
        );

    \I__11807\ : ClkMux
    port map (
            O => \N__49876\,
            I => \N__49482\
        );

    \I__11806\ : ClkMux
    port map (
            O => \N__49875\,
            I => \N__49482\
        );

    \I__11805\ : ClkMux
    port map (
            O => \N__49874\,
            I => \N__49482\
        );

    \I__11804\ : ClkMux
    port map (
            O => \N__49873\,
            I => \N__49482\
        );

    \I__11803\ : ClkMux
    port map (
            O => \N__49872\,
            I => \N__49482\
        );

    \I__11802\ : ClkMux
    port map (
            O => \N__49871\,
            I => \N__49482\
        );

    \I__11801\ : ClkMux
    port map (
            O => \N__49870\,
            I => \N__49482\
        );

    \I__11800\ : ClkMux
    port map (
            O => \N__49869\,
            I => \N__49482\
        );

    \I__11799\ : ClkMux
    port map (
            O => \N__49868\,
            I => \N__49482\
        );

    \I__11798\ : ClkMux
    port map (
            O => \N__49867\,
            I => \N__49482\
        );

    \I__11797\ : ClkMux
    port map (
            O => \N__49866\,
            I => \N__49482\
        );

    \I__11796\ : ClkMux
    port map (
            O => \N__49865\,
            I => \N__49482\
        );

    \I__11795\ : ClkMux
    port map (
            O => \N__49864\,
            I => \N__49482\
        );

    \I__11794\ : ClkMux
    port map (
            O => \N__49863\,
            I => \N__49482\
        );

    \I__11793\ : ClkMux
    port map (
            O => \N__49862\,
            I => \N__49482\
        );

    \I__11792\ : ClkMux
    port map (
            O => \N__49861\,
            I => \N__49482\
        );

    \I__11791\ : ClkMux
    port map (
            O => \N__49860\,
            I => \N__49482\
        );

    \I__11790\ : ClkMux
    port map (
            O => \N__49859\,
            I => \N__49482\
        );

    \I__11789\ : ClkMux
    port map (
            O => \N__49858\,
            I => \N__49482\
        );

    \I__11788\ : ClkMux
    port map (
            O => \N__49857\,
            I => \N__49482\
        );

    \I__11787\ : ClkMux
    port map (
            O => \N__49856\,
            I => \N__49482\
        );

    \I__11786\ : ClkMux
    port map (
            O => \N__49855\,
            I => \N__49482\
        );

    \I__11785\ : ClkMux
    port map (
            O => \N__49854\,
            I => \N__49482\
        );

    \I__11784\ : ClkMux
    port map (
            O => \N__49853\,
            I => \N__49482\
        );

    \I__11783\ : ClkMux
    port map (
            O => \N__49852\,
            I => \N__49482\
        );

    \I__11782\ : ClkMux
    port map (
            O => \N__49851\,
            I => \N__49482\
        );

    \I__11781\ : ClkMux
    port map (
            O => \N__49850\,
            I => \N__49482\
        );

    \I__11780\ : ClkMux
    port map (
            O => \N__49849\,
            I => \N__49482\
        );

    \I__11779\ : ClkMux
    port map (
            O => \N__49848\,
            I => \N__49482\
        );

    \I__11778\ : ClkMux
    port map (
            O => \N__49847\,
            I => \N__49482\
        );

    \I__11777\ : ClkMux
    port map (
            O => \N__49846\,
            I => \N__49482\
        );

    \I__11776\ : ClkMux
    port map (
            O => \N__49845\,
            I => \N__49482\
        );

    \I__11775\ : ClkMux
    port map (
            O => \N__49844\,
            I => \N__49482\
        );

    \I__11774\ : ClkMux
    port map (
            O => \N__49843\,
            I => \N__49482\
        );

    \I__11773\ : ClkMux
    port map (
            O => \N__49842\,
            I => \N__49482\
        );

    \I__11772\ : ClkMux
    port map (
            O => \N__49841\,
            I => \N__49482\
        );

    \I__11771\ : ClkMux
    port map (
            O => \N__49840\,
            I => \N__49482\
        );

    \I__11770\ : ClkMux
    port map (
            O => \N__49839\,
            I => \N__49482\
        );

    \I__11769\ : ClkMux
    port map (
            O => \N__49838\,
            I => \N__49482\
        );

    \I__11768\ : ClkMux
    port map (
            O => \N__49837\,
            I => \N__49482\
        );

    \I__11767\ : ClkMux
    port map (
            O => \N__49836\,
            I => \N__49482\
        );

    \I__11766\ : ClkMux
    port map (
            O => \N__49835\,
            I => \N__49482\
        );

    \I__11765\ : ClkMux
    port map (
            O => \N__49834\,
            I => \N__49482\
        );

    \I__11764\ : ClkMux
    port map (
            O => \N__49833\,
            I => \N__49482\
        );

    \I__11763\ : ClkMux
    port map (
            O => \N__49832\,
            I => \N__49482\
        );

    \I__11762\ : ClkMux
    port map (
            O => \N__49831\,
            I => \N__49482\
        );

    \I__11761\ : ClkMux
    port map (
            O => \N__49830\,
            I => \N__49482\
        );

    \I__11760\ : ClkMux
    port map (
            O => \N__49829\,
            I => \N__49482\
        );

    \I__11759\ : ClkMux
    port map (
            O => \N__49828\,
            I => \N__49482\
        );

    \I__11758\ : ClkMux
    port map (
            O => \N__49827\,
            I => \N__49482\
        );

    \I__11757\ : ClkMux
    port map (
            O => \N__49826\,
            I => \N__49482\
        );

    \I__11756\ : ClkMux
    port map (
            O => \N__49825\,
            I => \N__49482\
        );

    \I__11755\ : ClkMux
    port map (
            O => \N__49824\,
            I => \N__49482\
        );

    \I__11754\ : ClkMux
    port map (
            O => \N__49823\,
            I => \N__49482\
        );

    \I__11753\ : ClkMux
    port map (
            O => \N__49822\,
            I => \N__49482\
        );

    \I__11752\ : ClkMux
    port map (
            O => \N__49821\,
            I => \N__49482\
        );

    \I__11751\ : ClkMux
    port map (
            O => \N__49820\,
            I => \N__49482\
        );

    \I__11750\ : ClkMux
    port map (
            O => \N__49819\,
            I => \N__49482\
        );

    \I__11749\ : ClkMux
    port map (
            O => \N__49818\,
            I => \N__49482\
        );

    \I__11748\ : ClkMux
    port map (
            O => \N__49817\,
            I => \N__49482\
        );

    \I__11747\ : ClkMux
    port map (
            O => \N__49816\,
            I => \N__49482\
        );

    \I__11746\ : ClkMux
    port map (
            O => \N__49815\,
            I => \N__49482\
        );

    \I__11745\ : ClkMux
    port map (
            O => \N__49814\,
            I => \N__49482\
        );

    \I__11744\ : ClkMux
    port map (
            O => \N__49813\,
            I => \N__49482\
        );

    \I__11743\ : ClkMux
    port map (
            O => \N__49812\,
            I => \N__49482\
        );

    \I__11742\ : ClkMux
    port map (
            O => \N__49811\,
            I => \N__49482\
        );

    \I__11741\ : ClkMux
    port map (
            O => \N__49810\,
            I => \N__49482\
        );

    \I__11740\ : ClkMux
    port map (
            O => \N__49809\,
            I => \N__49482\
        );

    \I__11739\ : ClkMux
    port map (
            O => \N__49808\,
            I => \N__49482\
        );

    \I__11738\ : ClkMux
    port map (
            O => \N__49807\,
            I => \N__49482\
        );

    \I__11737\ : ClkMux
    port map (
            O => \N__49806\,
            I => \N__49482\
        );

    \I__11736\ : ClkMux
    port map (
            O => \N__49805\,
            I => \N__49482\
        );

    \I__11735\ : ClkMux
    port map (
            O => \N__49804\,
            I => \N__49482\
        );

    \I__11734\ : ClkMux
    port map (
            O => \N__49803\,
            I => \N__49482\
        );

    \I__11733\ : ClkMux
    port map (
            O => \N__49802\,
            I => \N__49482\
        );

    \I__11732\ : ClkMux
    port map (
            O => \N__49801\,
            I => \N__49482\
        );

    \I__11731\ : ClkMux
    port map (
            O => \N__49800\,
            I => \N__49482\
        );

    \I__11730\ : ClkMux
    port map (
            O => \N__49799\,
            I => \N__49482\
        );

    \I__11729\ : GlobalMux
    port map (
            O => \N__49482\,
            I => clk_100mhz_0
        );

    \I__11728\ : InMux
    port map (
            O => \N__49479\,
            I => \N__49473\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49478\,
            I => \N__49470\
        );

    \I__11726\ : InMux
    port map (
            O => \N__49477\,
            I => \N__49467\
        );

    \I__11725\ : InMux
    port map (
            O => \N__49476\,
            I => \N__49464\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__49473\,
            I => \N__49461\
        );

    \I__11723\ : LocalMux
    port map (
            O => \N__49470\,
            I => \N__49458\
        );

    \I__11722\ : LocalMux
    port map (
            O => \N__49467\,
            I => \N__49455\
        );

    \I__11721\ : LocalMux
    port map (
            O => \N__49464\,
            I => \N__49447\
        );

    \I__11720\ : Glb2LocalMux
    port map (
            O => \N__49461\,
            I => \N__48960\
        );

    \I__11719\ : Glb2LocalMux
    port map (
            O => \N__49458\,
            I => \N__48960\
        );

    \I__11718\ : Glb2LocalMux
    port map (
            O => \N__49455\,
            I => \N__48960\
        );

    \I__11717\ : SRMux
    port map (
            O => \N__49454\,
            I => \N__48960\
        );

    \I__11716\ : SRMux
    port map (
            O => \N__49453\,
            I => \N__48960\
        );

    \I__11715\ : SRMux
    port map (
            O => \N__49452\,
            I => \N__48960\
        );

    \I__11714\ : SRMux
    port map (
            O => \N__49451\,
            I => \N__48960\
        );

    \I__11713\ : SRMux
    port map (
            O => \N__49450\,
            I => \N__48960\
        );

    \I__11712\ : Glb2LocalMux
    port map (
            O => \N__49447\,
            I => \N__48960\
        );

    \I__11711\ : SRMux
    port map (
            O => \N__49446\,
            I => \N__48960\
        );

    \I__11710\ : SRMux
    port map (
            O => \N__49445\,
            I => \N__48960\
        );

    \I__11709\ : SRMux
    port map (
            O => \N__49444\,
            I => \N__48960\
        );

    \I__11708\ : SRMux
    port map (
            O => \N__49443\,
            I => \N__48960\
        );

    \I__11707\ : SRMux
    port map (
            O => \N__49442\,
            I => \N__48960\
        );

    \I__11706\ : SRMux
    port map (
            O => \N__49441\,
            I => \N__48960\
        );

    \I__11705\ : SRMux
    port map (
            O => \N__49440\,
            I => \N__48960\
        );

    \I__11704\ : SRMux
    port map (
            O => \N__49439\,
            I => \N__48960\
        );

    \I__11703\ : SRMux
    port map (
            O => \N__49438\,
            I => \N__48960\
        );

    \I__11702\ : SRMux
    port map (
            O => \N__49437\,
            I => \N__48960\
        );

    \I__11701\ : SRMux
    port map (
            O => \N__49436\,
            I => \N__48960\
        );

    \I__11700\ : SRMux
    port map (
            O => \N__49435\,
            I => \N__48960\
        );

    \I__11699\ : SRMux
    port map (
            O => \N__49434\,
            I => \N__48960\
        );

    \I__11698\ : SRMux
    port map (
            O => \N__49433\,
            I => \N__48960\
        );

    \I__11697\ : SRMux
    port map (
            O => \N__49432\,
            I => \N__48960\
        );

    \I__11696\ : SRMux
    port map (
            O => \N__49431\,
            I => \N__48960\
        );

    \I__11695\ : SRMux
    port map (
            O => \N__49430\,
            I => \N__48960\
        );

    \I__11694\ : SRMux
    port map (
            O => \N__49429\,
            I => \N__48960\
        );

    \I__11693\ : SRMux
    port map (
            O => \N__49428\,
            I => \N__48960\
        );

    \I__11692\ : SRMux
    port map (
            O => \N__49427\,
            I => \N__48960\
        );

    \I__11691\ : SRMux
    port map (
            O => \N__49426\,
            I => \N__48960\
        );

    \I__11690\ : SRMux
    port map (
            O => \N__49425\,
            I => \N__48960\
        );

    \I__11689\ : SRMux
    port map (
            O => \N__49424\,
            I => \N__48960\
        );

    \I__11688\ : SRMux
    port map (
            O => \N__49423\,
            I => \N__48960\
        );

    \I__11687\ : SRMux
    port map (
            O => \N__49422\,
            I => \N__48960\
        );

    \I__11686\ : SRMux
    port map (
            O => \N__49421\,
            I => \N__48960\
        );

    \I__11685\ : SRMux
    port map (
            O => \N__49420\,
            I => \N__48960\
        );

    \I__11684\ : SRMux
    port map (
            O => \N__49419\,
            I => \N__48960\
        );

    \I__11683\ : SRMux
    port map (
            O => \N__49418\,
            I => \N__48960\
        );

    \I__11682\ : SRMux
    port map (
            O => \N__49417\,
            I => \N__48960\
        );

    \I__11681\ : SRMux
    port map (
            O => \N__49416\,
            I => \N__48960\
        );

    \I__11680\ : SRMux
    port map (
            O => \N__49415\,
            I => \N__48960\
        );

    \I__11679\ : SRMux
    port map (
            O => \N__49414\,
            I => \N__48960\
        );

    \I__11678\ : SRMux
    port map (
            O => \N__49413\,
            I => \N__48960\
        );

    \I__11677\ : SRMux
    port map (
            O => \N__49412\,
            I => \N__48960\
        );

    \I__11676\ : SRMux
    port map (
            O => \N__49411\,
            I => \N__48960\
        );

    \I__11675\ : SRMux
    port map (
            O => \N__49410\,
            I => \N__48960\
        );

    \I__11674\ : SRMux
    port map (
            O => \N__49409\,
            I => \N__48960\
        );

    \I__11673\ : SRMux
    port map (
            O => \N__49408\,
            I => \N__48960\
        );

    \I__11672\ : SRMux
    port map (
            O => \N__49407\,
            I => \N__48960\
        );

    \I__11671\ : SRMux
    port map (
            O => \N__49406\,
            I => \N__48960\
        );

    \I__11670\ : SRMux
    port map (
            O => \N__49405\,
            I => \N__48960\
        );

    \I__11669\ : SRMux
    port map (
            O => \N__49404\,
            I => \N__48960\
        );

    \I__11668\ : SRMux
    port map (
            O => \N__49403\,
            I => \N__48960\
        );

    \I__11667\ : SRMux
    port map (
            O => \N__49402\,
            I => \N__48960\
        );

    \I__11666\ : SRMux
    port map (
            O => \N__49401\,
            I => \N__48960\
        );

    \I__11665\ : SRMux
    port map (
            O => \N__49400\,
            I => \N__48960\
        );

    \I__11664\ : SRMux
    port map (
            O => \N__49399\,
            I => \N__48960\
        );

    \I__11663\ : SRMux
    port map (
            O => \N__49398\,
            I => \N__48960\
        );

    \I__11662\ : SRMux
    port map (
            O => \N__49397\,
            I => \N__48960\
        );

    \I__11661\ : SRMux
    port map (
            O => \N__49396\,
            I => \N__48960\
        );

    \I__11660\ : SRMux
    port map (
            O => \N__49395\,
            I => \N__48960\
        );

    \I__11659\ : SRMux
    port map (
            O => \N__49394\,
            I => \N__48960\
        );

    \I__11658\ : SRMux
    port map (
            O => \N__49393\,
            I => \N__48960\
        );

    \I__11657\ : SRMux
    port map (
            O => \N__49392\,
            I => \N__48960\
        );

    \I__11656\ : SRMux
    port map (
            O => \N__49391\,
            I => \N__48960\
        );

    \I__11655\ : SRMux
    port map (
            O => \N__49390\,
            I => \N__48960\
        );

    \I__11654\ : SRMux
    port map (
            O => \N__49389\,
            I => \N__48960\
        );

    \I__11653\ : SRMux
    port map (
            O => \N__49388\,
            I => \N__48960\
        );

    \I__11652\ : SRMux
    port map (
            O => \N__49387\,
            I => \N__48960\
        );

    \I__11651\ : SRMux
    port map (
            O => \N__49386\,
            I => \N__48960\
        );

    \I__11650\ : SRMux
    port map (
            O => \N__49385\,
            I => \N__48960\
        );

    \I__11649\ : SRMux
    port map (
            O => \N__49384\,
            I => \N__48960\
        );

    \I__11648\ : SRMux
    port map (
            O => \N__49383\,
            I => \N__48960\
        );

    \I__11647\ : SRMux
    port map (
            O => \N__49382\,
            I => \N__48960\
        );

    \I__11646\ : SRMux
    port map (
            O => \N__49381\,
            I => \N__48960\
        );

    \I__11645\ : SRMux
    port map (
            O => \N__49380\,
            I => \N__48960\
        );

    \I__11644\ : SRMux
    port map (
            O => \N__49379\,
            I => \N__48960\
        );

    \I__11643\ : SRMux
    port map (
            O => \N__49378\,
            I => \N__48960\
        );

    \I__11642\ : SRMux
    port map (
            O => \N__49377\,
            I => \N__48960\
        );

    \I__11641\ : SRMux
    port map (
            O => \N__49376\,
            I => \N__48960\
        );

    \I__11640\ : SRMux
    port map (
            O => \N__49375\,
            I => \N__48960\
        );

    \I__11639\ : SRMux
    port map (
            O => \N__49374\,
            I => \N__48960\
        );

    \I__11638\ : SRMux
    port map (
            O => \N__49373\,
            I => \N__48960\
        );

    \I__11637\ : SRMux
    port map (
            O => \N__49372\,
            I => \N__48960\
        );

    \I__11636\ : SRMux
    port map (
            O => \N__49371\,
            I => \N__48960\
        );

    \I__11635\ : SRMux
    port map (
            O => \N__49370\,
            I => \N__48960\
        );

    \I__11634\ : SRMux
    port map (
            O => \N__49369\,
            I => \N__48960\
        );

    \I__11633\ : SRMux
    port map (
            O => \N__49368\,
            I => \N__48960\
        );

    \I__11632\ : SRMux
    port map (
            O => \N__49367\,
            I => \N__48960\
        );

    \I__11631\ : SRMux
    port map (
            O => \N__49366\,
            I => \N__48960\
        );

    \I__11630\ : SRMux
    port map (
            O => \N__49365\,
            I => \N__48960\
        );

    \I__11629\ : SRMux
    port map (
            O => \N__49364\,
            I => \N__48960\
        );

    \I__11628\ : SRMux
    port map (
            O => \N__49363\,
            I => \N__48960\
        );

    \I__11627\ : SRMux
    port map (
            O => \N__49362\,
            I => \N__48960\
        );

    \I__11626\ : SRMux
    port map (
            O => \N__49361\,
            I => \N__48960\
        );

    \I__11625\ : SRMux
    port map (
            O => \N__49360\,
            I => \N__48960\
        );

    \I__11624\ : SRMux
    port map (
            O => \N__49359\,
            I => \N__48960\
        );

    \I__11623\ : SRMux
    port map (
            O => \N__49358\,
            I => \N__48960\
        );

    \I__11622\ : SRMux
    port map (
            O => \N__49357\,
            I => \N__48960\
        );

    \I__11621\ : SRMux
    port map (
            O => \N__49356\,
            I => \N__48960\
        );

    \I__11620\ : SRMux
    port map (
            O => \N__49355\,
            I => \N__48960\
        );

    \I__11619\ : SRMux
    port map (
            O => \N__49354\,
            I => \N__48960\
        );

    \I__11618\ : SRMux
    port map (
            O => \N__49353\,
            I => \N__48960\
        );

    \I__11617\ : SRMux
    port map (
            O => \N__49352\,
            I => \N__48960\
        );

    \I__11616\ : SRMux
    port map (
            O => \N__49351\,
            I => \N__48960\
        );

    \I__11615\ : SRMux
    port map (
            O => \N__49350\,
            I => \N__48960\
        );

    \I__11614\ : SRMux
    port map (
            O => \N__49349\,
            I => \N__48960\
        );

    \I__11613\ : SRMux
    port map (
            O => \N__49348\,
            I => \N__48960\
        );

    \I__11612\ : SRMux
    port map (
            O => \N__49347\,
            I => \N__48960\
        );

    \I__11611\ : SRMux
    port map (
            O => \N__49346\,
            I => \N__48960\
        );

    \I__11610\ : SRMux
    port map (
            O => \N__49345\,
            I => \N__48960\
        );

    \I__11609\ : SRMux
    port map (
            O => \N__49344\,
            I => \N__48960\
        );

    \I__11608\ : SRMux
    port map (
            O => \N__49343\,
            I => \N__48960\
        );

    \I__11607\ : SRMux
    port map (
            O => \N__49342\,
            I => \N__48960\
        );

    \I__11606\ : SRMux
    port map (
            O => \N__49341\,
            I => \N__48960\
        );

    \I__11605\ : SRMux
    port map (
            O => \N__49340\,
            I => \N__48960\
        );

    \I__11604\ : SRMux
    port map (
            O => \N__49339\,
            I => \N__48960\
        );

    \I__11603\ : SRMux
    port map (
            O => \N__49338\,
            I => \N__48960\
        );

    \I__11602\ : SRMux
    port map (
            O => \N__49337\,
            I => \N__48960\
        );

    \I__11601\ : SRMux
    port map (
            O => \N__49336\,
            I => \N__48960\
        );

    \I__11600\ : SRMux
    port map (
            O => \N__49335\,
            I => \N__48960\
        );

    \I__11599\ : SRMux
    port map (
            O => \N__49334\,
            I => \N__48960\
        );

    \I__11598\ : SRMux
    port map (
            O => \N__49333\,
            I => \N__48960\
        );

    \I__11597\ : SRMux
    port map (
            O => \N__49332\,
            I => \N__48960\
        );

    \I__11596\ : SRMux
    port map (
            O => \N__49331\,
            I => \N__48960\
        );

    \I__11595\ : SRMux
    port map (
            O => \N__49330\,
            I => \N__48960\
        );

    \I__11594\ : SRMux
    port map (
            O => \N__49329\,
            I => \N__48960\
        );

    \I__11593\ : SRMux
    port map (
            O => \N__49328\,
            I => \N__48960\
        );

    \I__11592\ : SRMux
    port map (
            O => \N__49327\,
            I => \N__48960\
        );

    \I__11591\ : SRMux
    port map (
            O => \N__49326\,
            I => \N__48960\
        );

    \I__11590\ : SRMux
    port map (
            O => \N__49325\,
            I => \N__48960\
        );

    \I__11589\ : SRMux
    port map (
            O => \N__49324\,
            I => \N__48960\
        );

    \I__11588\ : SRMux
    port map (
            O => \N__49323\,
            I => \N__48960\
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49322\,
            I => \N__48960\
        );

    \I__11586\ : SRMux
    port map (
            O => \N__49321\,
            I => \N__48960\
        );

    \I__11585\ : SRMux
    port map (
            O => \N__49320\,
            I => \N__48960\
        );

    \I__11584\ : SRMux
    port map (
            O => \N__49319\,
            I => \N__48960\
        );

    \I__11583\ : SRMux
    port map (
            O => \N__49318\,
            I => \N__48960\
        );

    \I__11582\ : SRMux
    port map (
            O => \N__49317\,
            I => \N__48960\
        );

    \I__11581\ : SRMux
    port map (
            O => \N__49316\,
            I => \N__48960\
        );

    \I__11580\ : SRMux
    port map (
            O => \N__49315\,
            I => \N__48960\
        );

    \I__11579\ : SRMux
    port map (
            O => \N__49314\,
            I => \N__48960\
        );

    \I__11578\ : SRMux
    port map (
            O => \N__49313\,
            I => \N__48960\
        );

    \I__11577\ : SRMux
    port map (
            O => \N__49312\,
            I => \N__48960\
        );

    \I__11576\ : SRMux
    port map (
            O => \N__49311\,
            I => \N__48960\
        );

    \I__11575\ : SRMux
    port map (
            O => \N__49310\,
            I => \N__48960\
        );

    \I__11574\ : SRMux
    port map (
            O => \N__49309\,
            I => \N__48960\
        );

    \I__11573\ : SRMux
    port map (
            O => \N__49308\,
            I => \N__48960\
        );

    \I__11572\ : SRMux
    port map (
            O => \N__49307\,
            I => \N__48960\
        );

    \I__11571\ : SRMux
    port map (
            O => \N__49306\,
            I => \N__48960\
        );

    \I__11570\ : SRMux
    port map (
            O => \N__49305\,
            I => \N__48960\
        );

    \I__11569\ : SRMux
    port map (
            O => \N__49304\,
            I => \N__48960\
        );

    \I__11568\ : SRMux
    port map (
            O => \N__49303\,
            I => \N__48960\
        );

    \I__11567\ : SRMux
    port map (
            O => \N__49302\,
            I => \N__48960\
        );

    \I__11566\ : SRMux
    port map (
            O => \N__49301\,
            I => \N__48960\
        );

    \I__11565\ : SRMux
    port map (
            O => \N__49300\,
            I => \N__48960\
        );

    \I__11564\ : SRMux
    port map (
            O => \N__49299\,
            I => \N__48960\
        );

    \I__11563\ : SRMux
    port map (
            O => \N__49298\,
            I => \N__48960\
        );

    \I__11562\ : SRMux
    port map (
            O => \N__49297\,
            I => \N__48960\
        );

    \I__11561\ : SRMux
    port map (
            O => \N__49296\,
            I => \N__48960\
        );

    \I__11560\ : SRMux
    port map (
            O => \N__49295\,
            I => \N__48960\
        );

    \I__11559\ : SRMux
    port map (
            O => \N__49294\,
            I => \N__48960\
        );

    \I__11558\ : SRMux
    port map (
            O => \N__49293\,
            I => \N__48960\
        );

    \I__11557\ : SRMux
    port map (
            O => \N__49292\,
            I => \N__48960\
        );

    \I__11556\ : SRMux
    port map (
            O => \N__49291\,
            I => \N__48960\
        );

    \I__11555\ : GlobalMux
    port map (
            O => \N__48960\,
            I => \N__48957\
        );

    \I__11554\ : gio2CtrlBuf
    port map (
            O => \N__48957\,
            I => red_c_g
        );

    \I__11553\ : InMux
    port map (
            O => \N__48954\,
            I => \N__48948\
        );

    \I__11552\ : CascadeMux
    port map (
            O => \N__48953\,
            I => \N__48945\
        );

    \I__11551\ : CascadeMux
    port map (
            O => \N__48952\,
            I => \N__48941\
        );

    \I__11550\ : CascadeMux
    port map (
            O => \N__48951\,
            I => \N__48937\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__48948\,
            I => \N__48933\
        );

    \I__11548\ : InMux
    port map (
            O => \N__48945\,
            I => \N__48919\
        );

    \I__11547\ : InMux
    port map (
            O => \N__48944\,
            I => \N__48919\
        );

    \I__11546\ : InMux
    port map (
            O => \N__48941\,
            I => \N__48919\
        );

    \I__11545\ : InMux
    port map (
            O => \N__48940\,
            I => \N__48919\
        );

    \I__11544\ : InMux
    port map (
            O => \N__48937\,
            I => \N__48919\
        );

    \I__11543\ : InMux
    port map (
            O => \N__48936\,
            I => \N__48919\
        );

    \I__11542\ : Span12Mux_s7_v
    port map (
            O => \N__48933\,
            I => \N__48916\
        );

    \I__11541\ : InMux
    port map (
            O => \N__48932\,
            I => \N__48913\
        );

    \I__11540\ : LocalMux
    port map (
            O => \N__48919\,
            I => \N__48910\
        );

    \I__11539\ : Span12Mux_h
    port map (
            O => \N__48916\,
            I => \N__48905\
        );

    \I__11538\ : LocalMux
    port map (
            O => \N__48913\,
            I => \N__48905\
        );

    \I__11537\ : Span4Mux_h
    port map (
            O => \N__48910\,
            I => \N__48902\
        );

    \I__11536\ : Span12Mux_h
    port map (
            O => \N__48905\,
            I => \N__48899\
        );

    \I__11535\ : Span4Mux_h
    port map (
            O => \N__48902\,
            I => \N__48896\
        );

    \I__11534\ : Odrv12
    port map (
            O => \N__48899\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__11533\ : Odrv4
    port map (
            O => \N__48896\,
            I => \pwm_generator_inst.un2_threshold_1_25\
        );

    \I__11532\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48888\
        );

    \I__11531\ : LocalMux
    port map (
            O => \N__48888\,
            I => \N__48885\
        );

    \I__11530\ : Span12Mux_v
    port map (
            O => \N__48885\,
            I => \N__48882\
        );

    \I__11529\ : Span12Mux_h
    port map (
            O => \N__48882\,
            I => \N__48878\
        );

    \I__11528\ : InMux
    port map (
            O => \N__48881\,
            I => \N__48875\
        );

    \I__11527\ : Odrv12
    port map (
            O => \N__48878\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__48875\,
            I => \pwm_generator_inst.un2_threshold_2_1_15\
        );

    \I__11525\ : CascadeMux
    port map (
            O => \N__48870\,
            I => \N__48846\
        );

    \I__11524\ : CascadeMux
    port map (
            O => \N__48869\,
            I => \N__48843\
        );

    \I__11523\ : InMux
    port map (
            O => \N__48868\,
            I => \N__48840\
        );

    \I__11522\ : InMux
    port map (
            O => \N__48867\,
            I => \N__48818\
        );

    \I__11521\ : InMux
    port map (
            O => \N__48866\,
            I => \N__48818\
        );

    \I__11520\ : InMux
    port map (
            O => \N__48865\,
            I => \N__48818\
        );

    \I__11519\ : InMux
    port map (
            O => \N__48864\,
            I => \N__48818\
        );

    \I__11518\ : InMux
    port map (
            O => \N__48863\,
            I => \N__48818\
        );

    \I__11517\ : InMux
    port map (
            O => \N__48862\,
            I => \N__48818\
        );

    \I__11516\ : InMux
    port map (
            O => \N__48861\,
            I => \N__48818\
        );

    \I__11515\ : InMux
    port map (
            O => \N__48860\,
            I => \N__48818\
        );

    \I__11514\ : InMux
    port map (
            O => \N__48859\,
            I => \N__48803\
        );

    \I__11513\ : InMux
    port map (
            O => \N__48858\,
            I => \N__48803\
        );

    \I__11512\ : InMux
    port map (
            O => \N__48857\,
            I => \N__48803\
        );

    \I__11511\ : InMux
    port map (
            O => \N__48856\,
            I => \N__48803\
        );

    \I__11510\ : InMux
    port map (
            O => \N__48855\,
            I => \N__48803\
        );

    \I__11509\ : InMux
    port map (
            O => \N__48854\,
            I => \N__48803\
        );

    \I__11508\ : InMux
    port map (
            O => \N__48853\,
            I => \N__48803\
        );

    \I__11507\ : CascadeMux
    port map (
            O => \N__48852\,
            I => \N__48800\
        );

    \I__11506\ : CascadeMux
    port map (
            O => \N__48851\,
            I => \N__48797\
        );

    \I__11505\ : CascadeMux
    port map (
            O => \N__48850\,
            I => \N__48793\
        );

    \I__11504\ : CascadeMux
    port map (
            O => \N__48849\,
            I => \N__48790\
        );

    \I__11503\ : InMux
    port map (
            O => \N__48846\,
            I => \N__48785\
        );

    \I__11502\ : InMux
    port map (
            O => \N__48843\,
            I => \N__48785\
        );

    \I__11501\ : LocalMux
    port map (
            O => \N__48840\,
            I => \N__48782\
        );

    \I__11500\ : InMux
    port map (
            O => \N__48839\,
            I => \N__48775\
        );

    \I__11499\ : InMux
    port map (
            O => \N__48838\,
            I => \N__48775\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48837\,
            I => \N__48768\
        );

    \I__11497\ : InMux
    port map (
            O => \N__48836\,
            I => \N__48768\
        );

    \I__11496\ : InMux
    port map (
            O => \N__48835\,
            I => \N__48768\
        );

    \I__11495\ : LocalMux
    port map (
            O => \N__48818\,
            I => \N__48763\
        );

    \I__11494\ : LocalMux
    port map (
            O => \N__48803\,
            I => \N__48763\
        );

    \I__11493\ : InMux
    port map (
            O => \N__48800\,
            I => \N__48758\
        );

    \I__11492\ : InMux
    port map (
            O => \N__48797\,
            I => \N__48758\
        );

    \I__11491\ : InMux
    port map (
            O => \N__48796\,
            I => \N__48751\
        );

    \I__11490\ : InMux
    port map (
            O => \N__48793\,
            I => \N__48751\
        );

    \I__11489\ : InMux
    port map (
            O => \N__48790\,
            I => \N__48751\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__48785\,
            I => \N__48748\
        );

    \I__11487\ : Span4Mux_s3_h
    port map (
            O => \N__48782\,
            I => \N__48745\
        );

    \I__11486\ : CascadeMux
    port map (
            O => \N__48781\,
            I => \N__48742\
        );

    \I__11485\ : InMux
    port map (
            O => \N__48780\,
            I => \N__48739\
        );

    \I__11484\ : LocalMux
    port map (
            O => \N__48775\,
            I => \N__48734\
        );

    \I__11483\ : LocalMux
    port map (
            O => \N__48768\,
            I => \N__48734\
        );

    \I__11482\ : Span4Mux_s3_h
    port map (
            O => \N__48763\,
            I => \N__48731\
        );

    \I__11481\ : LocalMux
    port map (
            O => \N__48758\,
            I => \N__48722\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__48751\,
            I => \N__48722\
        );

    \I__11479\ : Span4Mux_h
    port map (
            O => \N__48748\,
            I => \N__48722\
        );

    \I__11478\ : Span4Mux_h
    port map (
            O => \N__48745\,
            I => \N__48719\
        );

    \I__11477\ : InMux
    port map (
            O => \N__48742\,
            I => \N__48716\
        );

    \I__11476\ : LocalMux
    port map (
            O => \N__48739\,
            I => \N__48713\
        );

    \I__11475\ : Span4Mux_s2_h
    port map (
            O => \N__48734\,
            I => \N__48710\
        );

    \I__11474\ : Span4Mux_h
    port map (
            O => \N__48731\,
            I => \N__48707\
        );

    \I__11473\ : CascadeMux
    port map (
            O => \N__48730\,
            I => \N__48704\
        );

    \I__11472\ : CascadeMux
    port map (
            O => \N__48729\,
            I => \N__48701\
        );

    \I__11471\ : Span4Mux_h
    port map (
            O => \N__48722\,
            I => \N__48696\
        );

    \I__11470\ : Span4Mux_h
    port map (
            O => \N__48719\,
            I => \N__48696\
        );

    \I__11469\ : LocalMux
    port map (
            O => \N__48716\,
            I => \N__48689\
        );

    \I__11468\ : Span4Mux_h
    port map (
            O => \N__48713\,
            I => \N__48689\
        );

    \I__11467\ : Span4Mux_h
    port map (
            O => \N__48710\,
            I => \N__48689\
        );

    \I__11466\ : Span4Mux_h
    port map (
            O => \N__48707\,
            I => \N__48686\
        );

    \I__11465\ : InMux
    port map (
            O => \N__48704\,
            I => \N__48683\
        );

    \I__11464\ : InMux
    port map (
            O => \N__48701\,
            I => \N__48680\
        );

    \I__11463\ : Span4Mux_h
    port map (
            O => \N__48696\,
            I => \N__48677\
        );

    \I__11462\ : Span4Mux_h
    port map (
            O => \N__48689\,
            I => \N__48672\
        );

    \I__11461\ : Span4Mux_h
    port map (
            O => \N__48686\,
            I => \N__48672\
        );

    \I__11460\ : LocalMux
    port map (
            O => \N__48683\,
            I => \N_19_1\
        );

    \I__11459\ : LocalMux
    port map (
            O => \N__48680\,
            I => \N_19_1\
        );

    \I__11458\ : Odrv4
    port map (
            O => \N__48677\,
            I => \N_19_1\
        );

    \I__11457\ : Odrv4
    port map (
            O => \N__48672\,
            I => \N_19_1\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48663\,
            I => \N__48660\
        );

    \I__11455\ : LocalMux
    port map (
            O => \N__48660\,
            I => \N__48657\
        );

    \I__11454\ : Span12Mux_s8_h
    port map (
            O => \N__48657\,
            I => \N__48654\
        );

    \I__11453\ : Span12Mux_h
    port map (
            O => \N__48654\,
            I => \N__48651\
        );

    \I__11452\ : Odrv12
    port map (
            O => \N__48651\,
            I => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\
        );

    \I__11451\ : InMux
    port map (
            O => \N__48648\,
            I => \N__48629\
        );

    \I__11450\ : InMux
    port map (
            O => \N__48647\,
            I => \N__48629\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48646\,
            I => \N__48629\
        );

    \I__11448\ : InMux
    port map (
            O => \N__48645\,
            I => \N__48629\
        );

    \I__11447\ : InMux
    port map (
            O => \N__48644\,
            I => \N__48619\
        );

    \I__11446\ : InMux
    port map (
            O => \N__48643\,
            I => \N__48612\
        );

    \I__11445\ : InMux
    port map (
            O => \N__48642\,
            I => \N__48612\
        );

    \I__11444\ : InMux
    port map (
            O => \N__48641\,
            I => \N__48612\
        );

    \I__11443\ : InMux
    port map (
            O => \N__48640\,
            I => \N__48607\
        );

    \I__11442\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48607\
        );

    \I__11441\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48604\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48629\,
            I => \N__48601\
        );

    \I__11439\ : InMux
    port map (
            O => \N__48628\,
            I => \N__48592\
        );

    \I__11438\ : InMux
    port map (
            O => \N__48627\,
            I => \N__48592\
        );

    \I__11437\ : InMux
    port map (
            O => \N__48626\,
            I => \N__48592\
        );

    \I__11436\ : InMux
    port map (
            O => \N__48625\,
            I => \N__48592\
        );

    \I__11435\ : InMux
    port map (
            O => \N__48624\,
            I => \N__48585\
        );

    \I__11434\ : InMux
    port map (
            O => \N__48623\,
            I => \N__48585\
        );

    \I__11433\ : InMux
    port map (
            O => \N__48622\,
            I => \N__48585\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__48619\,
            I => \N__48577\
        );

    \I__11431\ : LocalMux
    port map (
            O => \N__48612\,
            I => \N__48574\
        );

    \I__11430\ : LocalMux
    port map (
            O => \N__48607\,
            I => \N__48563\
        );

    \I__11429\ : LocalMux
    port map (
            O => \N__48604\,
            I => \N__48563\
        );

    \I__11428\ : Span4Mux_v
    port map (
            O => \N__48601\,
            I => \N__48563\
        );

    \I__11427\ : LocalMux
    port map (
            O => \N__48592\,
            I => \N__48563\
        );

    \I__11426\ : LocalMux
    port map (
            O => \N__48585\,
            I => \N__48563\
        );

    \I__11425\ : InMux
    port map (
            O => \N__48584\,
            I => \N__48552\
        );

    \I__11424\ : InMux
    port map (
            O => \N__48583\,
            I => \N__48552\
        );

    \I__11423\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48552\
        );

    \I__11422\ : InMux
    port map (
            O => \N__48581\,
            I => \N__48552\
        );

    \I__11421\ : InMux
    port map (
            O => \N__48580\,
            I => \N__48552\
        );

    \I__11420\ : Span4Mux_h
    port map (
            O => \N__48577\,
            I => \N__48545\
        );

    \I__11419\ : Span4Mux_v
    port map (
            O => \N__48574\,
            I => \N__48545\
        );

    \I__11418\ : Span4Mux_v
    port map (
            O => \N__48563\,
            I => \N__48540\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48552\,
            I => \N__48540\
        );

    \I__11416\ : InMux
    port map (
            O => \N__48551\,
            I => \N__48537\
        );

    \I__11415\ : InMux
    port map (
            O => \N__48550\,
            I => \N__48534\
        );

    \I__11414\ : Odrv4
    port map (
            O => \N__48545\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11413\ : Odrv4
    port map (
            O => \N__48540\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48537\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__48534\,
            I => \current_shift_inst.elapsed_time_ns_s1_31_rep1\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48525\,
            I => \N__48520\
        );

    \I__11409\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48517\
        );

    \I__11408\ : InMux
    port map (
            O => \N__48523\,
            I => \N__48514\
        );

    \I__11407\ : LocalMux
    port map (
            O => \N__48520\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__48517\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__11405\ : LocalMux
    port map (
            O => \N__48514\,
            I => \current_shift_inst.un4_control_input1_2\
        );

    \I__11404\ : InMux
    port map (
            O => \N__48507\,
            I => \N__48504\
        );

    \I__11403\ : LocalMux
    port map (
            O => \N__48504\,
            I => \N__48498\
        );

    \I__11402\ : InMux
    port map (
            O => \N__48503\,
            I => \N__48491\
        );

    \I__11401\ : InMux
    port map (
            O => \N__48502\,
            I => \N__48491\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48501\,
            I => \N__48491\
        );

    \I__11399\ : Odrv4
    port map (
            O => \N__48498\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48491\,
            I => \current_shift_inst.elapsed_time_ns_s1_2\
        );

    \I__11397\ : CascadeMux
    port map (
            O => \N__48486\,
            I => \N__48483\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48480\
        );

    \I__11395\ : LocalMux
    port map (
            O => \N__48480\,
            I => \N__48477\
        );

    \I__11394\ : Span4Mux_v
    port map (
            O => \N__48477\,
            I => \N__48474\
        );

    \I__11393\ : Span4Mux_h
    port map (
            O => \N__48474\,
            I => \N__48471\
        );

    \I__11392\ : Odrv4
    port map (
            O => \N__48471\,
            I => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\
        );

    \I__11391\ : InMux
    port map (
            O => \N__48468\,
            I => \N__48464\
        );

    \I__11390\ : InMux
    port map (
            O => \N__48467\,
            I => \N__48461\
        );

    \I__11389\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48457\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__48461\,
            I => \N__48454\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48460\,
            I => \N__48451\
        );

    \I__11386\ : Span4Mux_h
    port map (
            O => \N__48457\,
            I => \N__48447\
        );

    \I__11385\ : Span4Mux_v
    port map (
            O => \N__48454\,
            I => \N__48442\
        );

    \I__11384\ : LocalMux
    port map (
            O => \N__48451\,
            I => \N__48442\
        );

    \I__11383\ : InMux
    port map (
            O => \N__48450\,
            I => \N__48439\
        );

    \I__11382\ : Odrv4
    port map (
            O => \N__48447\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__11381\ : Odrv4
    port map (
            O => \N__48442\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__48439\,
            I => \current_shift_inst.elapsed_time_ns_s1_13\
        );

    \I__11379\ : CascadeMux
    port map (
            O => \N__48432\,
            I => \N__48429\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48429\,
            I => \N__48426\
        );

    \I__11377\ : LocalMux
    port map (
            O => \N__48426\,
            I => \N__48422\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48425\,
            I => \N__48418\
        );

    \I__11375\ : Span4Mux_v
    port map (
            O => \N__48422\,
            I => \N__48415\
        );

    \I__11374\ : InMux
    port map (
            O => \N__48421\,
            I => \N__48412\
        );

    \I__11373\ : LocalMux
    port map (
            O => \N__48418\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__11372\ : Odrv4
    port map (
            O => \N__48415\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__11371\ : LocalMux
    port map (
            O => \N__48412\,
            I => \current_shift_inst.un4_control_input1_13\
        );

    \I__11370\ : CascadeMux
    port map (
            O => \N__48405\,
            I => \N__48402\
        );

    \I__11369\ : InMux
    port map (
            O => \N__48402\,
            I => \N__48399\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__48399\,
            I => \N__48396\
        );

    \I__11367\ : Odrv12
    port map (
            O => \N__48396\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\
        );

    \I__11366\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48389\
        );

    \I__11365\ : InMux
    port map (
            O => \N__48392\,
            I => \N__48386\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__48389\,
            I => \N__48381\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__48386\,
            I => \N__48378\
        );

    \I__11362\ : InMux
    port map (
            O => \N__48385\,
            I => \N__48373\
        );

    \I__11361\ : InMux
    port map (
            O => \N__48384\,
            I => \N__48373\
        );

    \I__11360\ : Span4Mux_v
    port map (
            O => \N__48381\,
            I => \N__48368\
        );

    \I__11359\ : Span4Mux_h
    port map (
            O => \N__48378\,
            I => \N__48368\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__48373\,
            I => \N__48365\
        );

    \I__11357\ : Odrv4
    port map (
            O => \N__48368\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__11356\ : Odrv4
    port map (
            O => \N__48365\,
            I => \current_shift_inst.elapsed_time_ns_s1_11\
        );

    \I__11355\ : InMux
    port map (
            O => \N__48360\,
            I => \N__48357\
        );

    \I__11354\ : LocalMux
    port map (
            O => \N__48357\,
            I => \N__48354\
        );

    \I__11353\ : Span4Mux_h
    port map (
            O => \N__48354\,
            I => \N__48349\
        );

    \I__11352\ : InMux
    port map (
            O => \N__48353\,
            I => \N__48346\
        );

    \I__11351\ : InMux
    port map (
            O => \N__48352\,
            I => \N__48343\
        );

    \I__11350\ : Odrv4
    port map (
            O => \N__48349\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__48346\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__48343\,
            I => \current_shift_inst.un4_control_input1_11\
        );

    \I__11347\ : CascadeMux
    port map (
            O => \N__48336\,
            I => \N__48333\
        );

    \I__11346\ : InMux
    port map (
            O => \N__48333\,
            I => \N__48330\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__48330\,
            I => \N__48327\
        );

    \I__11344\ : Span4Mux_h
    port map (
            O => \N__48327\,
            I => \N__48324\
        );

    \I__11343\ : Odrv4
    port map (
            O => \N__48324\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\
        );

    \I__11342\ : CascadeMux
    port map (
            O => \N__48321\,
            I => \N__48318\
        );

    \I__11341\ : InMux
    port map (
            O => \N__48318\,
            I => \N__48315\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__48315\,
            I => \N__48310\
        );

    \I__11339\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48305\
        );

    \I__11338\ : InMux
    port map (
            O => \N__48313\,
            I => \N__48305\
        );

    \I__11337\ : Span4Mux_h
    port map (
            O => \N__48310\,
            I => \N__48299\
        );

    \I__11336\ : LocalMux
    port map (
            O => \N__48305\,
            I => \N__48299\
        );

    \I__11335\ : InMux
    port map (
            O => \N__48304\,
            I => \N__48296\
        );

    \I__11334\ : Odrv4
    port map (
            O => \N__48299\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11333\ : LocalMux
    port map (
            O => \N__48296\,
            I => \current_shift_inst.elapsed_time_ns_s1_21\
        );

    \I__11332\ : CascadeMux
    port map (
            O => \N__48291\,
            I => \N__48288\
        );

    \I__11331\ : InMux
    port map (
            O => \N__48288\,
            I => \N__48283\
        );

    \I__11330\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48280\
        );

    \I__11329\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48277\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__48283\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__11327\ : LocalMux
    port map (
            O => \N__48280\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__11326\ : LocalMux
    port map (
            O => \N__48277\,
            I => \current_shift_inst.un4_control_input1_21\
        );

    \I__11325\ : CascadeMux
    port map (
            O => \N__48270\,
            I => \N__48267\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48267\,
            I => \N__48264\
        );

    \I__11323\ : LocalMux
    port map (
            O => \N__48264\,
            I => \N__48261\
        );

    \I__11322\ : Span4Mux_h
    port map (
            O => \N__48261\,
            I => \N__48258\
        );

    \I__11321\ : Odrv4
    port map (
            O => \N__48258\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\
        );

    \I__11320\ : InMux
    port map (
            O => \N__48255\,
            I => \N__48248\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48254\,
            I => \N__48245\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48253\,
            I => \N__48229\
        );

    \I__11317\ : InMux
    port map (
            O => \N__48252\,
            I => \N__48229\
        );

    \I__11316\ : CascadeMux
    port map (
            O => \N__48251\,
            I => \N__48217\
        );

    \I__11315\ : LocalMux
    port map (
            O => \N__48248\,
            I => \N__48202\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__48245\,
            I => \N__48199\
        );

    \I__11313\ : InMux
    port map (
            O => \N__48244\,
            I => \N__48191\
        );

    \I__11312\ : InMux
    port map (
            O => \N__48243\,
            I => \N__48191\
        );

    \I__11311\ : InMux
    port map (
            O => \N__48242\,
            I => \N__48188\
        );

    \I__11310\ : InMux
    port map (
            O => \N__48241\,
            I => \N__48170\
        );

    \I__11309\ : InMux
    port map (
            O => \N__48240\,
            I => \N__48170\
        );

    \I__11308\ : InMux
    port map (
            O => \N__48239\,
            I => \N__48170\
        );

    \I__11307\ : InMux
    port map (
            O => \N__48238\,
            I => \N__48170\
        );

    \I__11306\ : InMux
    port map (
            O => \N__48237\,
            I => \N__48159\
        );

    \I__11305\ : InMux
    port map (
            O => \N__48236\,
            I => \N__48159\
        );

    \I__11304\ : InMux
    port map (
            O => \N__48235\,
            I => \N__48154\
        );

    \I__11303\ : InMux
    port map (
            O => \N__48234\,
            I => \N__48154\
        );

    \I__11302\ : LocalMux
    port map (
            O => \N__48229\,
            I => \N__48151\
        );

    \I__11301\ : InMux
    port map (
            O => \N__48228\,
            I => \N__48142\
        );

    \I__11300\ : InMux
    port map (
            O => \N__48227\,
            I => \N__48142\
        );

    \I__11299\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48142\
        );

    \I__11298\ : InMux
    port map (
            O => \N__48225\,
            I => \N__48142\
        );

    \I__11297\ : InMux
    port map (
            O => \N__48224\,
            I => \N__48127\
        );

    \I__11296\ : InMux
    port map (
            O => \N__48223\,
            I => \N__48127\
        );

    \I__11295\ : InMux
    port map (
            O => \N__48222\,
            I => \N__48127\
        );

    \I__11294\ : InMux
    port map (
            O => \N__48221\,
            I => \N__48127\
        );

    \I__11293\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48127\
        );

    \I__11292\ : InMux
    port map (
            O => \N__48217\,
            I => \N__48127\
        );

    \I__11291\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48127\
        );

    \I__11290\ : InMux
    port map (
            O => \N__48215\,
            I => \N__48110\
        );

    \I__11289\ : InMux
    port map (
            O => \N__48214\,
            I => \N__48110\
        );

    \I__11288\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48110\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48212\,
            I => \N__48110\
        );

    \I__11286\ : InMux
    port map (
            O => \N__48211\,
            I => \N__48110\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48210\,
            I => \N__48110\
        );

    \I__11284\ : InMux
    port map (
            O => \N__48209\,
            I => \N__48110\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48208\,
            I => \N__48110\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48207\,
            I => \N__48107\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48206\,
            I => \N__48104\
        );

    \I__11280\ : InMux
    port map (
            O => \N__48205\,
            I => \N__48101\
        );

    \I__11279\ : Span4Mux_v
    port map (
            O => \N__48202\,
            I => \N__48098\
        );

    \I__11278\ : Span4Mux_v
    port map (
            O => \N__48199\,
            I => \N__48095\
        );

    \I__11277\ : CascadeMux
    port map (
            O => \N__48198\,
            I => \N__48088\
        );

    \I__11276\ : InMux
    port map (
            O => \N__48197\,
            I => \N__48074\
        );

    \I__11275\ : InMux
    port map (
            O => \N__48196\,
            I => \N__48074\
        );

    \I__11274\ : LocalMux
    port map (
            O => \N__48191\,
            I => \N__48071\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__48188\,
            I => \N__48068\
        );

    \I__11272\ : InMux
    port map (
            O => \N__48187\,
            I => \N__48061\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48186\,
            I => \N__48061\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48061\
        );

    \I__11269\ : InMux
    port map (
            O => \N__48184\,
            I => \N__48056\
        );

    \I__11268\ : InMux
    port map (
            O => \N__48183\,
            I => \N__48056\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48182\,
            I => \N__48047\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48047\
        );

    \I__11265\ : InMux
    port map (
            O => \N__48180\,
            I => \N__48047\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48179\,
            I => \N__48047\
        );

    \I__11263\ : LocalMux
    port map (
            O => \N__48170\,
            I => \N__48044\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48169\,
            I => \N__48031\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48168\,
            I => \N__48031\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48167\,
            I => \N__48031\
        );

    \I__11259\ : InMux
    port map (
            O => \N__48166\,
            I => \N__48031\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48165\,
            I => \N__48031\
        );

    \I__11257\ : InMux
    port map (
            O => \N__48164\,
            I => \N__48031\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__48159\,
            I => \N__48016\
        );

    \I__11255\ : LocalMux
    port map (
            O => \N__48154\,
            I => \N__48016\
        );

    \I__11254\ : Span4Mux_v
    port map (
            O => \N__48151\,
            I => \N__48016\
        );

    \I__11253\ : LocalMux
    port map (
            O => \N__48142\,
            I => \N__48016\
        );

    \I__11252\ : LocalMux
    port map (
            O => \N__48127\,
            I => \N__48016\
        );

    \I__11251\ : LocalMux
    port map (
            O => \N__48110\,
            I => \N__48016\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__48107\,
            I => \N__48016\
        );

    \I__11249\ : LocalMux
    port map (
            O => \N__48104\,
            I => \N__48011\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__48101\,
            I => \N__48011\
        );

    \I__11247\ : Span4Mux_h
    port map (
            O => \N__48098\,
            I => \N__48003\
        );

    \I__11246\ : Span4Mux_h
    port map (
            O => \N__48095\,
            I => \N__48003\
        );

    \I__11245\ : InMux
    port map (
            O => \N__48094\,
            I => \N__47998\
        );

    \I__11244\ : InMux
    port map (
            O => \N__48093\,
            I => \N__47998\
        );

    \I__11243\ : InMux
    port map (
            O => \N__48092\,
            I => \N__47995\
        );

    \I__11242\ : InMux
    port map (
            O => \N__48091\,
            I => \N__47990\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48088\,
            I => \N__47990\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48087\,
            I => \N__47987\
        );

    \I__11239\ : InMux
    port map (
            O => \N__48086\,
            I => \N__47984\
        );

    \I__11238\ : InMux
    port map (
            O => \N__48085\,
            I => \N__47969\
        );

    \I__11237\ : InMux
    port map (
            O => \N__48084\,
            I => \N__47969\
        );

    \I__11236\ : InMux
    port map (
            O => \N__48083\,
            I => \N__47969\
        );

    \I__11235\ : InMux
    port map (
            O => \N__48082\,
            I => \N__47969\
        );

    \I__11234\ : InMux
    port map (
            O => \N__48081\,
            I => \N__47969\
        );

    \I__11233\ : InMux
    port map (
            O => \N__48080\,
            I => \N__47969\
        );

    \I__11232\ : InMux
    port map (
            O => \N__48079\,
            I => \N__47969\
        );

    \I__11231\ : LocalMux
    port map (
            O => \N__48074\,
            I => \N__47956\
        );

    \I__11230\ : Sp12to4
    port map (
            O => \N__48071\,
            I => \N__47956\
        );

    \I__11229\ : Sp12to4
    port map (
            O => \N__48068\,
            I => \N__47956\
        );

    \I__11228\ : LocalMux
    port map (
            O => \N__48061\,
            I => \N__47956\
        );

    \I__11227\ : LocalMux
    port map (
            O => \N__48056\,
            I => \N__47956\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__48047\,
            I => \N__47956\
        );

    \I__11225\ : Span4Mux_v
    port map (
            O => \N__48044\,
            I => \N__47947\
        );

    \I__11224\ : LocalMux
    port map (
            O => \N__48031\,
            I => \N__47947\
        );

    \I__11223\ : Span4Mux_v
    port map (
            O => \N__48016\,
            I => \N__47947\
        );

    \I__11222\ : Span4Mux_v
    port map (
            O => \N__48011\,
            I => \N__47947\
        );

    \I__11221\ : InMux
    port map (
            O => \N__48010\,
            I => \N__47940\
        );

    \I__11220\ : InMux
    port map (
            O => \N__48009\,
            I => \N__47940\
        );

    \I__11219\ : InMux
    port map (
            O => \N__48008\,
            I => \N__47940\
        );

    \I__11218\ : Odrv4
    port map (
            O => \N__48003\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11217\ : LocalMux
    port map (
            O => \N__47998\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11216\ : LocalMux
    port map (
            O => \N__47995\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11215\ : LocalMux
    port map (
            O => \N__47990\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__47987\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__47984\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11212\ : LocalMux
    port map (
            O => \N__47969\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11211\ : Odrv12
    port map (
            O => \N__47956\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11210\ : Odrv4
    port map (
            O => \N__47947\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__47940\,
            I => \current_shift_inst.elapsed_time_ns_s1_31\
        );

    \I__11208\ : InMux
    port map (
            O => \N__47919\,
            I => \N__47915\
        );

    \I__11207\ : CascadeMux
    port map (
            O => \N__47918\,
            I => \N__47912\
        );

    \I__11206\ : LocalMux
    port map (
            O => \N__47915\,
            I => \N__47908\
        );

    \I__11205\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47905\
        );

    \I__11204\ : InMux
    port map (
            O => \N__47911\,
            I => \N__47902\
        );

    \I__11203\ : Span4Mux_h
    port map (
            O => \N__47908\,
            I => \N__47898\
        );

    \I__11202\ : LocalMux
    port map (
            O => \N__47905\,
            I => \N__47895\
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__47902\,
            I => \N__47892\
        );

    \I__11200\ : InMux
    port map (
            O => \N__47901\,
            I => \N__47889\
        );

    \I__11199\ : Odrv4
    port map (
            O => \N__47898\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__11198\ : Odrv12
    port map (
            O => \N__47895\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__11197\ : Odrv4
    port map (
            O => \N__47892\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__11196\ : LocalMux
    port map (
            O => \N__47889\,
            I => \current_shift_inst.elapsed_time_ns_s1_14\
        );

    \I__11195\ : CascadeMux
    port map (
            O => \N__47880\,
            I => \N__47867\
        );

    \I__11194\ : CascadeMux
    port map (
            O => \N__47879\,
            I => \N__47858\
        );

    \I__11193\ : CascadeMux
    port map (
            O => \N__47878\,
            I => \N__47854\
        );

    \I__11192\ : CascadeMux
    port map (
            O => \N__47877\,
            I => \N__47850\
        );

    \I__11191\ : CascadeMux
    port map (
            O => \N__47876\,
            I => \N__47843\
        );

    \I__11190\ : CascadeMux
    port map (
            O => \N__47875\,
            I => \N__47840\
        );

    \I__11189\ : CascadeMux
    port map (
            O => \N__47874\,
            I => \N__47831\
        );

    \I__11188\ : CascadeMux
    port map (
            O => \N__47873\,
            I => \N__47827\
        );

    \I__11187\ : CascadeMux
    port map (
            O => \N__47872\,
            I => \N__47823\
        );

    \I__11186\ : InMux
    port map (
            O => \N__47871\,
            I => \N__47802\
        );

    \I__11185\ : InMux
    port map (
            O => \N__47870\,
            I => \N__47802\
        );

    \I__11184\ : InMux
    port map (
            O => \N__47867\,
            I => \N__47792\
        );

    \I__11183\ : CascadeMux
    port map (
            O => \N__47866\,
            I => \N__47788\
        );

    \I__11182\ : CascadeMux
    port map (
            O => \N__47865\,
            I => \N__47785\
        );

    \I__11181\ : CascadeMux
    port map (
            O => \N__47864\,
            I => \N__47782\
        );

    \I__11180\ : InMux
    port map (
            O => \N__47863\,
            I => \N__47769\
        );

    \I__11179\ : InMux
    port map (
            O => \N__47862\,
            I => \N__47769\
        );

    \I__11178\ : InMux
    port map (
            O => \N__47861\,
            I => \N__47769\
        );

    \I__11177\ : InMux
    port map (
            O => \N__47858\,
            I => \N__47769\
        );

    \I__11176\ : InMux
    port map (
            O => \N__47857\,
            I => \N__47769\
        );

    \I__11175\ : InMux
    port map (
            O => \N__47854\,
            I => \N__47769\
        );

    \I__11174\ : InMux
    port map (
            O => \N__47853\,
            I => \N__47763\
        );

    \I__11173\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47763\
        );

    \I__11172\ : InMux
    port map (
            O => \N__47849\,
            I => \N__47758\
        );

    \I__11171\ : InMux
    port map (
            O => \N__47848\,
            I => \N__47758\
        );

    \I__11170\ : CascadeMux
    port map (
            O => \N__47847\,
            I => \N__47751\
        );

    \I__11169\ : CascadeMux
    port map (
            O => \N__47846\,
            I => \N__47747\
        );

    \I__11168\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47736\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47840\,
            I => \N__47733\
        );

    \I__11166\ : CascadeMux
    port map (
            O => \N__47839\,
            I => \N__47730\
        );

    \I__11165\ : CascadeMux
    port map (
            O => \N__47838\,
            I => \N__47726\
        );

    \I__11164\ : CascadeMux
    port map (
            O => \N__47837\,
            I => \N__47722\
        );

    \I__11163\ : CascadeMux
    port map (
            O => \N__47836\,
            I => \N__47718\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47835\,
            I => \N__47701\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47834\,
            I => \N__47701\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47701\
        );

    \I__11159\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47701\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47827\,
            I => \N__47701\
        );

    \I__11157\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47701\
        );

    \I__11156\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47701\
        );

    \I__11155\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47701\
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__47821\,
            I => \N__47698\
        );

    \I__11153\ : CascadeMux
    port map (
            O => \N__47820\,
            I => \N__47694\
        );

    \I__11152\ : CascadeMux
    port map (
            O => \N__47819\,
            I => \N__47690\
        );

    \I__11151\ : CascadeMux
    port map (
            O => \N__47818\,
            I => \N__47686\
        );

    \I__11150\ : CascadeMux
    port map (
            O => \N__47817\,
            I => \N__47682\
        );

    \I__11149\ : CascadeMux
    port map (
            O => \N__47816\,
            I => \N__47678\
        );

    \I__11148\ : CascadeMux
    port map (
            O => \N__47815\,
            I => \N__47674\
        );

    \I__11147\ : CascadeMux
    port map (
            O => \N__47814\,
            I => \N__47670\
        );

    \I__11146\ : CascadeMux
    port map (
            O => \N__47813\,
            I => \N__47666\
        );

    \I__11145\ : CascadeMux
    port map (
            O => \N__47812\,
            I => \N__47662\
        );

    \I__11144\ : CascadeMux
    port map (
            O => \N__47811\,
            I => \N__47658\
        );

    \I__11143\ : CascadeMux
    port map (
            O => \N__47810\,
            I => \N__47654\
        );

    \I__11142\ : CascadeMux
    port map (
            O => \N__47809\,
            I => \N__47650\
        );

    \I__11141\ : CascadeMux
    port map (
            O => \N__47808\,
            I => \N__47646\
        );

    \I__11140\ : CascadeMux
    port map (
            O => \N__47807\,
            I => \N__47642\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__47802\,
            I => \N__47638\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47801\,
            I => \N__47631\
        );

    \I__11137\ : InMux
    port map (
            O => \N__47800\,
            I => \N__47631\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47799\,
            I => \N__47631\
        );

    \I__11135\ : InMux
    port map (
            O => \N__47798\,
            I => \N__47624\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47797\,
            I => \N__47624\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47796\,
            I => \N__47624\
        );

    \I__11132\ : CascadeMux
    port map (
            O => \N__47795\,
            I => \N__47620\
        );

    \I__11131\ : LocalMux
    port map (
            O => \N__47792\,
            I => \N__47607\
        );

    \I__11130\ : InMux
    port map (
            O => \N__47791\,
            I => \N__47604\
        );

    \I__11129\ : InMux
    port map (
            O => \N__47788\,
            I => \N__47597\
        );

    \I__11128\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47597\
        );

    \I__11127\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47597\
        );

    \I__11126\ : LocalMux
    port map (
            O => \N__47769\,
            I => \N__47594\
        );

    \I__11125\ : InMux
    port map (
            O => \N__47768\,
            I => \N__47591\
        );

    \I__11124\ : LocalMux
    port map (
            O => \N__47763\,
            I => \N__47579\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__47758\,
            I => \N__47579\
        );

    \I__11122\ : InMux
    port map (
            O => \N__47757\,
            I => \N__47564\
        );

    \I__11121\ : InMux
    port map (
            O => \N__47756\,
            I => \N__47564\
        );

    \I__11120\ : InMux
    port map (
            O => \N__47755\,
            I => \N__47564\
        );

    \I__11119\ : InMux
    port map (
            O => \N__47754\,
            I => \N__47564\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47751\,
            I => \N__47564\
        );

    \I__11117\ : InMux
    port map (
            O => \N__47750\,
            I => \N__47564\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47747\,
            I => \N__47564\
        );

    \I__11115\ : InMux
    port map (
            O => \N__47746\,
            I => \N__47547\
        );

    \I__11114\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47547\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47744\,
            I => \N__47547\
        );

    \I__11112\ : InMux
    port map (
            O => \N__47743\,
            I => \N__47547\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47547\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47741\,
            I => \N__47547\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47740\,
            I => \N__47547\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47739\,
            I => \N__47547\
        );

    \I__11107\ : LocalMux
    port map (
            O => \N__47736\,
            I => \N__47542\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47733\,
            I => \N__47542\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47527\
        );

    \I__11104\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47527\
        );

    \I__11103\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47527\
        );

    \I__11102\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47527\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47722\,
            I => \N__47527\
        );

    \I__11100\ : InMux
    port map (
            O => \N__47721\,
            I => \N__47527\
        );

    \I__11099\ : InMux
    port map (
            O => \N__47718\,
            I => \N__47527\
        );

    \I__11098\ : LocalMux
    port map (
            O => \N__47701\,
            I => \N__47524\
        );

    \I__11097\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47507\
        );

    \I__11096\ : InMux
    port map (
            O => \N__47697\,
            I => \N__47507\
        );

    \I__11095\ : InMux
    port map (
            O => \N__47694\,
            I => \N__47507\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47693\,
            I => \N__47507\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47690\,
            I => \N__47507\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47689\,
            I => \N__47507\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47686\,
            I => \N__47507\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47685\,
            I => \N__47507\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47682\,
            I => \N__47490\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47681\,
            I => \N__47490\
        );

    \I__11087\ : InMux
    port map (
            O => \N__47678\,
            I => \N__47490\
        );

    \I__11086\ : InMux
    port map (
            O => \N__47677\,
            I => \N__47490\
        );

    \I__11085\ : InMux
    port map (
            O => \N__47674\,
            I => \N__47490\
        );

    \I__11084\ : InMux
    port map (
            O => \N__47673\,
            I => \N__47490\
        );

    \I__11083\ : InMux
    port map (
            O => \N__47670\,
            I => \N__47490\
        );

    \I__11082\ : InMux
    port map (
            O => \N__47669\,
            I => \N__47490\
        );

    \I__11081\ : InMux
    port map (
            O => \N__47666\,
            I => \N__47473\
        );

    \I__11080\ : InMux
    port map (
            O => \N__47665\,
            I => \N__47473\
        );

    \I__11079\ : InMux
    port map (
            O => \N__47662\,
            I => \N__47473\
        );

    \I__11078\ : InMux
    port map (
            O => \N__47661\,
            I => \N__47473\
        );

    \I__11077\ : InMux
    port map (
            O => \N__47658\,
            I => \N__47473\
        );

    \I__11076\ : InMux
    port map (
            O => \N__47657\,
            I => \N__47473\
        );

    \I__11075\ : InMux
    port map (
            O => \N__47654\,
            I => \N__47473\
        );

    \I__11074\ : InMux
    port map (
            O => \N__47653\,
            I => \N__47473\
        );

    \I__11073\ : InMux
    port map (
            O => \N__47650\,
            I => \N__47460\
        );

    \I__11072\ : InMux
    port map (
            O => \N__47649\,
            I => \N__47460\
        );

    \I__11071\ : InMux
    port map (
            O => \N__47646\,
            I => \N__47460\
        );

    \I__11070\ : InMux
    port map (
            O => \N__47645\,
            I => \N__47460\
        );

    \I__11069\ : InMux
    port map (
            O => \N__47642\,
            I => \N__47460\
        );

    \I__11068\ : InMux
    port map (
            O => \N__47641\,
            I => \N__47460\
        );

    \I__11067\ : Span12Mux_v
    port map (
            O => \N__47638\,
            I => \N__47455\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47631\,
            I => \N__47455\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__47624\,
            I => \N__47452\
        );

    \I__11064\ : InMux
    port map (
            O => \N__47623\,
            I => \N__47445\
        );

    \I__11063\ : InMux
    port map (
            O => \N__47620\,
            I => \N__47445\
        );

    \I__11062\ : InMux
    port map (
            O => \N__47619\,
            I => \N__47445\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47618\,
            I => \N__47430\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47617\,
            I => \N__47430\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47616\,
            I => \N__47430\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47615\,
            I => \N__47430\
        );

    \I__11057\ : InMux
    port map (
            O => \N__47614\,
            I => \N__47430\
        );

    \I__11056\ : InMux
    port map (
            O => \N__47613\,
            I => \N__47430\
        );

    \I__11055\ : InMux
    port map (
            O => \N__47612\,
            I => \N__47430\
        );

    \I__11054\ : CascadeMux
    port map (
            O => \N__47611\,
            I => \N__47423\
        );

    \I__11053\ : CascadeMux
    port map (
            O => \N__47610\,
            I => \N__47420\
        );

    \I__11052\ : Span4Mux_v
    port map (
            O => \N__47607\,
            I => \N__47407\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__47604\,
            I => \N__47407\
        );

    \I__11050\ : LocalMux
    port map (
            O => \N__47597\,
            I => \N__47407\
        );

    \I__11049\ : Span4Mux_h
    port map (
            O => \N__47594\,
            I => \N__47407\
        );

    \I__11048\ : LocalMux
    port map (
            O => \N__47591\,
            I => \N__47407\
        );

    \I__11047\ : CascadeMux
    port map (
            O => \N__47590\,
            I => \N__47404\
        );

    \I__11046\ : CascadeMux
    port map (
            O => \N__47589\,
            I => \N__47400\
        );

    \I__11045\ : CascadeMux
    port map (
            O => \N__47588\,
            I => \N__47396\
        );

    \I__11044\ : CascadeMux
    port map (
            O => \N__47587\,
            I => \N__47392\
        );

    \I__11043\ : CascadeMux
    port map (
            O => \N__47586\,
            I => \N__47388\
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__47585\,
            I => \N__47384\
        );

    \I__11041\ : CascadeMux
    port map (
            O => \N__47584\,
            I => \N__47380\
        );

    \I__11040\ : Span4Mux_h
    port map (
            O => \N__47579\,
            I => \N__47358\
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47564\,
            I => \N__47358\
        );

    \I__11038\ : LocalMux
    port map (
            O => \N__47547\,
            I => \N__47358\
        );

    \I__11037\ : Span4Mux_h
    port map (
            O => \N__47542\,
            I => \N__47358\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47527\,
            I => \N__47358\
        );

    \I__11035\ : Span4Mux_v
    port map (
            O => \N__47524\,
            I => \N__47358\
        );

    \I__11034\ : LocalMux
    port map (
            O => \N__47507\,
            I => \N__47358\
        );

    \I__11033\ : LocalMux
    port map (
            O => \N__47490\,
            I => \N__47358\
        );

    \I__11032\ : LocalMux
    port map (
            O => \N__47473\,
            I => \N__47358\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47460\,
            I => \N__47358\
        );

    \I__11030\ : Span12Mux_s11_h
    port map (
            O => \N__47455\,
            I => \N__47355\
        );

    \I__11029\ : Span4Mux_h
    port map (
            O => \N__47452\,
            I => \N__47348\
        );

    \I__11028\ : LocalMux
    port map (
            O => \N__47445\,
            I => \N__47348\
        );

    \I__11027\ : LocalMux
    port map (
            O => \N__47430\,
            I => \N__47348\
        );

    \I__11026\ : InMux
    port map (
            O => \N__47429\,
            I => \N__47335\
        );

    \I__11025\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47335\
        );

    \I__11024\ : InMux
    port map (
            O => \N__47427\,
            I => \N__47335\
        );

    \I__11023\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47335\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47423\,
            I => \N__47335\
        );

    \I__11021\ : InMux
    port map (
            O => \N__47420\,
            I => \N__47335\
        );

    \I__11020\ : InMux
    port map (
            O => \N__47419\,
            I => \N__47330\
        );

    \I__11019\ : InMux
    port map (
            O => \N__47418\,
            I => \N__47330\
        );

    \I__11018\ : Span4Mux_v
    port map (
            O => \N__47407\,
            I => \N__47327\
        );

    \I__11017\ : InMux
    port map (
            O => \N__47404\,
            I => \N__47310\
        );

    \I__11016\ : InMux
    port map (
            O => \N__47403\,
            I => \N__47310\
        );

    \I__11015\ : InMux
    port map (
            O => \N__47400\,
            I => \N__47310\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47399\,
            I => \N__47310\
        );

    \I__11013\ : InMux
    port map (
            O => \N__47396\,
            I => \N__47310\
        );

    \I__11012\ : InMux
    port map (
            O => \N__47395\,
            I => \N__47310\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47392\,
            I => \N__47310\
        );

    \I__11010\ : InMux
    port map (
            O => \N__47391\,
            I => \N__47310\
        );

    \I__11009\ : InMux
    port map (
            O => \N__47388\,
            I => \N__47297\
        );

    \I__11008\ : InMux
    port map (
            O => \N__47387\,
            I => \N__47297\
        );

    \I__11007\ : InMux
    port map (
            O => \N__47384\,
            I => \N__47297\
        );

    \I__11006\ : InMux
    port map (
            O => \N__47383\,
            I => \N__47297\
        );

    \I__11005\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47297\
        );

    \I__11004\ : InMux
    port map (
            O => \N__47379\,
            I => \N__47297\
        );

    \I__11003\ : Span4Mux_v
    port map (
            O => \N__47358\,
            I => \N__47294\
        );

    \I__11002\ : Odrv12
    port map (
            O => \N__47355\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11001\ : Odrv4
    port map (
            O => \N__47348\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__11000\ : LocalMux
    port map (
            O => \N__47335\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10999\ : LocalMux
    port map (
            O => \N__47330\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10998\ : Odrv4
    port map (
            O => \N__47327\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__47310\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10996\ : LocalMux
    port map (
            O => \N__47297\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10995\ : Odrv4
    port map (
            O => \N__47294\,
            I => \current_shift_inst.un38_control_input_5_2\
        );

    \I__10994\ : InMux
    port map (
            O => \N__47277\,
            I => \N__47274\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__47274\,
            I => \N__47269\
        );

    \I__10992\ : InMux
    port map (
            O => \N__47273\,
            I => \N__47266\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47272\,
            I => \N__47263\
        );

    \I__10990\ : Span4Mux_v
    port map (
            O => \N__47269\,
            I => \N__47260\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47266\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10988\ : LocalMux
    port map (
            O => \N__47263\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10987\ : Odrv4
    port map (
            O => \N__47260\,
            I => \current_shift_inst.un4_control_input1_14\
        );

    \I__10986\ : InMux
    port map (
            O => \N__47253\,
            I => \N__47250\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47250\,
            I => \N__47247\
        );

    \I__10984\ : Odrv12
    port map (
            O => \N__47247\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\
        );

    \I__10983\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47240\
        );

    \I__10982\ : CascadeMux
    port map (
            O => \N__47243\,
            I => \N__47237\
        );

    \I__10981\ : LocalMux
    port map (
            O => \N__47240\,
            I => \N__47234\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47237\,
            I => \N__47229\
        );

    \I__10979\ : Span4Mux_h
    port map (
            O => \N__47234\,
            I => \N__47226\
        );

    \I__10978\ : InMux
    port map (
            O => \N__47233\,
            I => \N__47221\
        );

    \I__10977\ : InMux
    port map (
            O => \N__47232\,
            I => \N__47221\
        );

    \I__10976\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47218\
        );

    \I__10975\ : Odrv4
    port map (
            O => \N__47226\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__47221\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10973\ : Odrv4
    port map (
            O => \N__47218\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\
        );

    \I__10972\ : InMux
    port map (
            O => \N__47211\,
            I => \N__47208\
        );

    \I__10971\ : LocalMux
    port map (
            O => \N__47208\,
            I => \N__47205\
        );

    \I__10970\ : Span4Mux_h
    port map (
            O => \N__47205\,
            I => \N__47202\
        );

    \I__10969\ : Span4Mux_h
    port map (
            O => \N__47202\,
            I => \N__47198\
        );

    \I__10968\ : InMux
    port map (
            O => \N__47201\,
            I => \N__47195\
        );

    \I__10967\ : Odrv4
    port map (
            O => \N__47198\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__47195\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18\
        );

    \I__10965\ : InMux
    port map (
            O => \N__47190\,
            I => \N__47184\
        );

    \I__10964\ : InMux
    port map (
            O => \N__47189\,
            I => \N__47184\
        );

    \I__10963\ : LocalMux
    port map (
            O => \N__47184\,
            I => \N__47181\
        );

    \I__10962\ : Odrv12
    port map (
            O => \N__47181\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\
        );

    \I__10961\ : CascadeMux
    port map (
            O => \N__47178\,
            I => \N__47175\
        );

    \I__10960\ : InMux
    port map (
            O => \N__47175\,
            I => \N__47169\
        );

    \I__10959\ : InMux
    port map (
            O => \N__47174\,
            I => \N__47169\
        );

    \I__10958\ : LocalMux
    port map (
            O => \N__47169\,
            I => \N__47166\
        );

    \I__10957\ : Odrv12
    port map (
            O => \N__47166\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\
        );

    \I__10956\ : CEMux
    port map (
            O => \N__47163\,
            I => \N__47127\
        );

    \I__10955\ : CEMux
    port map (
            O => \N__47162\,
            I => \N__47127\
        );

    \I__10954\ : CEMux
    port map (
            O => \N__47161\,
            I => \N__47127\
        );

    \I__10953\ : CEMux
    port map (
            O => \N__47160\,
            I => \N__47127\
        );

    \I__10952\ : CEMux
    port map (
            O => \N__47159\,
            I => \N__47127\
        );

    \I__10951\ : CEMux
    port map (
            O => \N__47158\,
            I => \N__47127\
        );

    \I__10950\ : CEMux
    port map (
            O => \N__47157\,
            I => \N__47127\
        );

    \I__10949\ : CEMux
    port map (
            O => \N__47156\,
            I => \N__47127\
        );

    \I__10948\ : CEMux
    port map (
            O => \N__47155\,
            I => \N__47127\
        );

    \I__10947\ : CEMux
    port map (
            O => \N__47154\,
            I => \N__47127\
        );

    \I__10946\ : CEMux
    port map (
            O => \N__47153\,
            I => \N__47127\
        );

    \I__10945\ : CEMux
    port map (
            O => \N__47152\,
            I => \N__47127\
        );

    \I__10944\ : GlobalMux
    port map (
            O => \N__47127\,
            I => \N__47124\
        );

    \I__10943\ : gio2CtrlBuf
    port map (
            O => \N__47124\,
            I => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \I__10942\ : InMux
    port map (
            O => \N__47121\,
            I => \N__47117\
        );

    \I__10941\ : InMux
    port map (
            O => \N__47120\,
            I => \N__47114\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__47117\,
            I => \N__47109\
        );

    \I__10939\ : LocalMux
    port map (
            O => \N__47114\,
            I => \N__47106\
        );

    \I__10938\ : InMux
    port map (
            O => \N__47113\,
            I => \N__47103\
        );

    \I__10937\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47100\
        );

    \I__10936\ : Span4Mux_v
    port map (
            O => \N__47109\,
            I => \N__47097\
        );

    \I__10935\ : Span4Mux_v
    port map (
            O => \N__47106\,
            I => \N__47092\
        );

    \I__10934\ : LocalMux
    port map (
            O => \N__47103\,
            I => \N__47092\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__47100\,
            I => \N__47089\
        );

    \I__10932\ : Span4Mux_h
    port map (
            O => \N__47097\,
            I => \N__47084\
        );

    \I__10931\ : Span4Mux_h
    port map (
            O => \N__47092\,
            I => \N__47084\
        );

    \I__10930\ : Span4Mux_v
    port map (
            O => \N__47089\,
            I => \N__47081\
        );

    \I__10929\ : Odrv4
    port map (
            O => \N__47084\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__10928\ : Odrv4
    port map (
            O => \N__47081\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\
        );

    \I__10927\ : InMux
    port map (
            O => \N__47076\,
            I => \N__47071\
        );

    \I__10926\ : InMux
    port map (
            O => \N__47075\,
            I => \N__47064\
        );

    \I__10925\ : InMux
    port map (
            O => \N__47074\,
            I => \N__47064\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__47071\,
            I => \N__47061\
        );

    \I__10923\ : InMux
    port map (
            O => \N__47070\,
            I => \N__47052\
        );

    \I__10922\ : InMux
    port map (
            O => \N__47069\,
            I => \N__47049\
        );

    \I__10921\ : LocalMux
    port map (
            O => \N__47064\,
            I => \N__47017\
        );

    \I__10920\ : Span4Mux_h
    port map (
            O => \N__47061\,
            I => \N__47014\
        );

    \I__10919\ : InMux
    port map (
            O => \N__47060\,
            I => \N__47007\
        );

    \I__10918\ : InMux
    port map (
            O => \N__47059\,
            I => \N__47007\
        );

    \I__10917\ : InMux
    port map (
            O => \N__47058\,
            I => \N__47007\
        );

    \I__10916\ : InMux
    port map (
            O => \N__47057\,
            I => \N__47000\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47056\,
            I => \N__47000\
        );

    \I__10914\ : InMux
    port map (
            O => \N__47055\,
            I => \N__47000\
        );

    \I__10913\ : LocalMux
    port map (
            O => \N__47052\,
            I => \N__46995\
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__47049\,
            I => \N__46995\
        );

    \I__10911\ : InMux
    port map (
            O => \N__47048\,
            I => \N__46992\
        );

    \I__10910\ : InMux
    port map (
            O => \N__47047\,
            I => \N__46988\
        );

    \I__10909\ : InMux
    port map (
            O => \N__47046\,
            I => \N__46979\
        );

    \I__10908\ : InMux
    port map (
            O => \N__47045\,
            I => \N__46979\
        );

    \I__10907\ : InMux
    port map (
            O => \N__47044\,
            I => \N__46979\
        );

    \I__10906\ : InMux
    port map (
            O => \N__47043\,
            I => \N__46979\
        );

    \I__10905\ : InMux
    port map (
            O => \N__47042\,
            I => \N__46972\
        );

    \I__10904\ : InMux
    port map (
            O => \N__47041\,
            I => \N__46972\
        );

    \I__10903\ : InMux
    port map (
            O => \N__47040\,
            I => \N__46972\
        );

    \I__10902\ : CascadeMux
    port map (
            O => \N__47039\,
            I => \N__46966\
        );

    \I__10901\ : InMux
    port map (
            O => \N__47038\,
            I => \N__46961\
        );

    \I__10900\ : InMux
    port map (
            O => \N__47037\,
            I => \N__46944\
        );

    \I__10899\ : InMux
    port map (
            O => \N__47036\,
            I => \N__46944\
        );

    \I__10898\ : InMux
    port map (
            O => \N__47035\,
            I => \N__46944\
        );

    \I__10897\ : InMux
    port map (
            O => \N__47034\,
            I => \N__46944\
        );

    \I__10896\ : InMux
    port map (
            O => \N__47033\,
            I => \N__46944\
        );

    \I__10895\ : InMux
    port map (
            O => \N__47032\,
            I => \N__46937\
        );

    \I__10894\ : InMux
    port map (
            O => \N__47031\,
            I => \N__46922\
        );

    \I__10893\ : InMux
    port map (
            O => \N__47030\,
            I => \N__46922\
        );

    \I__10892\ : InMux
    port map (
            O => \N__47029\,
            I => \N__46922\
        );

    \I__10891\ : InMux
    port map (
            O => \N__47028\,
            I => \N__46922\
        );

    \I__10890\ : InMux
    port map (
            O => \N__47027\,
            I => \N__46922\
        );

    \I__10889\ : InMux
    port map (
            O => \N__47026\,
            I => \N__46903\
        );

    \I__10888\ : InMux
    port map (
            O => \N__47025\,
            I => \N__46903\
        );

    \I__10887\ : InMux
    port map (
            O => \N__47024\,
            I => \N__46903\
        );

    \I__10886\ : InMux
    port map (
            O => \N__47023\,
            I => \N__46903\
        );

    \I__10885\ : InMux
    port map (
            O => \N__47022\,
            I => \N__46896\
        );

    \I__10884\ : InMux
    port map (
            O => \N__47021\,
            I => \N__46896\
        );

    \I__10883\ : InMux
    port map (
            O => \N__47020\,
            I => \N__46896\
        );

    \I__10882\ : Span4Mux_h
    port map (
            O => \N__47017\,
            I => \N__46889\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__47014\,
            I => \N__46889\
        );

    \I__10880\ : LocalMux
    port map (
            O => \N__47007\,
            I => \N__46889\
        );

    \I__10879\ : LocalMux
    port map (
            O => \N__47000\,
            I => \N__46882\
        );

    \I__10878\ : Span4Mux_v
    port map (
            O => \N__46995\,
            I => \N__46882\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__46992\,
            I => \N__46882\
        );

    \I__10876\ : CascadeMux
    port map (
            O => \N__46991\,
            I => \N__46876\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__46988\,
            I => \N__46867\
        );

    \I__10874\ : LocalMux
    port map (
            O => \N__46979\,
            I => \N__46867\
        );

    \I__10873\ : LocalMux
    port map (
            O => \N__46972\,
            I => \N__46867\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46971\,
            I => \N__46854\
        );

    \I__10871\ : InMux
    port map (
            O => \N__46970\,
            I => \N__46854\
        );

    \I__10870\ : InMux
    port map (
            O => \N__46969\,
            I => \N__46854\
        );

    \I__10869\ : InMux
    port map (
            O => \N__46966\,
            I => \N__46854\
        );

    \I__10868\ : InMux
    port map (
            O => \N__46965\,
            I => \N__46854\
        );

    \I__10867\ : InMux
    port map (
            O => \N__46964\,
            I => \N__46854\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__46961\,
            I => \N__46846\
        );

    \I__10865\ : InMux
    port map (
            O => \N__46960\,
            I => \N__46835\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46959\,
            I => \N__46835\
        );

    \I__10863\ : InMux
    port map (
            O => \N__46958\,
            I => \N__46835\
        );

    \I__10862\ : InMux
    port map (
            O => \N__46957\,
            I => \N__46835\
        );

    \I__10861\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46835\
        );

    \I__10860\ : InMux
    port map (
            O => \N__46955\,
            I => \N__46832\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__46944\,
            I => \N__46827\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46943\,
            I => \N__46818\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46818\
        );

    \I__10856\ : InMux
    port map (
            O => \N__46941\,
            I => \N__46818\
        );

    \I__10855\ : InMux
    port map (
            O => \N__46940\,
            I => \N__46818\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46937\,
            I => \N__46808\
        );

    \I__10853\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46805\
        );

    \I__10852\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46798\
        );

    \I__10851\ : InMux
    port map (
            O => \N__46934\,
            I => \N__46798\
        );

    \I__10850\ : InMux
    port map (
            O => \N__46933\,
            I => \N__46798\
        );

    \I__10849\ : LocalMux
    port map (
            O => \N__46922\,
            I => \N__46795\
        );

    \I__10848\ : InMux
    port map (
            O => \N__46921\,
            I => \N__46782\
        );

    \I__10847\ : InMux
    port map (
            O => \N__46920\,
            I => \N__46782\
        );

    \I__10846\ : InMux
    port map (
            O => \N__46919\,
            I => \N__46782\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46918\,
            I => \N__46782\
        );

    \I__10844\ : InMux
    port map (
            O => \N__46917\,
            I => \N__46782\
        );

    \I__10843\ : InMux
    port map (
            O => \N__46916\,
            I => \N__46782\
        );

    \I__10842\ : InMux
    port map (
            O => \N__46915\,
            I => \N__46775\
        );

    \I__10841\ : InMux
    port map (
            O => \N__46914\,
            I => \N__46775\
        );

    \I__10840\ : InMux
    port map (
            O => \N__46913\,
            I => \N__46775\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46912\,
            I => \N__46772\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46903\,
            I => \N__46763\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__46896\,
            I => \N__46763\
        );

    \I__10836\ : Span4Mux_h
    port map (
            O => \N__46889\,
            I => \N__46763\
        );

    \I__10835\ : Span4Mux_h
    port map (
            O => \N__46882\,
            I => \N__46763\
        );

    \I__10834\ : InMux
    port map (
            O => \N__46881\,
            I => \N__46760\
        );

    \I__10833\ : InMux
    port map (
            O => \N__46880\,
            I => \N__46749\
        );

    \I__10832\ : InMux
    port map (
            O => \N__46879\,
            I => \N__46749\
        );

    \I__10831\ : InMux
    port map (
            O => \N__46876\,
            I => \N__46749\
        );

    \I__10830\ : InMux
    port map (
            O => \N__46875\,
            I => \N__46749\
        );

    \I__10829\ : InMux
    port map (
            O => \N__46874\,
            I => \N__46749\
        );

    \I__10828\ : Span4Mux_v
    port map (
            O => \N__46867\,
            I => \N__46744\
        );

    \I__10827\ : LocalMux
    port map (
            O => \N__46854\,
            I => \N__46744\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46853\,
            I => \N__46733\
        );

    \I__10825\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46733\
        );

    \I__10824\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46733\
        );

    \I__10823\ : InMux
    port map (
            O => \N__46850\,
            I => \N__46733\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46849\,
            I => \N__46733\
        );

    \I__10821\ : Span4Mux_h
    port map (
            O => \N__46846\,
            I => \N__46728\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46835\,
            I => \N__46728\
        );

    \I__10819\ : LocalMux
    port map (
            O => \N__46832\,
            I => \N__46725\
        );

    \I__10818\ : InMux
    port map (
            O => \N__46831\,
            I => \N__46717\
        );

    \I__10817\ : InMux
    port map (
            O => \N__46830\,
            I => \N__46717\
        );

    \I__10816\ : Span4Mux_v
    port map (
            O => \N__46827\,
            I => \N__46712\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46818\,
            I => \N__46712\
        );

    \I__10814\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46703\
        );

    \I__10813\ : InMux
    port map (
            O => \N__46816\,
            I => \N__46703\
        );

    \I__10812\ : InMux
    port map (
            O => \N__46815\,
            I => \N__46703\
        );

    \I__10811\ : InMux
    port map (
            O => \N__46814\,
            I => \N__46703\
        );

    \I__10810\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46696\
        );

    \I__10809\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46696\
        );

    \I__10808\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46696\
        );

    \I__10807\ : Span4Mux_v
    port map (
            O => \N__46808\,
            I => \N__46689\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46805\,
            I => \N__46689\
        );

    \I__10805\ : LocalMux
    port map (
            O => \N__46798\,
            I => \N__46689\
        );

    \I__10804\ : Span4Mux_h
    port map (
            O => \N__46795\,
            I => \N__46686\
        );

    \I__10803\ : LocalMux
    port map (
            O => \N__46782\,
            I => \N__46681\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__46775\,
            I => \N__46681\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46772\,
            I => \N__46676\
        );

    \I__10800\ : Span4Mux_v
    port map (
            O => \N__46763\,
            I => \N__46676\
        );

    \I__10799\ : LocalMux
    port map (
            O => \N__46760\,
            I => \N__46671\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46749\,
            I => \N__46671\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__46744\,
            I => \N__46664\
        );

    \I__10796\ : LocalMux
    port map (
            O => \N__46733\,
            I => \N__46664\
        );

    \I__10795\ : Span4Mux_v
    port map (
            O => \N__46728\,
            I => \N__46664\
        );

    \I__10794\ : Span4Mux_h
    port map (
            O => \N__46725\,
            I => \N__46661\
        );

    \I__10793\ : InMux
    port map (
            O => \N__46724\,
            I => \N__46658\
        );

    \I__10792\ : InMux
    port map (
            O => \N__46723\,
            I => \N__46653\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46722\,
            I => \N__46653\
        );

    \I__10790\ : LocalMux
    port map (
            O => \N__46717\,
            I => \N__46648\
        );

    \I__10789\ : Span4Mux_v
    port map (
            O => \N__46712\,
            I => \N__46648\
        );

    \I__10788\ : LocalMux
    port map (
            O => \N__46703\,
            I => \N__46639\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46696\,
            I => \N__46639\
        );

    \I__10786\ : Span4Mux_h
    port map (
            O => \N__46689\,
            I => \N__46639\
        );

    \I__10785\ : Span4Mux_v
    port map (
            O => \N__46686\,
            I => \N__46639\
        );

    \I__10784\ : Span4Mux_v
    port map (
            O => \N__46681\,
            I => \N__46634\
        );

    \I__10783\ : Span4Mux_h
    port map (
            O => \N__46676\,
            I => \N__46634\
        );

    \I__10782\ : Span4Mux_h
    port map (
            O => \N__46671\,
            I => \N__46629\
        );

    \I__10781\ : Span4Mux_v
    port map (
            O => \N__46664\,
            I => \N__46629\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__46661\,
            I => \N__46626\
        );

    \I__10779\ : LocalMux
    port map (
            O => \N__46658\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__46653\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10777\ : Odrv4
    port map (
            O => \N__46648\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10776\ : Odrv4
    port map (
            O => \N__46639\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10775\ : Odrv4
    port map (
            O => \N__46634\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10774\ : Odrv4
    port map (
            O => \N__46629\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10773\ : Odrv4
    port map (
            O => \N__46626\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46611\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_28\
        );

    \I__10771\ : InMux
    port map (
            O => \N__46608\,
            I => \N__46605\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46605\,
            I => \N__46601\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46604\,
            I => \N__46598\
        );

    \I__10768\ : Span4Mux_h
    port map (
            O => \N__46601\,
            I => \N__46595\
        );

    \I__10767\ : LocalMux
    port map (
            O => \N__46598\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10766\ : Odrv4
    port map (
            O => \N__46595\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\
        );

    \I__10765\ : InMux
    port map (
            O => \N__46590\,
            I => \N__46587\
        );

    \I__10764\ : LocalMux
    port map (
            O => \N__46587\,
            I => \N__46584\
        );

    \I__10763\ : Span4Mux_h
    port map (
            O => \N__46584\,
            I => \N__46581\
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__46581\,
            I => \current_shift_inst.un38_control_input_axb_31_s0\
        );

    \I__10761\ : CascadeMux
    port map (
            O => \N__46578\,
            I => \N__46573\
        );

    \I__10760\ : InMux
    port map (
            O => \N__46577\,
            I => \N__46570\
        );

    \I__10759\ : InMux
    port map (
            O => \N__46576\,
            I => \N__46567\
        );

    \I__10758\ : InMux
    port map (
            O => \N__46573\,
            I => \N__46564\
        );

    \I__10757\ : LocalMux
    port map (
            O => \N__46570\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10756\ : LocalMux
    port map (
            O => \N__46567\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10755\ : LocalMux
    port map (
            O => \N__46564\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1\
        );

    \I__10754\ : CascadeMux
    port map (
            O => \N__46557\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__46554\,
            I => \N__46550\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46553\,
            I => \N__46547\
        );

    \I__10751\ : InMux
    port map (
            O => \N__46550\,
            I => \N__46544\
        );

    \I__10750\ : LocalMux
    port map (
            O => \N__46547\,
            I => \N__46539\
        );

    \I__10749\ : LocalMux
    port map (
            O => \N__46544\,
            I => \N__46539\
        );

    \I__10748\ : Span4Mux_h
    port map (
            O => \N__46539\,
            I => \N__46536\
        );

    \I__10747\ : Span4Mux_v
    port map (
            O => \N__46536\,
            I => \N__46533\
        );

    \I__10746\ : Odrv4
    port map (
            O => \N__46533\,
            I => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\
        );

    \I__10745\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46526\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46529\,
            I => \N__46522\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46526\,
            I => \N__46519\
        );

    \I__10742\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46516\
        );

    \I__10741\ : LocalMux
    port map (
            O => \N__46522\,
            I => \N__46513\
        );

    \I__10740\ : Span4Mux_v
    port map (
            O => \N__46519\,
            I => \N__46510\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46516\,
            I => \N__46507\
        );

    \I__10738\ : Span12Mux_v
    port map (
            O => \N__46513\,
            I => \N__46504\
        );

    \I__10737\ : Span4Mux_v
    port map (
            O => \N__46510\,
            I => \N__46499\
        );

    \I__10736\ : Span4Mux_v
    port map (
            O => \N__46507\,
            I => \N__46499\
        );

    \I__10735\ : Odrv12
    port map (
            O => \N__46504\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10734\ : Odrv4
    port map (
            O => \N__46499\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\
        );

    \I__10733\ : InMux
    port map (
            O => \N__46494\,
            I => \N__46491\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__46491\,
            I => \N__46487\
        );

    \I__10731\ : InMux
    port map (
            O => \N__46490\,
            I => \N__46484\
        );

    \I__10730\ : Span4Mux_h
    port map (
            O => \N__46487\,
            I => \N__46480\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__46484\,
            I => \N__46477\
        );

    \I__10728\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46474\
        );

    \I__10727\ : Span4Mux_v
    port map (
            O => \N__46480\,
            I => \N__46469\
        );

    \I__10726\ : Span4Mux_h
    port map (
            O => \N__46477\,
            I => \N__46469\
        );

    \I__10725\ : LocalMux
    port map (
            O => \N__46474\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10724\ : Odrv4
    port map (
            O => \N__46469\,
            I => \current_shift_inst.timer_s1.counterZ0Z_0\
        );

    \I__10723\ : InMux
    port map (
            O => \N__46464\,
            I => \N__46461\
        );

    \I__10722\ : LocalMux
    port map (
            O => \N__46461\,
            I => \N__46455\
        );

    \I__10721\ : InMux
    port map (
            O => \N__46460\,
            I => \N__46452\
        );

    \I__10720\ : InMux
    port map (
            O => \N__46459\,
            I => \N__46447\
        );

    \I__10719\ : InMux
    port map (
            O => \N__46458\,
            I => \N__46447\
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__46455\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10717\ : LocalMux
    port map (
            O => \N__46452\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46447\,
            I => \current_shift_inst.elapsed_time_ns_s1_1\
        );

    \I__10715\ : InMux
    port map (
            O => \N__46440\,
            I => \N__46436\
        );

    \I__10714\ : InMux
    port map (
            O => \N__46439\,
            I => \N__46433\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__46436\,
            I => \N__46429\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__46433\,
            I => \N__46426\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46432\,
            I => \N__46423\
        );

    \I__10710\ : Span4Mux_v
    port map (
            O => \N__46429\,
            I => \N__46418\
        );

    \I__10709\ : Span4Mux_h
    port map (
            O => \N__46426\,
            I => \N__46418\
        );

    \I__10708\ : LocalMux
    port map (
            O => \N__46423\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10707\ : Odrv4
    port map (
            O => \N__46418\,
            I => \current_shift_inst.timer_s1.counterZ0Z_1\
        );

    \I__10706\ : CEMux
    port map (
            O => \N__46413\,
            I => \N__46389\
        );

    \I__10705\ : CEMux
    port map (
            O => \N__46412\,
            I => \N__46389\
        );

    \I__10704\ : CEMux
    port map (
            O => \N__46411\,
            I => \N__46389\
        );

    \I__10703\ : CEMux
    port map (
            O => \N__46410\,
            I => \N__46389\
        );

    \I__10702\ : CEMux
    port map (
            O => \N__46409\,
            I => \N__46389\
        );

    \I__10701\ : CEMux
    port map (
            O => \N__46408\,
            I => \N__46389\
        );

    \I__10700\ : CEMux
    port map (
            O => \N__46407\,
            I => \N__46389\
        );

    \I__10699\ : CEMux
    port map (
            O => \N__46406\,
            I => \N__46389\
        );

    \I__10698\ : GlobalMux
    port map (
            O => \N__46389\,
            I => \N__46386\
        );

    \I__10697\ : gio2CtrlBuf
    port map (
            O => \N__46386\,
            I => \current_shift_inst.timer_s1.N_161_i_g\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46383\,
            I => \N__46380\
        );

    \I__10695\ : LocalMux
    port map (
            O => \N__46380\,
            I => \current_shift_inst.un4_control_input_1_axb_1\
        );

    \I__10694\ : CascadeMux
    port map (
            O => \N__46377\,
            I => \N__46373\
        );

    \I__10693\ : CascadeMux
    port map (
            O => \N__46376\,
            I => \N__46370\
        );

    \I__10692\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46366\
        );

    \I__10691\ : InMux
    port map (
            O => \N__46370\,
            I => \N__46363\
        );

    \I__10690\ : InMux
    port map (
            O => \N__46369\,
            I => \N__46360\
        );

    \I__10689\ : LocalMux
    port map (
            O => \N__46366\,
            I => \N__46354\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__46363\,
            I => \N__46354\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__46360\,
            I => \N__46351\
        );

    \I__10686\ : InMux
    port map (
            O => \N__46359\,
            I => \N__46348\
        );

    \I__10685\ : Span4Mux_v
    port map (
            O => \N__46354\,
            I => \N__46343\
        );

    \I__10684\ : Span4Mux_v
    port map (
            O => \N__46351\,
            I => \N__46343\
        );

    \I__10683\ : LocalMux
    port map (
            O => \N__46348\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10682\ : Odrv4
    port map (
            O => \N__46343\,
            I => \current_shift_inst.un38_control_input_5_1\
        );

    \I__10681\ : CascadeMux
    port map (
            O => \N__46338\,
            I => \N__46335\
        );

    \I__10680\ : InMux
    port map (
            O => \N__46335\,
            I => \N__46332\
        );

    \I__10679\ : LocalMux
    port map (
            O => \N__46332\,
            I => \N__46329\
        );

    \I__10678\ : Odrv12
    port map (
            O => \N__46329\,
            I => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\
        );

    \I__10677\ : CascadeMux
    port map (
            O => \N__46326\,
            I => \N__46323\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46323\,
            I => \N__46319\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46322\,
            I => \N__46316\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__46319\,
            I => \N__46310\
        );

    \I__10673\ : LocalMux
    port map (
            O => \N__46316\,
            I => \N__46310\
        );

    \I__10672\ : InMux
    port map (
            O => \N__46315\,
            I => \N__46307\
        );

    \I__10671\ : Span4Mux_h
    port map (
            O => \N__46310\,
            I => \N__46304\
        );

    \I__10670\ : LocalMux
    port map (
            O => \N__46307\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10669\ : Odrv4
    port map (
            O => \N__46304\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\
        );

    \I__10668\ : InMux
    port map (
            O => \N__46299\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_20\
        );

    \I__10667\ : CascadeMux
    port map (
            O => \N__46296\,
            I => \N__46293\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46289\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46292\,
            I => \N__46286\
        );

    \I__10664\ : LocalMux
    port map (
            O => \N__46289\,
            I => \N__46280\
        );

    \I__10663\ : LocalMux
    port map (
            O => \N__46286\,
            I => \N__46280\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46285\,
            I => \N__46277\
        );

    \I__10661\ : Span4Mux_v
    port map (
            O => \N__46280\,
            I => \N__46274\
        );

    \I__10660\ : LocalMux
    port map (
            O => \N__46277\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__46274\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\
        );

    \I__10658\ : InMux
    port map (
            O => \N__46269\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_21\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46266\,
            I => \N__46260\
        );

    \I__10656\ : InMux
    port map (
            O => \N__46265\,
            I => \N__46260\
        );

    \I__10655\ : LocalMux
    port map (
            O => \N__46260\,
            I => \N__46256\
        );

    \I__10654\ : InMux
    port map (
            O => \N__46259\,
            I => \N__46253\
        );

    \I__10653\ : Span4Mux_h
    port map (
            O => \N__46256\,
            I => \N__46250\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__46253\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__46250\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\
        );

    \I__10650\ : InMux
    port map (
            O => \N__46245\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_22\
        );

    \I__10649\ : CascadeMux
    port map (
            O => \N__46242\,
            I => \N__46239\
        );

    \I__10648\ : InMux
    port map (
            O => \N__46239\,
            I => \N__46234\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46238\,
            I => \N__46231\
        );

    \I__10646\ : InMux
    port map (
            O => \N__46237\,
            I => \N__46228\
        );

    \I__10645\ : LocalMux
    port map (
            O => \N__46234\,
            I => \N__46225\
        );

    \I__10644\ : LocalMux
    port map (
            O => \N__46231\,
            I => \N__46222\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46228\,
            I => \N__46217\
        );

    \I__10642\ : Span4Mux_v
    port map (
            O => \N__46225\,
            I => \N__46217\
        );

    \I__10641\ : Span4Mux_h
    port map (
            O => \N__46222\,
            I => \N__46214\
        );

    \I__10640\ : Odrv4
    port map (
            O => \N__46217\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10639\ : Odrv4
    port map (
            O => \N__46214\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\
        );

    \I__10638\ : InMux
    port map (
            O => \N__46209\,
            I => \bfn_18_14_0_\
        );

    \I__10637\ : CascadeMux
    port map (
            O => \N__46206\,
            I => \N__46202\
        );

    \I__10636\ : CascadeMux
    port map (
            O => \N__46205\,
            I => \N__46199\
        );

    \I__10635\ : InMux
    port map (
            O => \N__46202\,
            I => \N__46196\
        );

    \I__10634\ : InMux
    port map (
            O => \N__46199\,
            I => \N__46193\
        );

    \I__10633\ : LocalMux
    port map (
            O => \N__46196\,
            I => \N__46189\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46193\,
            I => \N__46186\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46192\,
            I => \N__46183\
        );

    \I__10630\ : Span4Mux_v
    port map (
            O => \N__46189\,
            I => \N__46180\
        );

    \I__10629\ : Span4Mux_h
    port map (
            O => \N__46186\,
            I => \N__46177\
        );

    \I__10628\ : LocalMux
    port map (
            O => \N__46183\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10627\ : Odrv4
    port map (
            O => \N__46180\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10626\ : Odrv4
    port map (
            O => \N__46177\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\
        );

    \I__10625\ : InMux
    port map (
            O => \N__46170\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_24\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46167\,
            I => \N__46161\
        );

    \I__10623\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46161\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__46161\,
            I => \N__46157\
        );

    \I__10621\ : InMux
    port map (
            O => \N__46160\,
            I => \N__46154\
        );

    \I__10620\ : Span4Mux_h
    port map (
            O => \N__46157\,
            I => \N__46151\
        );

    \I__10619\ : LocalMux
    port map (
            O => \N__46154\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10618\ : Odrv4
    port map (
            O => \N__46151\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\
        );

    \I__10617\ : InMux
    port map (
            O => \N__46146\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_25\
        );

    \I__10616\ : CascadeMux
    port map (
            O => \N__46143\,
            I => \N__46140\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46140\,
            I => \N__46136\
        );

    \I__10614\ : InMux
    port map (
            O => \N__46139\,
            I => \N__46133\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__46136\,
            I => \N__46127\
        );

    \I__10612\ : LocalMux
    port map (
            O => \N__46133\,
            I => \N__46127\
        );

    \I__10611\ : InMux
    port map (
            O => \N__46132\,
            I => \N__46124\
        );

    \I__10610\ : Span4Mux_h
    port map (
            O => \N__46127\,
            I => \N__46121\
        );

    \I__10609\ : LocalMux
    port map (
            O => \N__46124\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10608\ : Odrv4
    port map (
            O => \N__46121\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46116\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_26\
        );

    \I__10606\ : CascadeMux
    port map (
            O => \N__46113\,
            I => \N__46110\
        );

    \I__10605\ : InMux
    port map (
            O => \N__46110\,
            I => \N__46107\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__46107\,
            I => \N__46103\
        );

    \I__10603\ : InMux
    port map (
            O => \N__46106\,
            I => \N__46100\
        );

    \I__10602\ : Span4Mux_h
    port map (
            O => \N__46103\,
            I => \N__46097\
        );

    \I__10601\ : LocalMux
    port map (
            O => \N__46100\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10600\ : Odrv4
    port map (
            O => \N__46097\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\
        );

    \I__10599\ : InMux
    port map (
            O => \N__46092\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_27\
        );

    \I__10598\ : CascadeMux
    port map (
            O => \N__46089\,
            I => \N__46086\
        );

    \I__10597\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46082\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46085\,
            I => \N__46079\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__46082\,
            I => \N__46073\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__46079\,
            I => \N__46073\
        );

    \I__10593\ : InMux
    port map (
            O => \N__46078\,
            I => \N__46070\
        );

    \I__10592\ : Span4Mux_h
    port map (
            O => \N__46073\,
            I => \N__46067\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__46070\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10590\ : Odrv4
    port map (
            O => \N__46067\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\
        );

    \I__10589\ : InMux
    port map (
            O => \N__46062\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_11\
        );

    \I__10588\ : CascadeMux
    port map (
            O => \N__46059\,
            I => \N__46055\
        );

    \I__10587\ : CascadeMux
    port map (
            O => \N__46058\,
            I => \N__46052\
        );

    \I__10586\ : InMux
    port map (
            O => \N__46055\,
            I => \N__46047\
        );

    \I__10585\ : InMux
    port map (
            O => \N__46052\,
            I => \N__46047\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__46047\,
            I => \N__46043\
        );

    \I__10583\ : InMux
    port map (
            O => \N__46046\,
            I => \N__46040\
        );

    \I__10582\ : Span4Mux_h
    port map (
            O => \N__46043\,
            I => \N__46037\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__46040\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10580\ : Odrv4
    port map (
            O => \N__46037\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\
        );

    \I__10579\ : InMux
    port map (
            O => \N__46032\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_12\
        );

    \I__10578\ : CascadeMux
    port map (
            O => \N__46029\,
            I => \N__46026\
        );

    \I__10577\ : InMux
    port map (
            O => \N__46026\,
            I => \N__46022\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46025\,
            I => \N__46019\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__46022\,
            I => \N__46013\
        );

    \I__10574\ : LocalMux
    port map (
            O => \N__46019\,
            I => \N__46013\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46018\,
            I => \N__46010\
        );

    \I__10572\ : Span4Mux_h
    port map (
            O => \N__46013\,
            I => \N__46007\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46010\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10570\ : Odrv4
    port map (
            O => \N__46007\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\
        );

    \I__10569\ : InMux
    port map (
            O => \N__46002\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_13\
        );

    \I__10568\ : InMux
    port map (
            O => \N__45999\,
            I => \N__45992\
        );

    \I__10567\ : InMux
    port map (
            O => \N__45998\,
            I => \N__45992\
        );

    \I__10566\ : InMux
    port map (
            O => \N__45997\,
            I => \N__45989\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__45992\,
            I => \N__45986\
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__45989\,
            I => \N__45981\
        );

    \I__10563\ : Span4Mux_v
    port map (
            O => \N__45986\,
            I => \N__45981\
        );

    \I__10562\ : Odrv4
    port map (
            O => \N__45981\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\
        );

    \I__10561\ : InMux
    port map (
            O => \N__45978\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_14\
        );

    \I__10560\ : CascadeMux
    port map (
            O => \N__45975\,
            I => \N__45972\
        );

    \I__10559\ : InMux
    port map (
            O => \N__45972\,
            I => \N__45968\
        );

    \I__10558\ : InMux
    port map (
            O => \N__45971\,
            I => \N__45965\
        );

    \I__10557\ : LocalMux
    port map (
            O => \N__45968\,
            I => \N__45961\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__45965\,
            I => \N__45958\
        );

    \I__10555\ : InMux
    port map (
            O => \N__45964\,
            I => \N__45955\
        );

    \I__10554\ : Span4Mux_v
    port map (
            O => \N__45961\,
            I => \N__45952\
        );

    \I__10553\ : Span4Mux_h
    port map (
            O => \N__45958\,
            I => \N__45949\
        );

    \I__10552\ : LocalMux
    port map (
            O => \N__45955\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10551\ : Odrv4
    port map (
            O => \N__45952\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10550\ : Odrv4
    port map (
            O => \N__45949\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\
        );

    \I__10549\ : InMux
    port map (
            O => \N__45942\,
            I => \bfn_18_13_0_\
        );

    \I__10548\ : CascadeMux
    port map (
            O => \N__45939\,
            I => \N__45935\
        );

    \I__10547\ : CascadeMux
    port map (
            O => \N__45938\,
            I => \N__45932\
        );

    \I__10546\ : InMux
    port map (
            O => \N__45935\,
            I => \N__45929\
        );

    \I__10545\ : InMux
    port map (
            O => \N__45932\,
            I => \N__45926\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__45929\,
            I => \N__45920\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__45926\,
            I => \N__45920\
        );

    \I__10542\ : InMux
    port map (
            O => \N__45925\,
            I => \N__45917\
        );

    \I__10541\ : Span4Mux_v
    port map (
            O => \N__45920\,
            I => \N__45914\
        );

    \I__10540\ : LocalMux
    port map (
            O => \N__45917\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10539\ : Odrv4
    port map (
            O => \N__45914\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\
        );

    \I__10538\ : InMux
    port map (
            O => \N__45909\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_16\
        );

    \I__10537\ : CascadeMux
    port map (
            O => \N__45906\,
            I => \N__45903\
        );

    \I__10536\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45899\
        );

    \I__10535\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45896\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__45899\,
            I => \N__45890\
        );

    \I__10533\ : LocalMux
    port map (
            O => \N__45896\,
            I => \N__45890\
        );

    \I__10532\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45887\
        );

    \I__10531\ : Span4Mux_h
    port map (
            O => \N__45890\,
            I => \N__45884\
        );

    \I__10530\ : LocalMux
    port map (
            O => \N__45887\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10529\ : Odrv4
    port map (
            O => \N__45884\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\
        );

    \I__10528\ : InMux
    port map (
            O => \N__45879\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_17\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__45876\,
            I => \N__45873\
        );

    \I__10526\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45869\
        );

    \I__10525\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45866\
        );

    \I__10524\ : LocalMux
    port map (
            O => \N__45869\,
            I => \N__45860\
        );

    \I__10523\ : LocalMux
    port map (
            O => \N__45866\,
            I => \N__45860\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45865\,
            I => \N__45857\
        );

    \I__10521\ : Span4Mux_h
    port map (
            O => \N__45860\,
            I => \N__45854\
        );

    \I__10520\ : LocalMux
    port map (
            O => \N__45857\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10519\ : Odrv4
    port map (
            O => \N__45854\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45849\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_18\
        );

    \I__10517\ : CascadeMux
    port map (
            O => \N__45846\,
            I => \N__45843\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45843\,
            I => \N__45839\
        );

    \I__10515\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45836\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__45839\,
            I => \N__45830\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__45836\,
            I => \N__45830\
        );

    \I__10512\ : InMux
    port map (
            O => \N__45835\,
            I => \N__45827\
        );

    \I__10511\ : Span4Mux_h
    port map (
            O => \N__45830\,
            I => \N__45824\
        );

    \I__10510\ : LocalMux
    port map (
            O => \N__45827\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10509\ : Odrv4
    port map (
            O => \N__45824\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\
        );

    \I__10508\ : InMux
    port map (
            O => \N__45819\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_19\
        );

    \I__10507\ : CascadeMux
    port map (
            O => \N__45816\,
            I => \N__45812\
        );

    \I__10506\ : CascadeMux
    port map (
            O => \N__45815\,
            I => \N__45809\
        );

    \I__10505\ : InMux
    port map (
            O => \N__45812\,
            I => \N__45804\
        );

    \I__10504\ : InMux
    port map (
            O => \N__45809\,
            I => \N__45804\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45804\,
            I => \N__45800\
        );

    \I__10502\ : InMux
    port map (
            O => \N__45803\,
            I => \N__45797\
        );

    \I__10501\ : Span4Mux_h
    port map (
            O => \N__45800\,
            I => \N__45794\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__45797\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__10499\ : Odrv4
    port map (
            O => \N__45794\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\
        );

    \I__10498\ : InMux
    port map (
            O => \N__45789\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_3\
        );

    \I__10497\ : CascadeMux
    port map (
            O => \N__45786\,
            I => \N__45782\
        );

    \I__10496\ : CascadeMux
    port map (
            O => \N__45785\,
            I => \N__45779\
        );

    \I__10495\ : InMux
    port map (
            O => \N__45782\,
            I => \N__45774\
        );

    \I__10494\ : InMux
    port map (
            O => \N__45779\,
            I => \N__45774\
        );

    \I__10493\ : LocalMux
    port map (
            O => \N__45774\,
            I => \N__45770\
        );

    \I__10492\ : InMux
    port map (
            O => \N__45773\,
            I => \N__45767\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__45770\,
            I => \N__45764\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45767\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__10489\ : Odrv4
    port map (
            O => \N__45764\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45759\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_4\
        );

    \I__10487\ : InMux
    port map (
            O => \N__45756\,
            I => \N__45750\
        );

    \I__10486\ : InMux
    port map (
            O => \N__45755\,
            I => \N__45750\
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45746\
        );

    \I__10484\ : InMux
    port map (
            O => \N__45749\,
            I => \N__45743\
        );

    \I__10483\ : Span4Mux_h
    port map (
            O => \N__45746\,
            I => \N__45740\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__45743\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__10481\ : Odrv4
    port map (
            O => \N__45740\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\
        );

    \I__10480\ : InMux
    port map (
            O => \N__45735\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_5\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45732\,
            I => \N__45726\
        );

    \I__10478\ : InMux
    port map (
            O => \N__45731\,
            I => \N__45726\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__45726\,
            I => \N__45722\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45725\,
            I => \N__45719\
        );

    \I__10475\ : Span4Mux_h
    port map (
            O => \N__45722\,
            I => \N__45716\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45719\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10473\ : Odrv4
    port map (
            O => \N__45716\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\
        );

    \I__10472\ : InMux
    port map (
            O => \N__45711\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_6\
        );

    \I__10471\ : CascadeMux
    port map (
            O => \N__45708\,
            I => \N__45704\
        );

    \I__10470\ : CascadeMux
    port map (
            O => \N__45707\,
            I => \N__45701\
        );

    \I__10469\ : InMux
    port map (
            O => \N__45704\,
            I => \N__45698\
        );

    \I__10468\ : InMux
    port map (
            O => \N__45701\,
            I => \N__45695\
        );

    \I__10467\ : LocalMux
    port map (
            O => \N__45698\,
            I => \N__45691\
        );

    \I__10466\ : LocalMux
    port map (
            O => \N__45695\,
            I => \N__45688\
        );

    \I__10465\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45685\
        );

    \I__10464\ : Span4Mux_v
    port map (
            O => \N__45691\,
            I => \N__45682\
        );

    \I__10463\ : Span4Mux_h
    port map (
            O => \N__45688\,
            I => \N__45679\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__45685\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__45682\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10460\ : Odrv4
    port map (
            O => \N__45679\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\
        );

    \I__10459\ : InMux
    port map (
            O => \N__45672\,
            I => \bfn_18_12_0_\
        );

    \I__10458\ : CascadeMux
    port map (
            O => \N__45669\,
            I => \N__45665\
        );

    \I__10457\ : CascadeMux
    port map (
            O => \N__45668\,
            I => \N__45662\
        );

    \I__10456\ : InMux
    port map (
            O => \N__45665\,
            I => \N__45659\
        );

    \I__10455\ : InMux
    port map (
            O => \N__45662\,
            I => \N__45656\
        );

    \I__10454\ : LocalMux
    port map (
            O => \N__45659\,
            I => \N__45652\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__45656\,
            I => \N__45649\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45646\
        );

    \I__10451\ : Span4Mux_v
    port map (
            O => \N__45652\,
            I => \N__45643\
        );

    \I__10450\ : Span4Mux_h
    port map (
            O => \N__45649\,
            I => \N__45640\
        );

    \I__10449\ : LocalMux
    port map (
            O => \N__45646\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10448\ : Odrv4
    port map (
            O => \N__45643\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10447\ : Odrv4
    port map (
            O => \N__45640\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\
        );

    \I__10446\ : InMux
    port map (
            O => \N__45633\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_8\
        );

    \I__10445\ : CascadeMux
    port map (
            O => \N__45630\,
            I => \N__45627\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45627\,
            I => \N__45623\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45626\,
            I => \N__45620\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__45623\,
            I => \N__45614\
        );

    \I__10441\ : LocalMux
    port map (
            O => \N__45620\,
            I => \N__45614\
        );

    \I__10440\ : InMux
    port map (
            O => \N__45619\,
            I => \N__45611\
        );

    \I__10439\ : Span4Mux_h
    port map (
            O => \N__45614\,
            I => \N__45608\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__45611\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10437\ : Odrv4
    port map (
            O => \N__45608\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45603\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_9\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45600\,
            I => \N__45594\
        );

    \I__10434\ : InMux
    port map (
            O => \N__45599\,
            I => \N__45594\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45594\,
            I => \N__45590\
        );

    \I__10432\ : InMux
    port map (
            O => \N__45593\,
            I => \N__45587\
        );

    \I__10431\ : Span4Mux_h
    port map (
            O => \N__45590\,
            I => \N__45584\
        );

    \I__10430\ : LocalMux
    port map (
            O => \N__45587\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10429\ : Odrv4
    port map (
            O => \N__45584\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\
        );

    \I__10428\ : InMux
    port map (
            O => \N__45579\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_10\
        );

    \I__10427\ : InMux
    port map (
            O => \N__45576\,
            I => \N__45570\
        );

    \I__10426\ : InMux
    port map (
            O => \N__45575\,
            I => \N__45570\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__45570\,
            I => \N__45567\
        );

    \I__10424\ : Odrv12
    port map (
            O => \N__45567\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\
        );

    \I__10423\ : CascadeMux
    port map (
            O => \N__45564\,
            I => \N__45559\
        );

    \I__10422\ : InMux
    port map (
            O => \N__45563\,
            I => \N__45556\
        );

    \I__10421\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45551\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45559\,
            I => \N__45551\
        );

    \I__10419\ : LocalMux
    port map (
            O => \N__45556\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45551\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__10417\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45541\
        );

    \I__10416\ : InMux
    port map (
            O => \N__45545\,
            I => \N__45536\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45544\,
            I => \N__45536\
        );

    \I__10414\ : LocalMux
    port map (
            O => \N__45541\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__10413\ : LocalMux
    port map (
            O => \N__45536\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__10412\ : CascadeMux
    port map (
            O => \N__45531\,
            I => \N__45528\
        );

    \I__10411\ : InMux
    port map (
            O => \N__45528\,
            I => \N__45525\
        );

    \I__10410\ : LocalMux
    port map (
            O => \N__45525\,
            I => \N__45522\
        );

    \I__10409\ : Span4Mux_v
    port map (
            O => \N__45522\,
            I => \N__45519\
        );

    \I__10408\ : Odrv4
    port map (
            O => \N__45519\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\
        );

    \I__10407\ : CascadeMux
    port map (
            O => \N__45516\,
            I => \N__45511\
        );

    \I__10406\ : InMux
    port map (
            O => \N__45515\,
            I => \N__45508\
        );

    \I__10405\ : CascadeMux
    port map (
            O => \N__45514\,
            I => \N__45504\
        );

    \I__10404\ : InMux
    port map (
            O => \N__45511\,
            I => \N__45501\
        );

    \I__10403\ : LocalMux
    port map (
            O => \N__45508\,
            I => \N__45498\
        );

    \I__10402\ : InMux
    port map (
            O => \N__45507\,
            I => \N__45493\
        );

    \I__10401\ : InMux
    port map (
            O => \N__45504\,
            I => \N__45493\
        );

    \I__10400\ : LocalMux
    port map (
            O => \N__45501\,
            I => \N__45490\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__45498\,
            I => \N__45487\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45493\,
            I => \N__45484\
        );

    \I__10397\ : Span4Mux_h
    port map (
            O => \N__45490\,
            I => \N__45481\
        );

    \I__10396\ : Odrv4
    port map (
            O => \N__45487\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__45484\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10394\ : Odrv4
    port map (
            O => \N__45481\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\
        );

    \I__10393\ : InMux
    port map (
            O => \N__45474\,
            I => \N__45471\
        );

    \I__10392\ : LocalMux
    port map (
            O => \N__45471\,
            I => \N__45468\
        );

    \I__10391\ : Span4Mux_h
    port map (
            O => \N__45468\,
            I => \N__45464\
        );

    \I__10390\ : InMux
    port map (
            O => \N__45467\,
            I => \N__45461\
        );

    \I__10389\ : Odrv4
    port map (
            O => \N__45464\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__45461\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21\
        );

    \I__10387\ : CascadeMux
    port map (
            O => \N__45456\,
            I => \N__45452\
        );

    \I__10386\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45447\
        );

    \I__10385\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45447\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45447\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\
        );

    \I__10383\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45436\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45436\
        );

    \I__10381\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45433\
        );

    \I__10380\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45430\
        );

    \I__10379\ : LocalMux
    port map (
            O => \N__45436\,
            I => \N__45425\
        );

    \I__10378\ : LocalMux
    port map (
            O => \N__45433\,
            I => \N__45425\
        );

    \I__10377\ : LocalMux
    port map (
            O => \N__45430\,
            I => \N__45422\
        );

    \I__10376\ : Span4Mux_v
    port map (
            O => \N__45425\,
            I => \N__45419\
        );

    \I__10375\ : Odrv12
    port map (
            O => \N__45422\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45419\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\
        );

    \I__10373\ : InMux
    port map (
            O => \N__45414\,
            I => \N__45411\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45411\,
            I => \N__45408\
        );

    \I__10371\ : Span12Mux_s10_v
    port map (
            O => \N__45408\,
            I => \N__45404\
        );

    \I__10370\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45401\
        );

    \I__10369\ : Odrv12
    port map (
            O => \N__45404\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__45401\,
            I => \elapsed_time_ns_1_RNII43T9_0_6\
        );

    \I__10367\ : InMux
    port map (
            O => \N__45396\,
            I => \N__45393\
        );

    \I__10366\ : LocalMux
    port map (
            O => \N__45393\,
            I => \N__45390\
        );

    \I__10365\ : Span4Mux_v
    port map (
            O => \N__45390\,
            I => \N__45387\
        );

    \I__10364\ : Odrv4
    port map (
            O => \N__45387\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\
        );

    \I__10363\ : InMux
    port map (
            O => \N__45384\,
            I => \N__45380\
        );

    \I__10362\ : InMux
    port map (
            O => \N__45383\,
            I => \N__45377\
        );

    \I__10361\ : LocalMux
    port map (
            O => \N__45380\,
            I => \N__45373\
        );

    \I__10360\ : LocalMux
    port map (
            O => \N__45377\,
            I => \N__45370\
        );

    \I__10359\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45367\
        );

    \I__10358\ : Span4Mux_h
    port map (
            O => \N__45373\,
            I => \N__45364\
        );

    \I__10357\ : Span4Mux_h
    port map (
            O => \N__45370\,
            I => \N__45361\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__45367\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__10355\ : Odrv4
    port map (
            O => \N__45364\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__10354\ : Odrv4
    port map (
            O => \N__45361\,
            I => \elapsed_time_ns_1_RNIJ53T9_0_7\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45354\,
            I => \N__45349\
        );

    \I__10352\ : InMux
    port map (
            O => \N__45353\,
            I => \N__45346\
        );

    \I__10351\ : InMux
    port map (
            O => \N__45352\,
            I => \N__45343\
        );

    \I__10350\ : LocalMux
    port map (
            O => \N__45349\,
            I => \N__45337\
        );

    \I__10349\ : LocalMux
    port map (
            O => \N__45346\,
            I => \N__45337\
        );

    \I__10348\ : LocalMux
    port map (
            O => \N__45343\,
            I => \N__45334\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45342\,
            I => \N__45331\
        );

    \I__10346\ : Span4Mux_v
    port map (
            O => \N__45337\,
            I => \N__45328\
        );

    \I__10345\ : Odrv4
    port map (
            O => \N__45334\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__45331\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__10343\ : Odrv4
    port map (
            O => \N__45328\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\
        );

    \I__10342\ : InMux
    port map (
            O => \N__45321\,
            I => \N__45318\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__45318\,
            I => \N__45315\
        );

    \I__10340\ : Span4Mux_v
    port map (
            O => \N__45315\,
            I => \N__45312\
        );

    \I__10339\ : Odrv4
    port map (
            O => \N__45312\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\
        );

    \I__10338\ : InMux
    port map (
            O => \N__45309\,
            I => \bfn_18_11_0_\
        );

    \I__10337\ : CascadeMux
    port map (
            O => \N__45306\,
            I => \N__45302\
        );

    \I__10336\ : InMux
    port map (
            O => \N__45305\,
            I => \N__45299\
        );

    \I__10335\ : InMux
    port map (
            O => \N__45302\,
            I => \N__45296\
        );

    \I__10334\ : LocalMux
    port map (
            O => \N__45299\,
            I => \N__45292\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__45296\,
            I => \N__45289\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45295\,
            I => \N__45286\
        );

    \I__10331\ : Span4Mux_v
    port map (
            O => \N__45292\,
            I => \N__45281\
        );

    \I__10330\ : Span4Mux_v
    port map (
            O => \N__45289\,
            I => \N__45281\
        );

    \I__10329\ : LocalMux
    port map (
            O => \N__45286\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__10328\ : Odrv4
    port map (
            O => \N__45281\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\
        );

    \I__10327\ : InMux
    port map (
            O => \N__45276\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_0\
        );

    \I__10326\ : InMux
    port map (
            O => \N__45273\,
            I => \N__45267\
        );

    \I__10325\ : InMux
    port map (
            O => \N__45272\,
            I => \N__45267\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__45267\,
            I => \N__45263\
        );

    \I__10323\ : InMux
    port map (
            O => \N__45266\,
            I => \N__45260\
        );

    \I__10322\ : Span4Mux_h
    port map (
            O => \N__45263\,
            I => \N__45257\
        );

    \I__10321\ : LocalMux
    port map (
            O => \N__45260\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__10320\ : Odrv4
    port map (
            O => \N__45257\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\
        );

    \I__10319\ : InMux
    port map (
            O => \N__45252\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_1\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45249\,
            I => \N__45243\
        );

    \I__10317\ : InMux
    port map (
            O => \N__45248\,
            I => \N__45243\
        );

    \I__10316\ : LocalMux
    port map (
            O => \N__45243\,
            I => \N__45239\
        );

    \I__10315\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45236\
        );

    \I__10314\ : Span4Mux_h
    port map (
            O => \N__45239\,
            I => \N__45233\
        );

    \I__10313\ : LocalMux
    port map (
            O => \N__45236\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__10312\ : Odrv4
    port map (
            O => \N__45233\,
            I => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\
        );

    \I__10311\ : InMux
    port map (
            O => \N__45228\,
            I => \delay_measurement_inst.delay_hc_timer.counter_cry_2\
        );

    \I__10310\ : InMux
    port map (
            O => \N__45225\,
            I => \N__45222\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__45222\,
            I => \N__45219\
        );

    \I__10308\ : Odrv4
    port map (
            O => \N__45219\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45216\,
            I => \N__45213\
        );

    \I__10306\ : LocalMux
    port map (
            O => \N__45213\,
            I => \N__45209\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45212\,
            I => \N__45205\
        );

    \I__10304\ : Span4Mux_h
    port map (
            O => \N__45209\,
            I => \N__45202\
        );

    \I__10303\ : InMux
    port map (
            O => \N__45208\,
            I => \N__45199\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__45205\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__10301\ : Odrv4
    port map (
            O => \N__45202\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45199\,
            I => \elapsed_time_ns_1_RNI24CN9_0_15\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45192\,
            I => \N__45187\
        );

    \I__10298\ : InMux
    port map (
            O => \N__45191\,
            I => \N__45184\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45190\,
            I => \N__45181\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45187\,
            I => \N__45178\
        );

    \I__10295\ : LocalMux
    port map (
            O => \N__45184\,
            I => \N__45173\
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__45181\,
            I => \N__45173\
        );

    \I__10293\ : Span4Mux_v
    port map (
            O => \N__45178\,
            I => \N__45167\
        );

    \I__10292\ : Span4Mux_v
    port map (
            O => \N__45173\,
            I => \N__45167\
        );

    \I__10291\ : InMux
    port map (
            O => \N__45172\,
            I => \N__45164\
        );

    \I__10290\ : Odrv4
    port map (
            O => \N__45167\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10289\ : LocalMux
    port map (
            O => \N__45164\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\
        );

    \I__10288\ : CascadeMux
    port map (
            O => \N__45159\,
            I => \N__45156\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45156\,
            I => \N__45153\
        );

    \I__10286\ : LocalMux
    port map (
            O => \N__45153\,
            I => \N__45150\
        );

    \I__10285\ : Odrv4
    port map (
            O => \N__45150\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\
        );

    \I__10284\ : InMux
    port map (
            O => \N__45147\,
            I => \N__45143\
        );

    \I__10283\ : InMux
    port map (
            O => \N__45146\,
            I => \N__45140\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__45143\,
            I => \N__45136\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__45140\,
            I => \N__45133\
        );

    \I__10280\ : InMux
    port map (
            O => \N__45139\,
            I => \N__45130\
        );

    \I__10279\ : Span4Mux_v
    port map (
            O => \N__45136\,
            I => \N__45127\
        );

    \I__10278\ : Span4Mux_h
    port map (
            O => \N__45133\,
            I => \N__45124\
        );

    \I__10277\ : LocalMux
    port map (
            O => \N__45130\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10276\ : Odrv4
    port map (
            O => \N__45127\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10275\ : Odrv4
    port map (
            O => \N__45124\,
            I => \elapsed_time_ns_1_RNIDV2T9_0_1\
        );

    \I__10274\ : InMux
    port map (
            O => \N__45117\,
            I => \N__45114\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__45114\,
            I => \N__45111\
        );

    \I__10272\ : Span4Mux_h
    port map (
            O => \N__45111\,
            I => \N__45108\
        );

    \I__10271\ : Odrv4
    port map (
            O => \N__45108\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\
        );

    \I__10270\ : InMux
    port map (
            O => \N__45105\,
            I => \N__45102\
        );

    \I__10269\ : LocalMux
    port map (
            O => \N__45102\,
            I => \N__45099\
        );

    \I__10268\ : Odrv4
    port map (
            O => \N__45099\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt24\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45096\,
            I => \N__45090\
        );

    \I__10266\ : InMux
    port map (
            O => \N__45095\,
            I => \N__45090\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__45090\,
            I => \N__45087\
        );

    \I__10264\ : Odrv4
    port map (
            O => \N__45087\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\
        );

    \I__10263\ : CascadeMux
    port map (
            O => \N__45084\,
            I => \N__45079\
        );

    \I__10262\ : InMux
    port map (
            O => \N__45083\,
            I => \N__45076\
        );

    \I__10261\ : InMux
    port map (
            O => \N__45082\,
            I => \N__45071\
        );

    \I__10260\ : InMux
    port map (
            O => \N__45079\,
            I => \N__45071\
        );

    \I__10259\ : LocalMux
    port map (
            O => \N__45076\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__10258\ : LocalMux
    port map (
            O => \N__45071\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__10257\ : InMux
    port map (
            O => \N__45066\,
            I => \N__45061\
        );

    \I__10256\ : InMux
    port map (
            O => \N__45065\,
            I => \N__45056\
        );

    \I__10255\ : InMux
    port map (
            O => \N__45064\,
            I => \N__45056\
        );

    \I__10254\ : LocalMux
    port map (
            O => \N__45061\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10253\ : LocalMux
    port map (
            O => \N__45056\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__10252\ : CascadeMux
    port map (
            O => \N__45051\,
            I => \N__45048\
        );

    \I__10251\ : InMux
    port map (
            O => \N__45048\,
            I => \N__45045\
        );

    \I__10250\ : LocalMux
    port map (
            O => \N__45045\,
            I => \N__45042\
        );

    \I__10249\ : Odrv12
    port map (
            O => \N__45042\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\
        );

    \I__10248\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45035\
        );

    \I__10247\ : InMux
    port map (
            O => \N__45038\,
            I => \N__45031\
        );

    \I__10246\ : LocalMux
    port map (
            O => \N__45035\,
            I => \N__45028\
        );

    \I__10245\ : InMux
    port map (
            O => \N__45034\,
            I => \N__45025\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__45031\,
            I => \N__45020\
        );

    \I__10243\ : Span4Mux_v
    port map (
            O => \N__45028\,
            I => \N__45020\
        );

    \I__10242\ : LocalMux
    port map (
            O => \N__45025\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__10241\ : Odrv4
    port map (
            O => \N__45020\,
            I => \elapsed_time_ns_1_RNI36DN9_0_25\
        );

    \I__10240\ : InMux
    port map (
            O => \N__45015\,
            I => \N__45010\
        );

    \I__10239\ : InMux
    port map (
            O => \N__45014\,
            I => \N__45007\
        );

    \I__10238\ : InMux
    port map (
            O => \N__45013\,
            I => \N__45004\
        );

    \I__10237\ : LocalMux
    port map (
            O => \N__45010\,
            I => \N__45000\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__45007\,
            I => \N__44997\
        );

    \I__10235\ : LocalMux
    port map (
            O => \N__45004\,
            I => \N__44994\
        );

    \I__10234\ : InMux
    port map (
            O => \N__45003\,
            I => \N__44991\
        );

    \I__10233\ : Span4Mux_v
    port map (
            O => \N__45000\,
            I => \N__44988\
        );

    \I__10232\ : Span12Mux_s11_v
    port map (
            O => \N__44997\,
            I => \N__44985\
        );

    \I__10231\ : Span4Mux_v
    port map (
            O => \N__44994\,
            I => \N__44980\
        );

    \I__10230\ : LocalMux
    port map (
            O => \N__44991\,
            I => \N__44980\
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__44988\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10228\ : Odrv12
    port map (
            O => \N__44985\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10227\ : Odrv4
    port map (
            O => \N__44980\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\
        );

    \I__10226\ : CascadeMux
    port map (
            O => \N__44973\,
            I => \N__44969\
        );

    \I__10225\ : InMux
    port map (
            O => \N__44972\,
            I => \N__44964\
        );

    \I__10224\ : InMux
    port map (
            O => \N__44969\,
            I => \N__44964\
        );

    \I__10223\ : LocalMux
    port map (
            O => \N__44964\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\
        );

    \I__10222\ : CascadeMux
    port map (
            O => \N__44961\,
            I => \N__44958\
        );

    \I__10221\ : InMux
    port map (
            O => \N__44958\,
            I => \N__44955\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__44955\,
            I => \N__44952\
        );

    \I__10219\ : Odrv12
    port map (
            O => \N__44952\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\
        );

    \I__10218\ : CascadeMux
    port map (
            O => \N__44949\,
            I => \N__44944\
        );

    \I__10217\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44941\
        );

    \I__10216\ : InMux
    port map (
            O => \N__44947\,
            I => \N__44938\
        );

    \I__10215\ : InMux
    port map (
            O => \N__44944\,
            I => \N__44935\
        );

    \I__10214\ : LocalMux
    port map (
            O => \N__44941\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__44938\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__10212\ : LocalMux
    port map (
            O => \N__44935\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__10211\ : InMux
    port map (
            O => \N__44928\,
            I => \N__44922\
        );

    \I__10210\ : InMux
    port map (
            O => \N__44927\,
            I => \N__44922\
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__44922\,
            I => \N__44919\
        );

    \I__10208\ : Odrv4
    port map (
            O => \N__44919\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\
        );

    \I__10207\ : InMux
    port map (
            O => \N__44916\,
            I => \N__44911\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44915\,
            I => \N__44908\
        );

    \I__10205\ : InMux
    port map (
            O => \N__44914\,
            I => \N__44905\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__44911\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__44908\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__44905\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__10201\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44895\
        );

    \I__10200\ : LocalMux
    port map (
            O => \N__44895\,
            I => \N__44892\
        );

    \I__10199\ : Odrv4
    port map (
            O => \N__44892\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt26\
        );

    \I__10198\ : InMux
    port map (
            O => \N__44889\,
            I => \N__44886\
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44886\,
            I => \N__44883\
        );

    \I__10196\ : Span4Mux_v
    port map (
            O => \N__44883\,
            I => \N__44880\
        );

    \I__10195\ : Odrv4
    port map (
            O => \N__44880\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt20\
        );

    \I__10194\ : InMux
    port map (
            O => \N__44877\,
            I => \current_shift_inst.timer_s1.counter_cry_27\
        );

    \I__10193\ : InMux
    port map (
            O => \N__44874\,
            I => \N__44854\
        );

    \I__10192\ : InMux
    port map (
            O => \N__44873\,
            I => \N__44854\
        );

    \I__10191\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44854\
        );

    \I__10190\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44854\
        );

    \I__10189\ : InMux
    port map (
            O => \N__44870\,
            I => \N__44837\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44869\,
            I => \N__44837\
        );

    \I__10187\ : InMux
    port map (
            O => \N__44868\,
            I => \N__44837\
        );

    \I__10186\ : InMux
    port map (
            O => \N__44867\,
            I => \N__44837\
        );

    \I__10185\ : InMux
    port map (
            O => \N__44866\,
            I => \N__44828\
        );

    \I__10184\ : InMux
    port map (
            O => \N__44865\,
            I => \N__44828\
        );

    \I__10183\ : InMux
    port map (
            O => \N__44864\,
            I => \N__44828\
        );

    \I__10182\ : InMux
    port map (
            O => \N__44863\,
            I => \N__44828\
        );

    \I__10181\ : LocalMux
    port map (
            O => \N__44854\,
            I => \N__44815\
        );

    \I__10180\ : InMux
    port map (
            O => \N__44853\,
            I => \N__44806\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44852\,
            I => \N__44806\
        );

    \I__10178\ : InMux
    port map (
            O => \N__44851\,
            I => \N__44806\
        );

    \I__10177\ : InMux
    port map (
            O => \N__44850\,
            I => \N__44806\
        );

    \I__10176\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44797\
        );

    \I__10175\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44797\
        );

    \I__10174\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44797\
        );

    \I__10173\ : InMux
    port map (
            O => \N__44846\,
            I => \N__44797\
        );

    \I__10172\ : LocalMux
    port map (
            O => \N__44837\,
            I => \N__44792\
        );

    \I__10171\ : LocalMux
    port map (
            O => \N__44828\,
            I => \N__44792\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44827\,
            I => \N__44787\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44826\,
            I => \N__44787\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44825\,
            I => \N__44778\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44824\,
            I => \N__44778\
        );

    \I__10166\ : InMux
    port map (
            O => \N__44823\,
            I => \N__44778\
        );

    \I__10165\ : InMux
    port map (
            O => \N__44822\,
            I => \N__44778\
        );

    \I__10164\ : InMux
    port map (
            O => \N__44821\,
            I => \N__44769\
        );

    \I__10163\ : InMux
    port map (
            O => \N__44820\,
            I => \N__44769\
        );

    \I__10162\ : InMux
    port map (
            O => \N__44819\,
            I => \N__44769\
        );

    \I__10161\ : InMux
    port map (
            O => \N__44818\,
            I => \N__44769\
        );

    \I__10160\ : Span4Mux_v
    port map (
            O => \N__44815\,
            I => \N__44762\
        );

    \I__10159\ : LocalMux
    port map (
            O => \N__44806\,
            I => \N__44762\
        );

    \I__10158\ : LocalMux
    port map (
            O => \N__44797\,
            I => \N__44762\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__44792\,
            I => \N__44755\
        );

    \I__10156\ : LocalMux
    port map (
            O => \N__44787\,
            I => \N__44755\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__44778\,
            I => \N__44755\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__44769\,
            I => \N__44752\
        );

    \I__10153\ : Span4Mux_h
    port map (
            O => \N__44762\,
            I => \N__44749\
        );

    \I__10152\ : Span4Mux_h
    port map (
            O => \N__44755\,
            I => \N__44746\
        );

    \I__10151\ : Odrv12
    port map (
            O => \N__44752\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10150\ : Odrv4
    port map (
            O => \N__44749\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10149\ : Odrv4
    port map (
            O => \N__44746\,
            I => \current_shift_inst.timer_s1.running_i\
        );

    \I__10148\ : InMux
    port map (
            O => \N__44739\,
            I => \current_shift_inst.timer_s1.counter_cry_28\
        );

    \I__10147\ : CascadeMux
    port map (
            O => \N__44736\,
            I => \N__44733\
        );

    \I__10146\ : InMux
    port map (
            O => \N__44733\,
            I => \N__44730\
        );

    \I__10145\ : LocalMux
    port map (
            O => \N__44730\,
            I => \N__44726\
        );

    \I__10144\ : InMux
    port map (
            O => \N__44729\,
            I => \N__44723\
        );

    \I__10143\ : Span4Mux_h
    port map (
            O => \N__44726\,
            I => \N__44720\
        );

    \I__10142\ : LocalMux
    port map (
            O => \N__44723\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10141\ : Odrv4
    port map (
            O => \N__44720\,
            I => \current_shift_inst.timer_s1.counterZ0Z_29\
        );

    \I__10140\ : CEMux
    port map (
            O => \N__44715\,
            I => \N__44710\
        );

    \I__10139\ : CEMux
    port map (
            O => \N__44714\,
            I => \N__44707\
        );

    \I__10138\ : CEMux
    port map (
            O => \N__44713\,
            I => \N__44703\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__44710\,
            I => \N__44700\
        );

    \I__10136\ : LocalMux
    port map (
            O => \N__44707\,
            I => \N__44697\
        );

    \I__10135\ : CEMux
    port map (
            O => \N__44706\,
            I => \N__44694\
        );

    \I__10134\ : LocalMux
    port map (
            O => \N__44703\,
            I => \N__44691\
        );

    \I__10133\ : Span4Mux_v
    port map (
            O => \N__44700\,
            I => \N__44686\
        );

    \I__10132\ : Span4Mux_h
    port map (
            O => \N__44697\,
            I => \N__44686\
        );

    \I__10131\ : LocalMux
    port map (
            O => \N__44694\,
            I => \N__44683\
        );

    \I__10130\ : Span4Mux_h
    port map (
            O => \N__44691\,
            I => \N__44680\
        );

    \I__10129\ : Span4Mux_h
    port map (
            O => \N__44686\,
            I => \N__44677\
        );

    \I__10128\ : Span4Mux_h
    port map (
            O => \N__44683\,
            I => \N__44674\
        );

    \I__10127\ : Odrv4
    port map (
            O => \N__44680\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__10126\ : Odrv4
    port map (
            O => \N__44677\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__10125\ : Odrv4
    port map (
            O => \N__44674\,
            I => \current_shift_inst.timer_s1.N_162_i\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44664\
        );

    \I__10123\ : LocalMux
    port map (
            O => \N__44664\,
            I => \N__44658\
        );

    \I__10122\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44655\
        );

    \I__10121\ : InMux
    port map (
            O => \N__44662\,
            I => \N__44650\
        );

    \I__10120\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44650\
        );

    \I__10119\ : Span4Mux_v
    port map (
            O => \N__44658\,
            I => \N__44647\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__44655\,
            I => \N__44644\
        );

    \I__10117\ : LocalMux
    port map (
            O => \N__44650\,
            I => \N__44641\
        );

    \I__10116\ : Span4Mux_v
    port map (
            O => \N__44647\,
            I => \N__44636\
        );

    \I__10115\ : Span4Mux_v
    port map (
            O => \N__44644\,
            I => \N__44636\
        );

    \I__10114\ : Odrv4
    port map (
            O => \N__44641\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10113\ : Odrv4
    port map (
            O => \N__44636\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44628\
        );

    \I__10111\ : LocalMux
    port map (
            O => \N__44628\,
            I => \N__44625\
        );

    \I__10110\ : Span4Mux_h
    port map (
            O => \N__44625\,
            I => \N__44621\
        );

    \I__10109\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44618\
        );

    \I__10108\ : Odrv4
    port map (
            O => \N__44621\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__10107\ : LocalMux
    port map (
            O => \N__44618\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20\
        );

    \I__10106\ : InMux
    port map (
            O => \N__44613\,
            I => \N__44608\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44612\,
            I => \N__44605\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44611\,
            I => \N__44602\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__44608\,
            I => \N__44599\
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44605\,
            I => \N__44596\
        );

    \I__10101\ : LocalMux
    port map (
            O => \N__44602\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10100\ : Odrv4
    port map (
            O => \N__44599\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10099\ : Odrv4
    port map (
            O => \N__44596\,
            I => \elapsed_time_ns_1_RNI46CN9_0_17\
        );

    \I__10098\ : InMux
    port map (
            O => \N__44589\,
            I => \N__44585\
        );

    \I__10097\ : InMux
    port map (
            O => \N__44588\,
            I => \N__44581\
        );

    \I__10096\ : LocalMux
    port map (
            O => \N__44585\,
            I => \N__44578\
        );

    \I__10095\ : InMux
    port map (
            O => \N__44584\,
            I => \N__44575\
        );

    \I__10094\ : LocalMux
    port map (
            O => \N__44581\,
            I => \N__44571\
        );

    \I__10093\ : Span4Mux_v
    port map (
            O => \N__44578\,
            I => \N__44566\
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__44575\,
            I => \N__44566\
        );

    \I__10091\ : InMux
    port map (
            O => \N__44574\,
            I => \N__44563\
        );

    \I__10090\ : Span12Mux_s10_v
    port map (
            O => \N__44571\,
            I => \N__44560\
        );

    \I__10089\ : Span4Mux_v
    port map (
            O => \N__44566\,
            I => \N__44557\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__44563\,
            I => \N__44554\
        );

    \I__10087\ : Odrv12
    port map (
            O => \N__44560\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10086\ : Odrv4
    port map (
            O => \N__44557\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10085\ : Odrv4
    port map (
            O => \N__44554\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44542\
        );

    \I__10083\ : InMux
    port map (
            O => \N__44546\,
            I => \N__44537\
        );

    \I__10082\ : InMux
    port map (
            O => \N__44545\,
            I => \N__44537\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__44542\,
            I => \N__44534\
        );

    \I__10080\ : LocalMux
    port map (
            O => \N__44537\,
            I => \N__44531\
        );

    \I__10079\ : Span4Mux_h
    port map (
            O => \N__44534\,
            I => \N__44525\
        );

    \I__10078\ : Span4Mux_h
    port map (
            O => \N__44531\,
            I => \N__44525\
        );

    \I__10077\ : InMux
    port map (
            O => \N__44530\,
            I => \N__44522\
        );

    \I__10076\ : Odrv4
    port map (
            O => \N__44525\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__44522\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\
        );

    \I__10074\ : InMux
    port map (
            O => \N__44517\,
            I => \N__44514\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__44514\,
            I => \N__44510\
        );

    \I__10072\ : InMux
    port map (
            O => \N__44513\,
            I => \N__44507\
        );

    \I__10071\ : Odrv4
    port map (
            O => \N__44510\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10070\ : LocalMux
    port map (
            O => \N__44507\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14\
        );

    \I__10069\ : InMux
    port map (
            O => \N__44502\,
            I => \N__44499\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44499\,
            I => \N__44496\
        );

    \I__10067\ : Span4Mux_h
    port map (
            O => \N__44496\,
            I => \N__44493\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__44493\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\
        );

    \I__10065\ : InMux
    port map (
            O => \N__44490\,
            I => \N__44487\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__44487\,
            I => \N__44484\
        );

    \I__10063\ : Span4Mux_v
    port map (
            O => \N__44484\,
            I => \N__44481\
        );

    \I__10062\ : Odrv4
    port map (
            O => \N__44481\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt16\
        );

    \I__10061\ : CascadeMux
    port map (
            O => \N__44478\,
            I => \N__44473\
        );

    \I__10060\ : InMux
    port map (
            O => \N__44477\,
            I => \N__44470\
        );

    \I__10059\ : InMux
    port map (
            O => \N__44476\,
            I => \N__44465\
        );

    \I__10058\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44465\
        );

    \I__10057\ : LocalMux
    port map (
            O => \N__44470\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__44465\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__10055\ : CascadeMux
    port map (
            O => \N__44460\,
            I => \N__44455\
        );

    \I__10054\ : InMux
    port map (
            O => \N__44459\,
            I => \N__44452\
        );

    \I__10053\ : InMux
    port map (
            O => \N__44458\,
            I => \N__44447\
        );

    \I__10052\ : InMux
    port map (
            O => \N__44455\,
            I => \N__44447\
        );

    \I__10051\ : LocalMux
    port map (
            O => \N__44452\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__44447\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__10049\ : InMux
    port map (
            O => \N__44442\,
            I => \N__44436\
        );

    \I__10048\ : InMux
    port map (
            O => \N__44441\,
            I => \N__44436\
        );

    \I__10047\ : LocalMux
    port map (
            O => \N__44436\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\
        );

    \I__10046\ : CascadeMux
    port map (
            O => \N__44433\,
            I => \N__44430\
        );

    \I__10045\ : InMux
    port map (
            O => \N__44430\,
            I => \N__44427\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__44427\,
            I => \N__44424\
        );

    \I__10043\ : Span4Mux_h
    port map (
            O => \N__44424\,
            I => \N__44421\
        );

    \I__10042\ : Odrv4
    port map (
            O => \N__44421\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\
        );

    \I__10041\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44413\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44417\,
            I => \N__44408\
        );

    \I__10039\ : InMux
    port map (
            O => \N__44416\,
            I => \N__44408\
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44413\,
            I => \N__44404\
        );

    \I__10037\ : LocalMux
    port map (
            O => \N__44408\,
            I => \N__44401\
        );

    \I__10036\ : CascadeMux
    port map (
            O => \N__44407\,
            I => \N__44398\
        );

    \I__10035\ : Span4Mux_v
    port map (
            O => \N__44404\,
            I => \N__44395\
        );

    \I__10034\ : Span4Mux_h
    port map (
            O => \N__44401\,
            I => \N__44392\
        );

    \I__10033\ : InMux
    port map (
            O => \N__44398\,
            I => \N__44389\
        );

    \I__10032\ : Odrv4
    port map (
            O => \N__44395\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10031\ : Odrv4
    port map (
            O => \N__44392\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10030\ : LocalMux
    port map (
            O => \N__44389\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\
        );

    \I__10029\ : InMux
    port map (
            O => \N__44382\,
            I => \N__44379\
        );

    \I__10028\ : LocalMux
    port map (
            O => \N__44379\,
            I => \N__44376\
        );

    \I__10027\ : Span4Mux_h
    port map (
            O => \N__44376\,
            I => \N__44372\
        );

    \I__10026\ : InMux
    port map (
            O => \N__44375\,
            I => \N__44369\
        );

    \I__10025\ : Odrv4
    port map (
            O => \N__44372\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__10024\ : LocalMux
    port map (
            O => \N__44369\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16\
        );

    \I__10023\ : InMux
    port map (
            O => \N__44364\,
            I => \N__44358\
        );

    \I__10022\ : InMux
    port map (
            O => \N__44363\,
            I => \N__44358\
        );

    \I__10021\ : LocalMux
    port map (
            O => \N__44358\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\
        );

    \I__10020\ : InMux
    port map (
            O => \N__44355\,
            I => \N__44351\
        );

    \I__10019\ : InMux
    port map (
            O => \N__44354\,
            I => \N__44348\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__44351\,
            I => \N__44344\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__44348\,
            I => \N__44341\
        );

    \I__10016\ : InMux
    port map (
            O => \N__44347\,
            I => \N__44338\
        );

    \I__10015\ : Span4Mux_v
    port map (
            O => \N__44344\,
            I => \N__44335\
        );

    \I__10014\ : Span4Mux_v
    port map (
            O => \N__44341\,
            I => \N__44332\
        );

    \I__10013\ : LocalMux
    port map (
            O => \N__44338\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__10012\ : Odrv4
    port map (
            O => \N__44335\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__44332\,
            I => \elapsed_time_ns_1_RNI02CN9_0_13\
        );

    \I__10010\ : InMux
    port map (
            O => \N__44325\,
            I => \N__44322\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__44322\,
            I => \N__44317\
        );

    \I__10008\ : InMux
    port map (
            O => \N__44321\,
            I => \N__44314\
        );

    \I__10007\ : InMux
    port map (
            O => \N__44320\,
            I => \N__44311\
        );

    \I__10006\ : Span4Mux_h
    port map (
            O => \N__44317\,
            I => \N__44307\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__44314\,
            I => \N__44304\
        );

    \I__10004\ : LocalMux
    port map (
            O => \N__44311\,
            I => \N__44301\
        );

    \I__10003\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44298\
        );

    \I__10002\ : Odrv4
    port map (
            O => \N__44307\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10001\ : Odrv12
    port map (
            O => \N__44304\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__10000\ : Odrv4
    port map (
            O => \N__44301\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__44298\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\
        );

    \I__9998\ : CascadeMux
    port map (
            O => \N__44289\,
            I => \N__44285\
        );

    \I__9997\ : CascadeMux
    port map (
            O => \N__44288\,
            I => \N__44282\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44285\,
            I => \N__44277\
        );

    \I__9995\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44277\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44277\,
            I => \N__44273\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44276\,
            I => \N__44270\
        );

    \I__9992\ : Span4Mux_h
    port map (
            O => \N__44273\,
            I => \N__44267\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__44270\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9990\ : Odrv4
    port map (
            O => \N__44267\,
            I => \current_shift_inst.timer_s1.counterZ0Z_20\
        );

    \I__9989\ : InMux
    port map (
            O => \N__44262\,
            I => \current_shift_inst.timer_s1.counter_cry_19\
        );

    \I__9988\ : CascadeMux
    port map (
            O => \N__44259\,
            I => \N__44255\
        );

    \I__9987\ : CascadeMux
    port map (
            O => \N__44258\,
            I => \N__44252\
        );

    \I__9986\ : InMux
    port map (
            O => \N__44255\,
            I => \N__44247\
        );

    \I__9985\ : InMux
    port map (
            O => \N__44252\,
            I => \N__44247\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44247\,
            I => \N__44243\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44246\,
            I => \N__44240\
        );

    \I__9982\ : Span4Mux_v
    port map (
            O => \N__44243\,
            I => \N__44237\
        );

    \I__9981\ : LocalMux
    port map (
            O => \N__44240\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9980\ : Odrv4
    port map (
            O => \N__44237\,
            I => \current_shift_inst.timer_s1.counterZ0Z_21\
        );

    \I__9979\ : InMux
    port map (
            O => \N__44232\,
            I => \current_shift_inst.timer_s1.counter_cry_20\
        );

    \I__9978\ : InMux
    port map (
            O => \N__44229\,
            I => \N__44223\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44228\,
            I => \N__44223\
        );

    \I__9976\ : LocalMux
    port map (
            O => \N__44223\,
            I => \N__44219\
        );

    \I__9975\ : InMux
    port map (
            O => \N__44222\,
            I => \N__44216\
        );

    \I__9974\ : Span4Mux_v
    port map (
            O => \N__44219\,
            I => \N__44213\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__44216\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9972\ : Odrv4
    port map (
            O => \N__44213\,
            I => \current_shift_inst.timer_s1.counterZ0Z_22\
        );

    \I__9971\ : InMux
    port map (
            O => \N__44208\,
            I => \current_shift_inst.timer_s1.counter_cry_21\
        );

    \I__9970\ : CascadeMux
    port map (
            O => \N__44205\,
            I => \N__44202\
        );

    \I__9969\ : InMux
    port map (
            O => \N__44202\,
            I => \N__44198\
        );

    \I__9968\ : InMux
    port map (
            O => \N__44201\,
            I => \N__44195\
        );

    \I__9967\ : LocalMux
    port map (
            O => \N__44198\,
            I => \N__44189\
        );

    \I__9966\ : LocalMux
    port map (
            O => \N__44195\,
            I => \N__44189\
        );

    \I__9965\ : InMux
    port map (
            O => \N__44194\,
            I => \N__44186\
        );

    \I__9964\ : Span4Mux_v
    port map (
            O => \N__44189\,
            I => \N__44183\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__44186\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__44183\,
            I => \current_shift_inst.timer_s1.counterZ0Z_23\
        );

    \I__9961\ : InMux
    port map (
            O => \N__44178\,
            I => \current_shift_inst.timer_s1.counter_cry_22\
        );

    \I__9960\ : CascadeMux
    port map (
            O => \N__44175\,
            I => \N__44171\
        );

    \I__9959\ : CascadeMux
    port map (
            O => \N__44174\,
            I => \N__44168\
        );

    \I__9958\ : InMux
    port map (
            O => \N__44171\,
            I => \N__44165\
        );

    \I__9957\ : InMux
    port map (
            O => \N__44168\,
            I => \N__44162\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__44165\,
            I => \N__44156\
        );

    \I__9955\ : LocalMux
    port map (
            O => \N__44162\,
            I => \N__44156\
        );

    \I__9954\ : InMux
    port map (
            O => \N__44161\,
            I => \N__44153\
        );

    \I__9953\ : Sp12to4
    port map (
            O => \N__44156\,
            I => \N__44150\
        );

    \I__9952\ : LocalMux
    port map (
            O => \N__44153\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9951\ : Odrv12
    port map (
            O => \N__44150\,
            I => \current_shift_inst.timer_s1.counterZ0Z_24\
        );

    \I__9950\ : InMux
    port map (
            O => \N__44145\,
            I => \bfn_17_26_0_\
        );

    \I__9949\ : CascadeMux
    port map (
            O => \N__44142\,
            I => \N__44139\
        );

    \I__9948\ : InMux
    port map (
            O => \N__44139\,
            I => \N__44135\
        );

    \I__9947\ : InMux
    port map (
            O => \N__44138\,
            I => \N__44132\
        );

    \I__9946\ : LocalMux
    port map (
            O => \N__44135\,
            I => \N__44128\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__44132\,
            I => \N__44125\
        );

    \I__9944\ : InMux
    port map (
            O => \N__44131\,
            I => \N__44122\
        );

    \I__9943\ : Span4Mux_h
    port map (
            O => \N__44128\,
            I => \N__44119\
        );

    \I__9942\ : Span4Mux_v
    port map (
            O => \N__44125\,
            I => \N__44116\
        );

    \I__9941\ : LocalMux
    port map (
            O => \N__44122\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__44119\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9939\ : Odrv4
    port map (
            O => \N__44116\,
            I => \current_shift_inst.timer_s1.counterZ0Z_25\
        );

    \I__9938\ : InMux
    port map (
            O => \N__44109\,
            I => \current_shift_inst.timer_s1.counter_cry_24\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__44106\,
            I => \N__44103\
        );

    \I__9936\ : InMux
    port map (
            O => \N__44103\,
            I => \N__44099\
        );

    \I__9935\ : InMux
    port map (
            O => \N__44102\,
            I => \N__44096\
        );

    \I__9934\ : LocalMux
    port map (
            O => \N__44099\,
            I => \N__44090\
        );

    \I__9933\ : LocalMux
    port map (
            O => \N__44096\,
            I => \N__44090\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44095\,
            I => \N__44087\
        );

    \I__9931\ : Span4Mux_h
    port map (
            O => \N__44090\,
            I => \N__44084\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__44087\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__9929\ : Odrv4
    port map (
            O => \N__44084\,
            I => \current_shift_inst.timer_s1.counterZ0Z_26\
        );

    \I__9928\ : InMux
    port map (
            O => \N__44079\,
            I => \current_shift_inst.timer_s1.counter_cry_25\
        );

    \I__9927\ : InMux
    port map (
            O => \N__44076\,
            I => \N__44070\
        );

    \I__9926\ : InMux
    port map (
            O => \N__44075\,
            I => \N__44070\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44070\,
            I => \N__44066\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44069\,
            I => \N__44063\
        );

    \I__9923\ : Span4Mux_h
    port map (
            O => \N__44066\,
            I => \N__44060\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__44063\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__9921\ : Odrv4
    port map (
            O => \N__44060\,
            I => \current_shift_inst.timer_s1.counterZ0Z_27\
        );

    \I__9920\ : InMux
    port map (
            O => \N__44055\,
            I => \current_shift_inst.timer_s1.counter_cry_26\
        );

    \I__9919\ : InMux
    port map (
            O => \N__44052\,
            I => \N__44049\
        );

    \I__9918\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__44045\
        );

    \I__9917\ : InMux
    port map (
            O => \N__44048\,
            I => \N__44042\
        );

    \I__9916\ : Span4Mux_h
    port map (
            O => \N__44045\,
            I => \N__44039\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__44042\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__9914\ : Odrv4
    port map (
            O => \N__44039\,
            I => \current_shift_inst.timer_s1.counterZ0Z_28\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44034\,
            I => \N__44028\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44033\,
            I => \N__44028\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__44028\,
            I => \N__44024\
        );

    \I__9910\ : InMux
    port map (
            O => \N__44027\,
            I => \N__44021\
        );

    \I__9909\ : Span4Mux_h
    port map (
            O => \N__44024\,
            I => \N__44018\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__44021\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__9907\ : Odrv4
    port map (
            O => \N__44018\,
            I => \current_shift_inst.timer_s1.counterZ0Z_12\
        );

    \I__9906\ : InMux
    port map (
            O => \N__44013\,
            I => \current_shift_inst.timer_s1.counter_cry_11\
        );

    \I__9905\ : CascadeMux
    port map (
            O => \N__44010\,
            I => \N__44006\
        );

    \I__9904\ : CascadeMux
    port map (
            O => \N__44009\,
            I => \N__44003\
        );

    \I__9903\ : InMux
    port map (
            O => \N__44006\,
            I => \N__43998\
        );

    \I__9902\ : InMux
    port map (
            O => \N__44003\,
            I => \N__43998\
        );

    \I__9901\ : LocalMux
    port map (
            O => \N__43998\,
            I => \N__43994\
        );

    \I__9900\ : InMux
    port map (
            O => \N__43997\,
            I => \N__43991\
        );

    \I__9899\ : Span4Mux_h
    port map (
            O => \N__43994\,
            I => \N__43988\
        );

    \I__9898\ : LocalMux
    port map (
            O => \N__43991\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__43988\,
            I => \current_shift_inst.timer_s1.counterZ0Z_13\
        );

    \I__9896\ : InMux
    port map (
            O => \N__43983\,
            I => \current_shift_inst.timer_s1.counter_cry_12\
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__43980\,
            I => \N__43976\
        );

    \I__9894\ : CascadeMux
    port map (
            O => \N__43979\,
            I => \N__43973\
        );

    \I__9893\ : InMux
    port map (
            O => \N__43976\,
            I => \N__43968\
        );

    \I__9892\ : InMux
    port map (
            O => \N__43973\,
            I => \N__43968\
        );

    \I__9891\ : LocalMux
    port map (
            O => \N__43968\,
            I => \N__43964\
        );

    \I__9890\ : InMux
    port map (
            O => \N__43967\,
            I => \N__43961\
        );

    \I__9889\ : Span4Mux_v
    port map (
            O => \N__43964\,
            I => \N__43958\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__43961\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__43958\,
            I => \current_shift_inst.timer_s1.counterZ0Z_14\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43953\,
            I => \current_shift_inst.timer_s1.counter_cry_13\
        );

    \I__9885\ : CascadeMux
    port map (
            O => \N__43950\,
            I => \N__43947\
        );

    \I__9884\ : InMux
    port map (
            O => \N__43947\,
            I => \N__43943\
        );

    \I__9883\ : InMux
    port map (
            O => \N__43946\,
            I => \N__43940\
        );

    \I__9882\ : LocalMux
    port map (
            O => \N__43943\,
            I => \N__43934\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43940\,
            I => \N__43934\
        );

    \I__9880\ : InMux
    port map (
            O => \N__43939\,
            I => \N__43931\
        );

    \I__9879\ : Span4Mux_v
    port map (
            O => \N__43934\,
            I => \N__43928\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__43931\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9877\ : Odrv4
    port map (
            O => \N__43928\,
            I => \current_shift_inst.timer_s1.counterZ0Z_15\
        );

    \I__9876\ : InMux
    port map (
            O => \N__43923\,
            I => \current_shift_inst.timer_s1.counter_cry_14\
        );

    \I__9875\ : CascadeMux
    port map (
            O => \N__43920\,
            I => \N__43917\
        );

    \I__9874\ : InMux
    port map (
            O => \N__43917\,
            I => \N__43913\
        );

    \I__9873\ : InMux
    port map (
            O => \N__43916\,
            I => \N__43910\
        );

    \I__9872\ : LocalMux
    port map (
            O => \N__43913\,
            I => \N__43904\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__43910\,
            I => \N__43904\
        );

    \I__9870\ : InMux
    port map (
            O => \N__43909\,
            I => \N__43901\
        );

    \I__9869\ : Span4Mux_v
    port map (
            O => \N__43904\,
            I => \N__43898\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__43901\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9867\ : Odrv4
    port map (
            O => \N__43898\,
            I => \current_shift_inst.timer_s1.counterZ0Z_16\
        );

    \I__9866\ : InMux
    port map (
            O => \N__43893\,
            I => \bfn_17_25_0_\
        );

    \I__9865\ : CascadeMux
    port map (
            O => \N__43890\,
            I => \N__43887\
        );

    \I__9864\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43883\
        );

    \I__9863\ : InMux
    port map (
            O => \N__43886\,
            I => \N__43880\
        );

    \I__9862\ : LocalMux
    port map (
            O => \N__43883\,
            I => \N__43876\
        );

    \I__9861\ : LocalMux
    port map (
            O => \N__43880\,
            I => \N__43873\
        );

    \I__9860\ : InMux
    port map (
            O => \N__43879\,
            I => \N__43870\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__43876\,
            I => \N__43867\
        );

    \I__9858\ : Span4Mux_v
    port map (
            O => \N__43873\,
            I => \N__43864\
        );

    \I__9857\ : LocalMux
    port map (
            O => \N__43870\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9856\ : Odrv4
    port map (
            O => \N__43867\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__43864\,
            I => \current_shift_inst.timer_s1.counterZ0Z_17\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43857\,
            I => \current_shift_inst.timer_s1.counter_cry_16\
        );

    \I__9853\ : InMux
    port map (
            O => \N__43854\,
            I => \N__43848\
        );

    \I__9852\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43848\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__43848\,
            I => \N__43844\
        );

    \I__9850\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43841\
        );

    \I__9849\ : Span4Mux_h
    port map (
            O => \N__43844\,
            I => \N__43838\
        );

    \I__9848\ : LocalMux
    port map (
            O => \N__43841\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__43838\,
            I => \current_shift_inst.timer_s1.counterZ0Z_18\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43833\,
            I => \current_shift_inst.timer_s1.counter_cry_17\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43830\,
            I => \N__43824\
        );

    \I__9844\ : InMux
    port map (
            O => \N__43829\,
            I => \N__43824\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__43824\,
            I => \N__43820\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43823\,
            I => \N__43817\
        );

    \I__9841\ : Span4Mux_h
    port map (
            O => \N__43820\,
            I => \N__43814\
        );

    \I__9840\ : LocalMux
    port map (
            O => \N__43817\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9839\ : Odrv4
    port map (
            O => \N__43814\,
            I => \current_shift_inst.timer_s1.counterZ0Z_19\
        );

    \I__9838\ : InMux
    port map (
            O => \N__43809\,
            I => \current_shift_inst.timer_s1.counter_cry_18\
        );

    \I__9837\ : CascadeMux
    port map (
            O => \N__43806\,
            I => \N__43802\
        );

    \I__9836\ : CascadeMux
    port map (
            O => \N__43805\,
            I => \N__43799\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43802\,
            I => \N__43794\
        );

    \I__9834\ : InMux
    port map (
            O => \N__43799\,
            I => \N__43794\
        );

    \I__9833\ : LocalMux
    port map (
            O => \N__43794\,
            I => \N__43790\
        );

    \I__9832\ : InMux
    port map (
            O => \N__43793\,
            I => \N__43787\
        );

    \I__9831\ : Span4Mux_h
    port map (
            O => \N__43790\,
            I => \N__43784\
        );

    \I__9830\ : LocalMux
    port map (
            O => \N__43787\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9829\ : Odrv4
    port map (
            O => \N__43784\,
            I => \current_shift_inst.timer_s1.counterZ0Z_3\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43779\,
            I => \current_shift_inst.timer_s1.counter_cry_2\
        );

    \I__9827\ : CascadeMux
    port map (
            O => \N__43776\,
            I => \N__43772\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__43775\,
            I => \N__43769\
        );

    \I__9825\ : InMux
    port map (
            O => \N__43772\,
            I => \N__43764\
        );

    \I__9824\ : InMux
    port map (
            O => \N__43769\,
            I => \N__43764\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43764\,
            I => \N__43760\
        );

    \I__9822\ : InMux
    port map (
            O => \N__43763\,
            I => \N__43757\
        );

    \I__9821\ : Span4Mux_v
    port map (
            O => \N__43760\,
            I => \N__43754\
        );

    \I__9820\ : LocalMux
    port map (
            O => \N__43757\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9819\ : Odrv4
    port map (
            O => \N__43754\,
            I => \current_shift_inst.timer_s1.counterZ0Z_4\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43749\,
            I => \current_shift_inst.timer_s1.counter_cry_3\
        );

    \I__9817\ : CascadeMux
    port map (
            O => \N__43746\,
            I => \N__43743\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43739\
        );

    \I__9815\ : InMux
    port map (
            O => \N__43742\,
            I => \N__43736\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__43739\,
            I => \N__43730\
        );

    \I__9813\ : LocalMux
    port map (
            O => \N__43736\,
            I => \N__43730\
        );

    \I__9812\ : InMux
    port map (
            O => \N__43735\,
            I => \N__43727\
        );

    \I__9811\ : Span4Mux_h
    port map (
            O => \N__43730\,
            I => \N__43724\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43727\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9809\ : Odrv4
    port map (
            O => \N__43724\,
            I => \current_shift_inst.timer_s1.counterZ0Z_5\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43719\,
            I => \current_shift_inst.timer_s1.counter_cry_4\
        );

    \I__9807\ : InMux
    port map (
            O => \N__43716\,
            I => \N__43710\
        );

    \I__9806\ : InMux
    port map (
            O => \N__43715\,
            I => \N__43710\
        );

    \I__9805\ : LocalMux
    port map (
            O => \N__43710\,
            I => \N__43706\
        );

    \I__9804\ : InMux
    port map (
            O => \N__43709\,
            I => \N__43703\
        );

    \I__9803\ : Span4Mux_v
    port map (
            O => \N__43706\,
            I => \N__43700\
        );

    \I__9802\ : LocalMux
    port map (
            O => \N__43703\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__43700\,
            I => \current_shift_inst.timer_s1.counterZ0Z_6\
        );

    \I__9800\ : InMux
    port map (
            O => \N__43695\,
            I => \current_shift_inst.timer_s1.counter_cry_5\
        );

    \I__9799\ : InMux
    port map (
            O => \N__43692\,
            I => \N__43686\
        );

    \I__9798\ : InMux
    port map (
            O => \N__43691\,
            I => \N__43686\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__43686\,
            I => \N__43682\
        );

    \I__9796\ : InMux
    port map (
            O => \N__43685\,
            I => \N__43679\
        );

    \I__9795\ : Span4Mux_v
    port map (
            O => \N__43682\,
            I => \N__43676\
        );

    \I__9794\ : LocalMux
    port map (
            O => \N__43679\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9793\ : Odrv4
    port map (
            O => \N__43676\,
            I => \current_shift_inst.timer_s1.counterZ0Z_7\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43671\,
            I => \current_shift_inst.timer_s1.counter_cry_6\
        );

    \I__9791\ : CascadeMux
    port map (
            O => \N__43668\,
            I => \N__43664\
        );

    \I__9790\ : CascadeMux
    port map (
            O => \N__43667\,
            I => \N__43661\
        );

    \I__9789\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43658\
        );

    \I__9788\ : InMux
    port map (
            O => \N__43661\,
            I => \N__43655\
        );

    \I__9787\ : LocalMux
    port map (
            O => \N__43658\,
            I => \N__43649\
        );

    \I__9786\ : LocalMux
    port map (
            O => \N__43655\,
            I => \N__43649\
        );

    \I__9785\ : InMux
    port map (
            O => \N__43654\,
            I => \N__43646\
        );

    \I__9784\ : Span4Mux_v
    port map (
            O => \N__43649\,
            I => \N__43643\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__43646\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9782\ : Odrv4
    port map (
            O => \N__43643\,
            I => \current_shift_inst.timer_s1.counterZ0Z_8\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43638\,
            I => \bfn_17_24_0_\
        );

    \I__9780\ : CascadeMux
    port map (
            O => \N__43635\,
            I => \N__43631\
        );

    \I__9779\ : CascadeMux
    port map (
            O => \N__43634\,
            I => \N__43628\
        );

    \I__9778\ : InMux
    port map (
            O => \N__43631\,
            I => \N__43625\
        );

    \I__9777\ : InMux
    port map (
            O => \N__43628\,
            I => \N__43622\
        );

    \I__9776\ : LocalMux
    port map (
            O => \N__43625\,
            I => \N__43619\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__43622\,
            I => \N__43615\
        );

    \I__9774\ : Span4Mux_v
    port map (
            O => \N__43619\,
            I => \N__43612\
        );

    \I__9773\ : InMux
    port map (
            O => \N__43618\,
            I => \N__43609\
        );

    \I__9772\ : Span4Mux_h
    port map (
            O => \N__43615\,
            I => \N__43604\
        );

    \I__9771\ : Span4Mux_h
    port map (
            O => \N__43612\,
            I => \N__43604\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__43609\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9769\ : Odrv4
    port map (
            O => \N__43604\,
            I => \current_shift_inst.timer_s1.counterZ0Z_9\
        );

    \I__9768\ : InMux
    port map (
            O => \N__43599\,
            I => \current_shift_inst.timer_s1.counter_cry_8\
        );

    \I__9767\ : CascadeMux
    port map (
            O => \N__43596\,
            I => \N__43593\
        );

    \I__9766\ : InMux
    port map (
            O => \N__43593\,
            I => \N__43589\
        );

    \I__9765\ : InMux
    port map (
            O => \N__43592\,
            I => \N__43586\
        );

    \I__9764\ : LocalMux
    port map (
            O => \N__43589\,
            I => \N__43580\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__43586\,
            I => \N__43580\
        );

    \I__9762\ : InMux
    port map (
            O => \N__43585\,
            I => \N__43577\
        );

    \I__9761\ : Span4Mux_h
    port map (
            O => \N__43580\,
            I => \N__43574\
        );

    \I__9760\ : LocalMux
    port map (
            O => \N__43577\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__9759\ : Odrv4
    port map (
            O => \N__43574\,
            I => \current_shift_inst.timer_s1.counterZ0Z_10\
        );

    \I__9758\ : InMux
    port map (
            O => \N__43569\,
            I => \current_shift_inst.timer_s1.counter_cry_9\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43566\,
            I => \N__43560\
        );

    \I__9756\ : InMux
    port map (
            O => \N__43565\,
            I => \N__43560\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__43560\,
            I => \N__43556\
        );

    \I__9754\ : InMux
    port map (
            O => \N__43559\,
            I => \N__43553\
        );

    \I__9753\ : Span4Mux_h
    port map (
            O => \N__43556\,
            I => \N__43550\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43553\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__9751\ : Odrv4
    port map (
            O => \N__43550\,
            I => \current_shift_inst.timer_s1.counterZ0Z_11\
        );

    \I__9750\ : InMux
    port map (
            O => \N__43545\,
            I => \current_shift_inst.timer_s1.counter_cry_10\
        );

    \I__9749\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43539\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__43539\,
            I => \N__43536\
        );

    \I__9747\ : Odrv12
    port map (
            O => \N__43536\,
            I => \current_shift_inst.un4_control_input_1_axb_20\
        );

    \I__9746\ : CascadeMux
    port map (
            O => \N__43533\,
            I => \N__43529\
        );

    \I__9745\ : CascadeMux
    port map (
            O => \N__43532\,
            I => \N__43526\
        );

    \I__9744\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43523\
        );

    \I__9743\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43520\
        );

    \I__9742\ : LocalMux
    port map (
            O => \N__43523\,
            I => \N__43514\
        );

    \I__9741\ : LocalMux
    port map (
            O => \N__43520\,
            I => \N__43514\
        );

    \I__9740\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43511\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__43514\,
            I => \N__43507\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__43511\,
            I => \N__43504\
        );

    \I__9737\ : InMux
    port map (
            O => \N__43510\,
            I => \N__43501\
        );

    \I__9736\ : Odrv4
    port map (
            O => \N__43507\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9735\ : Odrv4
    port map (
            O => \N__43504\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9734\ : LocalMux
    port map (
            O => \N__43501\,
            I => \current_shift_inst.elapsed_time_ns_s1_30\
        );

    \I__9733\ : InMux
    port map (
            O => \N__43494\,
            I => \N__43491\
        );

    \I__9732\ : LocalMux
    port map (
            O => \N__43491\,
            I => \N__43488\
        );

    \I__9731\ : Odrv12
    port map (
            O => \N__43488\,
            I => \current_shift_inst.un4_control_input_1_axb_29\
        );

    \I__9730\ : InMux
    port map (
            O => \N__43485\,
            I => \N__43481\
        );

    \I__9729\ : InMux
    port map (
            O => \N__43484\,
            I => \N__43477\
        );

    \I__9728\ : LocalMux
    port map (
            O => \N__43481\,
            I => \N__43474\
        );

    \I__9727\ : InMux
    port map (
            O => \N__43480\,
            I => \N__43471\
        );

    \I__9726\ : LocalMux
    port map (
            O => \N__43477\,
            I => \N__43465\
        );

    \I__9725\ : Span4Mux_v
    port map (
            O => \N__43474\,
            I => \N__43465\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__43471\,
            I => \N__43462\
        );

    \I__9723\ : InMux
    port map (
            O => \N__43470\,
            I => \N__43459\
        );

    \I__9722\ : Odrv4
    port map (
            O => \N__43465\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9721\ : Odrv4
    port map (
            O => \N__43462\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9720\ : LocalMux
    port map (
            O => \N__43459\,
            I => \current_shift_inst.elapsed_time_ns_s1_15\
        );

    \I__9719\ : CascadeMux
    port map (
            O => \N__43452\,
            I => \N__43449\
        );

    \I__9718\ : InMux
    port map (
            O => \N__43449\,
            I => \N__43445\
        );

    \I__9717\ : CascadeMux
    port map (
            O => \N__43448\,
            I => \N__43442\
        );

    \I__9716\ : LocalMux
    port map (
            O => \N__43445\,
            I => \N__43438\
        );

    \I__9715\ : InMux
    port map (
            O => \N__43442\,
            I => \N__43435\
        );

    \I__9714\ : InMux
    port map (
            O => \N__43441\,
            I => \N__43432\
        );

    \I__9713\ : Span4Mux_v
    port map (
            O => \N__43438\,
            I => \N__43429\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__43435\,
            I => \N__43426\
        );

    \I__9711\ : LocalMux
    port map (
            O => \N__43432\,
            I => \N__43423\
        );

    \I__9710\ : Span4Mux_h
    port map (
            O => \N__43429\,
            I => \N__43420\
        );

    \I__9709\ : Span4Mux_h
    port map (
            O => \N__43426\,
            I => \N__43417\
        );

    \I__9708\ : Span4Mux_v
    port map (
            O => \N__43423\,
            I => \N__43414\
        );

    \I__9707\ : Odrv4
    port map (
            O => \N__43420\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9706\ : Odrv4
    port map (
            O => \N__43417\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9705\ : Odrv4
    port map (
            O => \N__43414\,
            I => \current_shift_inst.un4_control_input1_15\
        );

    \I__9704\ : CascadeMux
    port map (
            O => \N__43407\,
            I => \N__43404\
        );

    \I__9703\ : InMux
    port map (
            O => \N__43404\,
            I => \N__43401\
        );

    \I__9702\ : LocalMux
    port map (
            O => \N__43401\,
            I => \N__43398\
        );

    \I__9701\ : Span4Mux_h
    port map (
            O => \N__43398\,
            I => \N__43395\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__43395\,
            I => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\
        );

    \I__9699\ : InMux
    port map (
            O => \N__43392\,
            I => \N__43389\
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__43389\,
            I => \N__43386\
        );

    \I__9697\ : Odrv4
    port map (
            O => \N__43386\,
            I => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\
        );

    \I__9696\ : CascadeMux
    port map (
            O => \N__43383\,
            I => \N__43379\
        );

    \I__9695\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43376\
        );

    \I__9694\ : InMux
    port map (
            O => \N__43379\,
            I => \N__43372\
        );

    \I__9693\ : LocalMux
    port map (
            O => \N__43376\,
            I => \N__43368\
        );

    \I__9692\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43365\
        );

    \I__9691\ : LocalMux
    port map (
            O => \N__43372\,
            I => \N__43362\
        );

    \I__9690\ : InMux
    port map (
            O => \N__43371\,
            I => \N__43359\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__43368\,
            I => \N__43354\
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__43365\,
            I => \N__43354\
        );

    \I__9687\ : Span4Mux_v
    port map (
            O => \N__43362\,
            I => \N__43349\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__43359\,
            I => \N__43349\
        );

    \I__9685\ : Odrv4
    port map (
            O => \N__43354\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__9684\ : Odrv4
    port map (
            O => \N__43349\,
            I => \current_shift_inst.elapsed_time_ns_s1_12\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43344\,
            I => \N__43340\
        );

    \I__9682\ : InMux
    port map (
            O => \N__43343\,
            I => \N__43337\
        );

    \I__9681\ : LocalMux
    port map (
            O => \N__43340\,
            I => \N__43333\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__43337\,
            I => \N__43330\
        );

    \I__9679\ : InMux
    port map (
            O => \N__43336\,
            I => \N__43327\
        );

    \I__9678\ : Span12Mux_h
    port map (
            O => \N__43333\,
            I => \N__43324\
        );

    \I__9677\ : Span12Mux_h
    port map (
            O => \N__43330\,
            I => \N__43319\
        );

    \I__9676\ : LocalMux
    port map (
            O => \N__43327\,
            I => \N__43319\
        );

    \I__9675\ : Odrv12
    port map (
            O => \N__43324\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9674\ : Odrv12
    port map (
            O => \N__43319\,
            I => \current_shift_inst.un4_control_input1_12\
        );

    \I__9673\ : InMux
    port map (
            O => \N__43314\,
            I => \N__43311\
        );

    \I__9672\ : LocalMux
    port map (
            O => \N__43311\,
            I => \N__43308\
        );

    \I__9671\ : Odrv12
    port map (
            O => \N__43308\,
            I => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\
        );

    \I__9670\ : InMux
    port map (
            O => \N__43305\,
            I => \bfn_17_23_0_\
        );

    \I__9669\ : InMux
    port map (
            O => \N__43302\,
            I => \current_shift_inst.timer_s1.counter_cry_0\
        );

    \I__9668\ : CascadeMux
    port map (
            O => \N__43299\,
            I => \N__43295\
        );

    \I__9667\ : InMux
    port map (
            O => \N__43298\,
            I => \N__43292\
        );

    \I__9666\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43289\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43292\,
            I => \N__43283\
        );

    \I__9664\ : LocalMux
    port map (
            O => \N__43289\,
            I => \N__43283\
        );

    \I__9663\ : InMux
    port map (
            O => \N__43288\,
            I => \N__43280\
        );

    \I__9662\ : Sp12to4
    port map (
            O => \N__43283\,
            I => \N__43277\
        );

    \I__9661\ : LocalMux
    port map (
            O => \N__43280\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9660\ : Odrv12
    port map (
            O => \N__43277\,
            I => \current_shift_inst.timer_s1.counterZ0Z_2\
        );

    \I__9659\ : InMux
    port map (
            O => \N__43272\,
            I => \current_shift_inst.timer_s1.counter_cry_1\
        );

    \I__9658\ : InMux
    port map (
            O => \N__43269\,
            I => \N__43266\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__43266\,
            I => \N__43263\
        );

    \I__9656\ : Odrv12
    port map (
            O => \N__43263\,
            I => \current_shift_inst.un4_control_input_1_axb_14\
        );

    \I__9655\ : CascadeMux
    port map (
            O => \N__43260\,
            I => \N__43257\
        );

    \I__9654\ : InMux
    port map (
            O => \N__43257\,
            I => \N__43253\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43256\,
            I => \N__43250\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43253\,
            I => \N__43246\
        );

    \I__9651\ : LocalMux
    port map (
            O => \N__43250\,
            I => \N__43243\
        );

    \I__9650\ : InMux
    port map (
            O => \N__43249\,
            I => \N__43240\
        );

    \I__9649\ : Span4Mux_h
    port map (
            O => \N__43246\,
            I => \N__43236\
        );

    \I__9648\ : Span4Mux_v
    port map (
            O => \N__43243\,
            I => \N__43233\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__43240\,
            I => \N__43230\
        );

    \I__9646\ : InMux
    port map (
            O => \N__43239\,
            I => \N__43227\
        );

    \I__9645\ : Odrv4
    port map (
            O => \N__43236\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9644\ : Odrv4
    port map (
            O => \N__43233\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9643\ : Odrv12
    port map (
            O => \N__43230\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9642\ : LocalMux
    port map (
            O => \N__43227\,
            I => \current_shift_inst.elapsed_time_ns_s1_17\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43215\
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__43215\,
            I => \N__43212\
        );

    \I__9639\ : Odrv12
    port map (
            O => \N__43212\,
            I => \current_shift_inst.un4_control_input_1_axb_16\
        );

    \I__9638\ : CascadeMux
    port map (
            O => \N__43209\,
            I => \N__43206\
        );

    \I__9637\ : InMux
    port map (
            O => \N__43206\,
            I => \N__43202\
        );

    \I__9636\ : InMux
    port map (
            O => \N__43205\,
            I => \N__43198\
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__43202\,
            I => \N__43195\
        );

    \I__9634\ : InMux
    port map (
            O => \N__43201\,
            I => \N__43192\
        );

    \I__9633\ : LocalMux
    port map (
            O => \N__43198\,
            I => \N__43188\
        );

    \I__9632\ : Span4Mux_v
    port map (
            O => \N__43195\,
            I => \N__43183\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__43192\,
            I => \N__43183\
        );

    \I__9630\ : InMux
    port map (
            O => \N__43191\,
            I => \N__43180\
        );

    \I__9629\ : Odrv4
    port map (
            O => \N__43188\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9628\ : Odrv4
    port map (
            O => \N__43183\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43180\,
            I => \current_shift_inst.elapsed_time_ns_s1_26\
        );

    \I__9626\ : InMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__9625\ : LocalMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__9624\ : Odrv4
    port map (
            O => \N__43167\,
            I => \current_shift_inst.un4_control_input_1_axb_25\
        );

    \I__9623\ : InMux
    port map (
            O => \N__43164\,
            I => \N__43160\
        );

    \I__9622\ : CascadeMux
    port map (
            O => \N__43163\,
            I => \N__43157\
        );

    \I__9621\ : LocalMux
    port map (
            O => \N__43160\,
            I => \N__43154\
        );

    \I__9620\ : InMux
    port map (
            O => \N__43157\,
            I => \N__43151\
        );

    \I__9619\ : Span4Mux_h
    port map (
            O => \N__43154\,
            I => \N__43147\
        );

    \I__9618\ : LocalMux
    port map (
            O => \N__43151\,
            I => \N__43144\
        );

    \I__9617\ : InMux
    port map (
            O => \N__43150\,
            I => \N__43141\
        );

    \I__9616\ : Span4Mux_h
    port map (
            O => \N__43147\,
            I => \N__43135\
        );

    \I__9615\ : Span4Mux_v
    port map (
            O => \N__43144\,
            I => \N__43135\
        );

    \I__9614\ : LocalMux
    port map (
            O => \N__43141\,
            I => \N__43132\
        );

    \I__9613\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43129\
        );

    \I__9612\ : Odrv4
    port map (
            O => \N__43135\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9611\ : Odrv4
    port map (
            O => \N__43132\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9610\ : LocalMux
    port map (
            O => \N__43129\,
            I => \current_shift_inst.elapsed_time_ns_s1_19\
        );

    \I__9609\ : CascadeMux
    port map (
            O => \N__43122\,
            I => \N__43119\
        );

    \I__9608\ : InMux
    port map (
            O => \N__43119\,
            I => \N__43116\
        );

    \I__9607\ : LocalMux
    port map (
            O => \N__43116\,
            I => \N__43113\
        );

    \I__9606\ : Odrv4
    port map (
            O => \N__43113\,
            I => \current_shift_inst.un4_control_input_1_axb_18\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__43110\,
            I => \N__43107\
        );

    \I__9604\ : InMux
    port map (
            O => \N__43107\,
            I => \N__43104\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__43104\,
            I => \N__43099\
        );

    \I__9602\ : InMux
    port map (
            O => \N__43103\,
            I => \N__43096\
        );

    \I__9601\ : InMux
    port map (
            O => \N__43102\,
            I => \N__43093\
        );

    \I__9600\ : Span12Mux_v
    port map (
            O => \N__43099\,
            I => \N__43089\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__43096\,
            I => \N__43084\
        );

    \I__9598\ : LocalMux
    port map (
            O => \N__43093\,
            I => \N__43084\
        );

    \I__9597\ : InMux
    port map (
            O => \N__43092\,
            I => \N__43081\
        );

    \I__9596\ : Odrv12
    port map (
            O => \N__43089\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9595\ : Odrv12
    port map (
            O => \N__43084\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__43081\,
            I => \current_shift_inst.elapsed_time_ns_s1_16\
        );

    \I__9593\ : InMux
    port map (
            O => \N__43074\,
            I => \N__43071\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__43071\,
            I => \N__43068\
        );

    \I__9591\ : Span4Mux_v
    port map (
            O => \N__43068\,
            I => \N__43065\
        );

    \I__9590\ : Odrv4
    port map (
            O => \N__43065\,
            I => \current_shift_inst.un4_control_input_1_axb_15\
        );

    \I__9589\ : CascadeMux
    port map (
            O => \N__43062\,
            I => \N__43058\
        );

    \I__9588\ : CascadeMux
    port map (
            O => \N__43061\,
            I => \N__43055\
        );

    \I__9587\ : InMux
    port map (
            O => \N__43058\,
            I => \N__43052\
        );

    \I__9586\ : InMux
    port map (
            O => \N__43055\,
            I => \N__43049\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43052\,
            I => \N__43043\
        );

    \I__9584\ : LocalMux
    port map (
            O => \N__43049\,
            I => \N__43043\
        );

    \I__9583\ : InMux
    port map (
            O => \N__43048\,
            I => \N__43040\
        );

    \I__9582\ : Span12Mux_v
    port map (
            O => \N__43043\,
            I => \N__43036\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43040\,
            I => \N__43033\
        );

    \I__9580\ : InMux
    port map (
            O => \N__43039\,
            I => \N__43030\
        );

    \I__9579\ : Odrv12
    port map (
            O => \N__43036\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9578\ : Odrv12
    port map (
            O => \N__43033\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9577\ : LocalMux
    port map (
            O => \N__43030\,
            I => \current_shift_inst.elapsed_time_ns_s1_25\
        );

    \I__9576\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__43020\,
            I => \N__43017\
        );

    \I__9574\ : Odrv12
    port map (
            O => \N__43017\,
            I => \current_shift_inst.un4_control_input_1_axb_24\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__43014\,
            I => \N__43010\
        );

    \I__9572\ : CascadeMux
    port map (
            O => \N__43013\,
            I => \N__43007\
        );

    \I__9571\ : InMux
    port map (
            O => \N__43010\,
            I => \N__43004\
        );

    \I__9570\ : InMux
    port map (
            O => \N__43007\,
            I => \N__43001\
        );

    \I__9569\ : LocalMux
    port map (
            O => \N__43004\,
            I => \N__42998\
        );

    \I__9568\ : LocalMux
    port map (
            O => \N__43001\,
            I => \N__42994\
        );

    \I__9567\ : Span4Mux_h
    port map (
            O => \N__42998\,
            I => \N__42991\
        );

    \I__9566\ : InMux
    port map (
            O => \N__42997\,
            I => \N__42988\
        );

    \I__9565\ : Span4Mux_h
    port map (
            O => \N__42994\,
            I => \N__42984\
        );

    \I__9564\ : Span4Mux_v
    port map (
            O => \N__42991\,
            I => \N__42979\
        );

    \I__9563\ : LocalMux
    port map (
            O => \N__42988\,
            I => \N__42979\
        );

    \I__9562\ : InMux
    port map (
            O => \N__42987\,
            I => \N__42976\
        );

    \I__9561\ : Odrv4
    port map (
            O => \N__42984\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9560\ : Odrv4
    port map (
            O => \N__42979\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9559\ : LocalMux
    port map (
            O => \N__42976\,
            I => \current_shift_inst.elapsed_time_ns_s1_29\
        );

    \I__9558\ : InMux
    port map (
            O => \N__42969\,
            I => \N__42966\
        );

    \I__9557\ : LocalMux
    port map (
            O => \N__42966\,
            I => \N__42963\
        );

    \I__9556\ : Odrv4
    port map (
            O => \N__42963\,
            I => \current_shift_inst.un4_control_input_1_axb_28\
        );

    \I__9555\ : CascadeMux
    port map (
            O => \N__42960\,
            I => \N__42956\
        );

    \I__9554\ : CascadeMux
    port map (
            O => \N__42959\,
            I => \N__42953\
        );

    \I__9553\ : InMux
    port map (
            O => \N__42956\,
            I => \N__42950\
        );

    \I__9552\ : InMux
    port map (
            O => \N__42953\,
            I => \N__42947\
        );

    \I__9551\ : LocalMux
    port map (
            O => \N__42950\,
            I => \N__42944\
        );

    \I__9550\ : LocalMux
    port map (
            O => \N__42947\,
            I => \N__42941\
        );

    \I__9549\ : Sp12to4
    port map (
            O => \N__42944\,
            I => \N__42934\
        );

    \I__9548\ : Span12Mux_h
    port map (
            O => \N__42941\,
            I => \N__42934\
        );

    \I__9547\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42931\
        );

    \I__9546\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42928\
        );

    \I__9545\ : Odrv12
    port map (
            O => \N__42934\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9544\ : LocalMux
    port map (
            O => \N__42931\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9543\ : LocalMux
    port map (
            O => \N__42928\,
            I => \current_shift_inst.elapsed_time_ns_s1_27\
        );

    \I__9542\ : InMux
    port map (
            O => \N__42921\,
            I => \N__42918\
        );

    \I__9541\ : LocalMux
    port map (
            O => \N__42918\,
            I => \N__42915\
        );

    \I__9540\ : Odrv4
    port map (
            O => \N__42915\,
            I => \current_shift_inst.un4_control_input_1_axb_26\
        );

    \I__9539\ : CascadeMux
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__9538\ : InMux
    port map (
            O => \N__42909\,
            I => \N__42905\
        );

    \I__9537\ : InMux
    port map (
            O => \N__42908\,
            I => \N__42902\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__42905\,
            I => \N__42897\
        );

    \I__9535\ : LocalMux
    port map (
            O => \N__42902\,
            I => \N__42897\
        );

    \I__9534\ : Span4Mux_h
    port map (
            O => \N__42897\,
            I => \N__42892\
        );

    \I__9533\ : InMux
    port map (
            O => \N__42896\,
            I => \N__42889\
        );

    \I__9532\ : InMux
    port map (
            O => \N__42895\,
            I => \N__42886\
        );

    \I__9531\ : Odrv4
    port map (
            O => \N__42892\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9530\ : LocalMux
    port map (
            O => \N__42889\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9529\ : LocalMux
    port map (
            O => \N__42886\,
            I => \current_shift_inst.elapsed_time_ns_s1_28\
        );

    \I__9528\ : InMux
    port map (
            O => \N__42879\,
            I => \N__42876\
        );

    \I__9527\ : LocalMux
    port map (
            O => \N__42876\,
            I => \N__42873\
        );

    \I__9526\ : Odrv4
    port map (
            O => \N__42873\,
            I => \current_shift_inst.un4_control_input_1_axb_27\
        );

    \I__9525\ : CascadeMux
    port map (
            O => \N__42870\,
            I => \N__42867\
        );

    \I__9524\ : InMux
    port map (
            O => \N__42867\,
            I => \N__42863\
        );

    \I__9523\ : InMux
    port map (
            O => \N__42866\,
            I => \N__42860\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__42863\,
            I => \N__42856\
        );

    \I__9521\ : LocalMux
    port map (
            O => \N__42860\,
            I => \N__42853\
        );

    \I__9520\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42850\
        );

    \I__9519\ : Span4Mux_v
    port map (
            O => \N__42856\,
            I => \N__42845\
        );

    \I__9518\ : Span4Mux_h
    port map (
            O => \N__42853\,
            I => \N__42845\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__42850\,
            I => \N__42841\
        );

    \I__9516\ : Span4Mux_v
    port map (
            O => \N__42845\,
            I => \N__42838\
        );

    \I__9515\ : InMux
    port map (
            O => \N__42844\,
            I => \N__42835\
        );

    \I__9514\ : Odrv12
    port map (
            O => \N__42841\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9513\ : Odrv4
    port map (
            O => \N__42838\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42835\,
            I => \current_shift_inst.elapsed_time_ns_s1_4\
        );

    \I__9511\ : InMux
    port map (
            O => \N__42828\,
            I => \N__42825\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__42825\,
            I => \N__42822\
        );

    \I__9509\ : Odrv12
    port map (
            O => \N__42822\,
            I => \current_shift_inst.un4_control_input_1_axb_3\
        );

    \I__9508\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42814\
        );

    \I__9507\ : CascadeMux
    port map (
            O => \N__42818\,
            I => \N__42811\
        );

    \I__9506\ : CascadeMux
    port map (
            O => \N__42817\,
            I => \N__42808\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__42814\,
            I => \N__42805\
        );

    \I__9504\ : InMux
    port map (
            O => \N__42811\,
            I => \N__42800\
        );

    \I__9503\ : InMux
    port map (
            O => \N__42808\,
            I => \N__42800\
        );

    \I__9502\ : Span4Mux_h
    port map (
            O => \N__42805\,
            I => \N__42794\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__42800\,
            I => \N__42794\
        );

    \I__9500\ : InMux
    port map (
            O => \N__42799\,
            I => \N__42791\
        );

    \I__9499\ : Odrv4
    port map (
            O => \N__42794\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42791\,
            I => \current_shift_inst.elapsed_time_ns_s1_6\
        );

    \I__9497\ : InMux
    port map (
            O => \N__42786\,
            I => \N__42783\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__42783\,
            I => \N__42780\
        );

    \I__9495\ : Odrv12
    port map (
            O => \N__42780\,
            I => \current_shift_inst.un4_control_input_1_axb_5\
        );

    \I__9494\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42774\
        );

    \I__9493\ : LocalMux
    port map (
            O => \N__42774\,
            I => \N__42771\
        );

    \I__9492\ : Odrv4
    port map (
            O => \N__42771\,
            I => \current_shift_inst.un4_control_input_1_axb_13\
        );

    \I__9491\ : InMux
    port map (
            O => \N__42768\,
            I => \N__42765\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__42765\,
            I => \N__42762\
        );

    \I__9489\ : Odrv4
    port map (
            O => \N__42762\,
            I => \current_shift_inst.un4_control_input_1_axb_12\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42759\,
            I => \N__42754\
        );

    \I__9487\ : InMux
    port map (
            O => \N__42758\,
            I => \N__42751\
        );

    \I__9486\ : CascadeMux
    port map (
            O => \N__42757\,
            I => \N__42748\
        );

    \I__9485\ : LocalMux
    port map (
            O => \N__42754\,
            I => \N__42745\
        );

    \I__9484\ : LocalMux
    port map (
            O => \N__42751\,
            I => \N__42742\
        );

    \I__9483\ : InMux
    port map (
            O => \N__42748\,
            I => \N__42739\
        );

    \I__9482\ : Sp12to4
    port map (
            O => \N__42745\,
            I => \N__42731\
        );

    \I__9481\ : Sp12to4
    port map (
            O => \N__42742\,
            I => \N__42731\
        );

    \I__9480\ : LocalMux
    port map (
            O => \N__42739\,
            I => \N__42731\
        );

    \I__9479\ : InMux
    port map (
            O => \N__42738\,
            I => \N__42728\
        );

    \I__9478\ : Odrv12
    port map (
            O => \N__42731\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42728\,
            I => \current_shift_inst.elapsed_time_ns_s1_7\
        );

    \I__9476\ : InMux
    port map (
            O => \N__42723\,
            I => \N__42720\
        );

    \I__9475\ : LocalMux
    port map (
            O => \N__42720\,
            I => \N__42717\
        );

    \I__9474\ : Odrv12
    port map (
            O => \N__42717\,
            I => \current_shift_inst.un4_control_input_1_axb_6\
        );

    \I__9473\ : CascadeMux
    port map (
            O => \N__42714\,
            I => \N__42710\
        );

    \I__9472\ : CascadeMux
    port map (
            O => \N__42713\,
            I => \N__42707\
        );

    \I__9471\ : InMux
    port map (
            O => \N__42710\,
            I => \N__42704\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42707\,
            I => \N__42701\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__42704\,
            I => \N__42698\
        );

    \I__9468\ : LocalMux
    port map (
            O => \N__42701\,
            I => \N__42694\
        );

    \I__9467\ : Span4Mux_h
    port map (
            O => \N__42698\,
            I => \N__42691\
        );

    \I__9466\ : InMux
    port map (
            O => \N__42697\,
            I => \N__42688\
        );

    \I__9465\ : Span4Mux_v
    port map (
            O => \N__42694\,
            I => \N__42684\
        );

    \I__9464\ : Sp12to4
    port map (
            O => \N__42691\,
            I => \N__42679\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__42688\,
            I => \N__42679\
        );

    \I__9462\ : InMux
    port map (
            O => \N__42687\,
            I => \N__42676\
        );

    \I__9461\ : Odrv4
    port map (
            O => \N__42684\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9460\ : Odrv12
    port map (
            O => \N__42679\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9459\ : LocalMux
    port map (
            O => \N__42676\,
            I => \current_shift_inst.elapsed_time_ns_s1_9\
        );

    \I__9458\ : InMux
    port map (
            O => \N__42669\,
            I => \N__42666\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42666\,
            I => \N__42663\
        );

    \I__9456\ : Span4Mux_v
    port map (
            O => \N__42663\,
            I => \N__42660\
        );

    \I__9455\ : Odrv4
    port map (
            O => \N__42660\,
            I => \current_shift_inst.un4_control_input_1_axb_8\
        );

    \I__9454\ : InMux
    port map (
            O => \N__42657\,
            I => \N__42653\
        );

    \I__9453\ : InMux
    port map (
            O => \N__42656\,
            I => \N__42650\
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42653\,
            I => \N__42647\
        );

    \I__9451\ : LocalMux
    port map (
            O => \N__42650\,
            I => \N__42644\
        );

    \I__9450\ : Span4Mux_v
    port map (
            O => \N__42647\,
            I => \N__42641\
        );

    \I__9449\ : Span4Mux_v
    port map (
            O => \N__42644\,
            I => \N__42637\
        );

    \I__9448\ : Span4Mux_h
    port map (
            O => \N__42641\,
            I => \N__42634\
        );

    \I__9447\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42631\
        );

    \I__9446\ : Span4Mux_v
    port map (
            O => \N__42637\,
            I => \N__42628\
        );

    \I__9445\ : Odrv4
    port map (
            O => \N__42634\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__42631\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9443\ : Odrv4
    port map (
            O => \N__42628\,
            I => \current_shift_inst.un4_control_input1_26\
        );

    \I__9442\ : InMux
    port map (
            O => \N__42621\,
            I => \N__42618\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__42618\,
            I => \N__42615\
        );

    \I__9440\ : Odrv12
    port map (
            O => \N__42615\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\
        );

    \I__9439\ : CascadeMux
    port map (
            O => \N__42612\,
            I => \N__42609\
        );

    \I__9438\ : InMux
    port map (
            O => \N__42609\,
            I => \N__42606\
        );

    \I__9437\ : LocalMux
    port map (
            O => \N__42606\,
            I => \N__42602\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42605\,
            I => \N__42599\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__42602\,
            I => \N__42593\
        );

    \I__9434\ : LocalMux
    port map (
            O => \N__42599\,
            I => \N__42593\
        );

    \I__9433\ : InMux
    port map (
            O => \N__42598\,
            I => \N__42590\
        );

    \I__9432\ : Sp12to4
    port map (
            O => \N__42593\,
            I => \N__42586\
        );

    \I__9431\ : LocalMux
    port map (
            O => \N__42590\,
            I => \N__42583\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42589\,
            I => \N__42580\
        );

    \I__9429\ : Odrv12
    port map (
            O => \N__42586\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9428\ : Odrv4
    port map (
            O => \N__42583\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9427\ : LocalMux
    port map (
            O => \N__42580\,
            I => \current_shift_inst.elapsed_time_ns_s1_20\
        );

    \I__9426\ : InMux
    port map (
            O => \N__42573\,
            I => \N__42570\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__42570\,
            I => \N__42567\
        );

    \I__9424\ : Odrv4
    port map (
            O => \N__42567\,
            I => \current_shift_inst.un4_control_input_1_axb_19\
        );

    \I__9423\ : InMux
    port map (
            O => \N__42564\,
            I => \N__42561\
        );

    \I__9422\ : LocalMux
    port map (
            O => \N__42561\,
            I => \current_shift_inst.un4_control_input_1_axb_22\
        );

    \I__9421\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42555\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__42555\,
            I => \N__42552\
        );

    \I__9419\ : Span4Mux_h
    port map (
            O => \N__42552\,
            I => \N__42547\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42551\,
            I => \N__42544\
        );

    \I__9417\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42541\
        );

    \I__9416\ : Odrv4
    port map (
            O => \N__42547\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9415\ : LocalMux
    port map (
            O => \N__42544\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42541\,
            I => \current_shift_inst.un4_control_input1_23\
        );

    \I__9413\ : InMux
    port map (
            O => \N__42534\,
            I => \current_shift_inst.un4_control_input_1_cry_21\
        );

    \I__9412\ : InMux
    port map (
            O => \N__42531\,
            I => \N__42528\
        );

    \I__9411\ : LocalMux
    port map (
            O => \N__42528\,
            I => \N__42525\
        );

    \I__9410\ : Span4Mux_h
    port map (
            O => \N__42525\,
            I => \N__42522\
        );

    \I__9409\ : Odrv4
    port map (
            O => \N__42522\,
            I => \current_shift_inst.un4_control_input_1_axb_23\
        );

    \I__9408\ : InMux
    port map (
            O => \N__42519\,
            I => \N__42516\
        );

    \I__9407\ : LocalMux
    port map (
            O => \N__42516\,
            I => \N__42512\
        );

    \I__9406\ : InMux
    port map (
            O => \N__42515\,
            I => \N__42509\
        );

    \I__9405\ : Span4Mux_v
    port map (
            O => \N__42512\,
            I => \N__42505\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__42509\,
            I => \N__42502\
        );

    \I__9403\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42499\
        );

    \I__9402\ : Odrv4
    port map (
            O => \N__42505\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9401\ : Odrv4
    port map (
            O => \N__42502\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9400\ : LocalMux
    port map (
            O => \N__42499\,
            I => \current_shift_inst.un4_control_input1_24\
        );

    \I__9399\ : InMux
    port map (
            O => \N__42492\,
            I => \current_shift_inst.un4_control_input_1_cry_22\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42486\
        );

    \I__9397\ : LocalMux
    port map (
            O => \N__42486\,
            I => \N__42482\
        );

    \I__9396\ : InMux
    port map (
            O => \N__42485\,
            I => \N__42479\
        );

    \I__9395\ : Span4Mux_v
    port map (
            O => \N__42482\,
            I => \N__42473\
        );

    \I__9394\ : LocalMux
    port map (
            O => \N__42479\,
            I => \N__42473\
        );

    \I__9393\ : InMux
    port map (
            O => \N__42478\,
            I => \N__42470\
        );

    \I__9392\ : Odrv4
    port map (
            O => \N__42473\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__42470\,
            I => \current_shift_inst.un4_control_input1_25\
        );

    \I__9390\ : InMux
    port map (
            O => \N__42465\,
            I => \current_shift_inst.un4_control_input_1_cry_23\
        );

    \I__9389\ : InMux
    port map (
            O => \N__42462\,
            I => \bfn_17_18_0_\
        );

    \I__9388\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42454\
        );

    \I__9387\ : InMux
    port map (
            O => \N__42458\,
            I => \N__42451\
        );

    \I__9386\ : InMux
    port map (
            O => \N__42457\,
            I => \N__42448\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__42454\,
            I => \N__42445\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__42451\,
            I => \N__42442\
        );

    \I__9383\ : LocalMux
    port map (
            O => \N__42448\,
            I => \N__42439\
        );

    \I__9382\ : Span4Mux_h
    port map (
            O => \N__42445\,
            I => \N__42436\
        );

    \I__9381\ : Span4Mux_v
    port map (
            O => \N__42442\,
            I => \N__42431\
        );

    \I__9380\ : Span4Mux_h
    port map (
            O => \N__42439\,
            I => \N__42431\
        );

    \I__9379\ : Span4Mux_v
    port map (
            O => \N__42436\,
            I => \N__42428\
        );

    \I__9378\ : Odrv4
    port map (
            O => \N__42431\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9377\ : Odrv4
    port map (
            O => \N__42428\,
            I => \current_shift_inst.un4_control_input1_27\
        );

    \I__9376\ : InMux
    port map (
            O => \N__42423\,
            I => \current_shift_inst.un4_control_input_1_cry_25\
        );

    \I__9375\ : InMux
    port map (
            O => \N__42420\,
            I => \N__42415\
        );

    \I__9374\ : InMux
    port map (
            O => \N__42419\,
            I => \N__42412\
        );

    \I__9373\ : InMux
    port map (
            O => \N__42418\,
            I => \N__42409\
        );

    \I__9372\ : LocalMux
    port map (
            O => \N__42415\,
            I => \N__42406\
        );

    \I__9371\ : LocalMux
    port map (
            O => \N__42412\,
            I => \N__42401\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__42409\,
            I => \N__42401\
        );

    \I__9369\ : Span4Mux_v
    port map (
            O => \N__42406\,
            I => \N__42398\
        );

    \I__9368\ : Odrv4
    port map (
            O => \N__42401\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9367\ : Odrv4
    port map (
            O => \N__42398\,
            I => \current_shift_inst.un4_control_input1_28\
        );

    \I__9366\ : InMux
    port map (
            O => \N__42393\,
            I => \current_shift_inst.un4_control_input_1_cry_26\
        );

    \I__9365\ : InMux
    port map (
            O => \N__42390\,
            I => \N__42385\
        );

    \I__9364\ : InMux
    port map (
            O => \N__42389\,
            I => \N__42382\
        );

    \I__9363\ : InMux
    port map (
            O => \N__42388\,
            I => \N__42379\
        );

    \I__9362\ : LocalMux
    port map (
            O => \N__42385\,
            I => \N__42376\
        );

    \I__9361\ : LocalMux
    port map (
            O => \N__42382\,
            I => \N__42373\
        );

    \I__9360\ : LocalMux
    port map (
            O => \N__42379\,
            I => \N__42370\
        );

    \I__9359\ : Span4Mux_h
    port map (
            O => \N__42376\,
            I => \N__42367\
        );

    \I__9358\ : Span4Mux_h
    port map (
            O => \N__42373\,
            I => \N__42362\
        );

    \I__9357\ : Span4Mux_v
    port map (
            O => \N__42370\,
            I => \N__42362\
        );

    \I__9356\ : Odrv4
    port map (
            O => \N__42367\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9355\ : Odrv4
    port map (
            O => \N__42362\,
            I => \current_shift_inst.un4_control_input1_29\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42357\,
            I => \current_shift_inst.un4_control_input_1_cry_27\
        );

    \I__9353\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42349\
        );

    \I__9352\ : InMux
    port map (
            O => \N__42353\,
            I => \N__42346\
        );

    \I__9351\ : InMux
    port map (
            O => \N__42352\,
            I => \N__42343\
        );

    \I__9350\ : LocalMux
    port map (
            O => \N__42349\,
            I => \N__42340\
        );

    \I__9349\ : LocalMux
    port map (
            O => \N__42346\,
            I => \N__42337\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__42343\,
            I => \N__42334\
        );

    \I__9347\ : Span4Mux_v
    port map (
            O => \N__42340\,
            I => \N__42331\
        );

    \I__9346\ : Odrv4
    port map (
            O => \N__42337\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9345\ : Odrv4
    port map (
            O => \N__42334\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9344\ : Odrv4
    port map (
            O => \N__42331\,
            I => \current_shift_inst.un4_control_input1_30\
        );

    \I__9343\ : InMux
    port map (
            O => \N__42324\,
            I => \current_shift_inst.un4_control_input_1_cry_28\
        );

    \I__9342\ : InMux
    port map (
            O => \N__42321\,
            I => \current_shift_inst.un4_control_input1_31\
        );

    \I__9341\ : CascadeMux
    port map (
            O => \N__42318\,
            I => \N__42315\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42311\
        );

    \I__9339\ : InMux
    port map (
            O => \N__42314\,
            I => \N__42307\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__42311\,
            I => \N__42304\
        );

    \I__9337\ : InMux
    port map (
            O => \N__42310\,
            I => \N__42301\
        );

    \I__9336\ : LocalMux
    port map (
            O => \N__42307\,
            I => \N__42298\
        );

    \I__9335\ : Span4Mux_h
    port map (
            O => \N__42304\,
            I => \N__42295\
        );

    \I__9334\ : LocalMux
    port map (
            O => \N__42301\,
            I => \N__42292\
        );

    \I__9333\ : Sp12to4
    port map (
            O => \N__42298\,
            I => \N__42289\
        );

    \I__9332\ : Odrv4
    port map (
            O => \N__42295\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9331\ : Odrv4
    port map (
            O => \N__42292\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9330\ : Odrv12
    port map (
            O => \N__42289\,
            I => \current_shift_inst.un4_control_input1_31_THRU_CO\
        );

    \I__9329\ : InMux
    port map (
            O => \N__42282\,
            I => \current_shift_inst.un4_control_input_1_cry_13\
        );

    \I__9328\ : InMux
    port map (
            O => \N__42279\,
            I => \N__42275\
        );

    \I__9327\ : CascadeMux
    port map (
            O => \N__42278\,
            I => \N__42272\
        );

    \I__9326\ : LocalMux
    port map (
            O => \N__42275\,
            I => \N__42269\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42272\,
            I => \N__42265\
        );

    \I__9324\ : Span4Mux_h
    port map (
            O => \N__42269\,
            I => \N__42262\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42268\,
            I => \N__42259\
        );

    \I__9322\ : LocalMux
    port map (
            O => \N__42265\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9321\ : Odrv4
    port map (
            O => \N__42262\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9320\ : LocalMux
    port map (
            O => \N__42259\,
            I => \current_shift_inst.un4_control_input1_16\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42252\,
            I => \current_shift_inst.un4_control_input_1_cry_14\
        );

    \I__9318\ : InMux
    port map (
            O => \N__42249\,
            I => \N__42245\
        );

    \I__9317\ : CascadeMux
    port map (
            O => \N__42248\,
            I => \N__42242\
        );

    \I__9316\ : LocalMux
    port map (
            O => \N__42245\,
            I => \N__42239\
        );

    \I__9315\ : InMux
    port map (
            O => \N__42242\,
            I => \N__42236\
        );

    \I__9314\ : Span4Mux_v
    port map (
            O => \N__42239\,
            I => \N__42230\
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42236\,
            I => \N__42230\
        );

    \I__9312\ : InMux
    port map (
            O => \N__42235\,
            I => \N__42227\
        );

    \I__9311\ : Odrv4
    port map (
            O => \N__42230\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9310\ : LocalMux
    port map (
            O => \N__42227\,
            I => \current_shift_inst.un4_control_input1_17\
        );

    \I__9309\ : InMux
    port map (
            O => \N__42222\,
            I => \current_shift_inst.un4_control_input_1_cry_15\
        );

    \I__9308\ : InMux
    port map (
            O => \N__42219\,
            I => \N__42216\
        );

    \I__9307\ : LocalMux
    port map (
            O => \N__42216\,
            I => \current_shift_inst.un4_control_input_1_axb_17\
        );

    \I__9306\ : InMux
    port map (
            O => \N__42213\,
            I => \N__42208\
        );

    \I__9305\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42205\
        );

    \I__9304\ : InMux
    port map (
            O => \N__42211\,
            I => \N__42202\
        );

    \I__9303\ : LocalMux
    port map (
            O => \N__42208\,
            I => \N__42199\
        );

    \I__9302\ : LocalMux
    port map (
            O => \N__42205\,
            I => \N__42196\
        );

    \I__9301\ : LocalMux
    port map (
            O => \N__42202\,
            I => \N__42193\
        );

    \I__9300\ : Span4Mux_h
    port map (
            O => \N__42199\,
            I => \N__42188\
        );

    \I__9299\ : Span4Mux_v
    port map (
            O => \N__42196\,
            I => \N__42188\
        );

    \I__9298\ : Odrv12
    port map (
            O => \N__42193\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9297\ : Odrv4
    port map (
            O => \N__42188\,
            I => \current_shift_inst.un4_control_input1_18\
        );

    \I__9296\ : InMux
    port map (
            O => \N__42183\,
            I => \bfn_17_17_0_\
        );

    \I__9295\ : CascadeMux
    port map (
            O => \N__42180\,
            I => \N__42177\
        );

    \I__9294\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42172\
        );

    \I__9293\ : InMux
    port map (
            O => \N__42176\,
            I => \N__42169\
        );

    \I__9292\ : InMux
    port map (
            O => \N__42175\,
            I => \N__42166\
        );

    \I__9291\ : LocalMux
    port map (
            O => \N__42172\,
            I => \N__42163\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__42169\,
            I => \N__42160\
        );

    \I__9289\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42157\
        );

    \I__9288\ : Span4Mux_h
    port map (
            O => \N__42163\,
            I => \N__42152\
        );

    \I__9287\ : Span4Mux_v
    port map (
            O => \N__42160\,
            I => \N__42152\
        );

    \I__9286\ : Span4Mux_v
    port map (
            O => \N__42157\,
            I => \N__42149\
        );

    \I__9285\ : Odrv4
    port map (
            O => \N__42152\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9284\ : Odrv4
    port map (
            O => \N__42149\,
            I => \current_shift_inst.un4_control_input1_19\
        );

    \I__9283\ : InMux
    port map (
            O => \N__42144\,
            I => \current_shift_inst.un4_control_input_1_cry_17\
        );

    \I__9282\ : CascadeMux
    port map (
            O => \N__42141\,
            I => \N__42137\
        );

    \I__9281\ : InMux
    port map (
            O => \N__42140\,
            I => \N__42133\
        );

    \I__9280\ : InMux
    port map (
            O => \N__42137\,
            I => \N__42130\
        );

    \I__9279\ : InMux
    port map (
            O => \N__42136\,
            I => \N__42127\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__42133\,
            I => \N__42124\
        );

    \I__9277\ : LocalMux
    port map (
            O => \N__42130\,
            I => \N__42121\
        );

    \I__9276\ : LocalMux
    port map (
            O => \N__42127\,
            I => \N__42118\
        );

    \I__9275\ : Span4Mux_h
    port map (
            O => \N__42124\,
            I => \N__42113\
        );

    \I__9274\ : Span4Mux_v
    port map (
            O => \N__42121\,
            I => \N__42113\
        );

    \I__9273\ : Span4Mux_v
    port map (
            O => \N__42118\,
            I => \N__42110\
        );

    \I__9272\ : Odrv4
    port map (
            O => \N__42113\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9271\ : Odrv4
    port map (
            O => \N__42110\,
            I => \current_shift_inst.un4_control_input1_20\
        );

    \I__9270\ : InMux
    port map (
            O => \N__42105\,
            I => \current_shift_inst.un4_control_input_1_cry_18\
        );

    \I__9269\ : InMux
    port map (
            O => \N__42102\,
            I => \current_shift_inst.un4_control_input_1_cry_19\
        );

    \I__9268\ : InMux
    port map (
            O => \N__42099\,
            I => \N__42096\
        );

    \I__9267\ : LocalMux
    port map (
            O => \N__42096\,
            I => \current_shift_inst.un4_control_input_1_axb_21\
        );

    \I__9266\ : CascadeMux
    port map (
            O => \N__42093\,
            I => \N__42090\
        );

    \I__9265\ : InMux
    port map (
            O => \N__42090\,
            I => \N__42086\
        );

    \I__9264\ : InMux
    port map (
            O => \N__42089\,
            I => \N__42082\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__42086\,
            I => \N__42079\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42085\,
            I => \N__42076\
        );

    \I__9261\ : LocalMux
    port map (
            O => \N__42082\,
            I => \N__42073\
        );

    \I__9260\ : Span4Mux_h
    port map (
            O => \N__42079\,
            I => \N__42068\
        );

    \I__9259\ : LocalMux
    port map (
            O => \N__42076\,
            I => \N__42068\
        );

    \I__9258\ : Span4Mux_v
    port map (
            O => \N__42073\,
            I => \N__42065\
        );

    \I__9257\ : Odrv4
    port map (
            O => \N__42068\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9256\ : Odrv4
    port map (
            O => \N__42065\,
            I => \current_shift_inst.un4_control_input1_22\
        );

    \I__9255\ : InMux
    port map (
            O => \N__42060\,
            I => \current_shift_inst.un4_control_input_1_cry_20\
        );

    \I__9254\ : InMux
    port map (
            O => \N__42057\,
            I => \current_shift_inst.un4_control_input_1_cry_4\
        );

    \I__9253\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42050\
        );

    \I__9252\ : InMux
    port map (
            O => \N__42053\,
            I => \N__42047\
        );

    \I__9251\ : LocalMux
    port map (
            O => \N__42050\,
            I => \N__42044\
        );

    \I__9250\ : LocalMux
    port map (
            O => \N__42047\,
            I => \N__42041\
        );

    \I__9249\ : Span4Mux_v
    port map (
            O => \N__42044\,
            I => \N__42037\
        );

    \I__9248\ : Span4Mux_h
    port map (
            O => \N__42041\,
            I => \N__42034\
        );

    \I__9247\ : InMux
    port map (
            O => \N__42040\,
            I => \N__42031\
        );

    \I__9246\ : Odrv4
    port map (
            O => \N__42037\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9245\ : Odrv4
    port map (
            O => \N__42034\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__42031\,
            I => \current_shift_inst.un4_control_input1_7\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42024\,
            I => \current_shift_inst.un4_control_input_1_cry_5\
        );

    \I__9242\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42018\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42018\,
            I => \N__42015\
        );

    \I__9240\ : Span4Mux_h
    port map (
            O => \N__42015\,
            I => \N__42012\
        );

    \I__9239\ : Odrv4
    port map (
            O => \N__42012\,
            I => \current_shift_inst.un4_control_input_1_axb_7\
        );

    \I__9238\ : InMux
    port map (
            O => \N__42009\,
            I => \N__42005\
        );

    \I__9237\ : InMux
    port map (
            O => \N__42008\,
            I => \N__42002\
        );

    \I__9236\ : LocalMux
    port map (
            O => \N__42005\,
            I => \N__41999\
        );

    \I__9235\ : LocalMux
    port map (
            O => \N__42002\,
            I => \N__41996\
        );

    \I__9234\ : Span4Mux_h
    port map (
            O => \N__41999\,
            I => \N__41992\
        );

    \I__9233\ : Span4Mux_h
    port map (
            O => \N__41996\,
            I => \N__41989\
        );

    \I__9232\ : InMux
    port map (
            O => \N__41995\,
            I => \N__41986\
        );

    \I__9231\ : Odrv4
    port map (
            O => \N__41992\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9230\ : Odrv4
    port map (
            O => \N__41989\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9229\ : LocalMux
    port map (
            O => \N__41986\,
            I => \current_shift_inst.un4_control_input1_8\
        );

    \I__9228\ : InMux
    port map (
            O => \N__41979\,
            I => \current_shift_inst.un4_control_input_1_cry_6\
        );

    \I__9227\ : InMux
    port map (
            O => \N__41976\,
            I => \N__41973\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__41973\,
            I => \N__41969\
        );

    \I__9225\ : InMux
    port map (
            O => \N__41972\,
            I => \N__41966\
        );

    \I__9224\ : Span4Mux_v
    port map (
            O => \N__41969\,
            I => \N__41960\
        );

    \I__9223\ : LocalMux
    port map (
            O => \N__41966\,
            I => \N__41960\
        );

    \I__9222\ : InMux
    port map (
            O => \N__41965\,
            I => \N__41957\
        );

    \I__9221\ : Odrv4
    port map (
            O => \N__41960\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9220\ : LocalMux
    port map (
            O => \N__41957\,
            I => \current_shift_inst.un4_control_input1_9\
        );

    \I__9219\ : InMux
    port map (
            O => \N__41952\,
            I => \current_shift_inst.un4_control_input_1_cry_7\
        );

    \I__9218\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41946\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__41946\,
            I => \current_shift_inst.un4_control_input_1_axb_9\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__9215\ : LocalMux
    port map (
            O => \N__41940\,
            I => \N__41937\
        );

    \I__9214\ : Span4Mux_v
    port map (
            O => \N__41937\,
            I => \N__41932\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41936\,
            I => \N__41929\
        );

    \I__9212\ : InMux
    port map (
            O => \N__41935\,
            I => \N__41926\
        );

    \I__9211\ : Odrv4
    port map (
            O => \N__41932\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41929\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9209\ : LocalMux
    port map (
            O => \N__41926\,
            I => \current_shift_inst.un4_control_input1_10\
        );

    \I__9208\ : InMux
    port map (
            O => \N__41919\,
            I => \bfn_17_16_0_\
        );

    \I__9207\ : InMux
    port map (
            O => \N__41916\,
            I => \N__41913\
        );

    \I__9206\ : LocalMux
    port map (
            O => \N__41913\,
            I => \current_shift_inst.un4_control_input_1_axb_10\
        );

    \I__9205\ : InMux
    port map (
            O => \N__41910\,
            I => \current_shift_inst.un4_control_input_1_cry_9\
        );

    \I__9204\ : InMux
    port map (
            O => \N__41907\,
            I => \N__41904\
        );

    \I__9203\ : LocalMux
    port map (
            O => \N__41904\,
            I => \current_shift_inst.un4_control_input_1_axb_11\
        );

    \I__9202\ : InMux
    port map (
            O => \N__41901\,
            I => \current_shift_inst.un4_control_input_1_cry_10\
        );

    \I__9201\ : InMux
    port map (
            O => \N__41898\,
            I => \current_shift_inst.un4_control_input_1_cry_11\
        );

    \I__9200\ : InMux
    port map (
            O => \N__41895\,
            I => \current_shift_inst.un4_control_input_1_cry_12\
        );

    \I__9199\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41889\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__41889\,
            I => \current_shift_inst.un4_control_input1_1\
        );

    \I__9197\ : CascadeMux
    port map (
            O => \N__41886\,
            I => \current_shift_inst.un4_control_input1_1_cascade_\
        );

    \I__9196\ : CascadeMux
    port map (
            O => \N__41883\,
            I => \N__41879\
        );

    \I__9195\ : InMux
    port map (
            O => \N__41882\,
            I => \N__41876\
        );

    \I__9194\ : InMux
    port map (
            O => \N__41879\,
            I => \N__41873\
        );

    \I__9193\ : LocalMux
    port map (
            O => \N__41876\,
            I => \N__41870\
        );

    \I__9192\ : LocalMux
    port map (
            O => \N__41873\,
            I => \N__41867\
        );

    \I__9191\ : Span4Mux_h
    port map (
            O => \N__41870\,
            I => \N__41864\
        );

    \I__9190\ : Span4Mux_h
    port map (
            O => \N__41867\,
            I => \N__41861\
        );

    \I__9189\ : Span4Mux_v
    port map (
            O => \N__41864\,
            I => \N__41856\
        );

    \I__9188\ : Span4Mux_h
    port map (
            O => \N__41861\,
            I => \N__41856\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__41856\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\
        );

    \I__9186\ : CascadeMux
    port map (
            O => \N__41853\,
            I => \N__41850\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41850\,
            I => \N__41847\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__9183\ : Span4Mux_h
    port map (
            O => \N__41844\,
            I => \N__41841\
        );

    \I__9182\ : Odrv4
    port map (
            O => \N__41841\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\
        );

    \I__9181\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41833\
        );

    \I__9180\ : InMux
    port map (
            O => \N__41837\,
            I => \N__41828\
        );

    \I__9179\ : InMux
    port map (
            O => \N__41836\,
            I => \N__41828\
        );

    \I__9178\ : LocalMux
    port map (
            O => \N__41833\,
            I => \N__41824\
        );

    \I__9177\ : LocalMux
    port map (
            O => \N__41828\,
            I => \N__41821\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41827\,
            I => \N__41818\
        );

    \I__9175\ : Span4Mux_v
    port map (
            O => \N__41824\,
            I => \N__41815\
        );

    \I__9174\ : Span4Mux_v
    port map (
            O => \N__41821\,
            I => \N__41812\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__41818\,
            I => \N__41809\
        );

    \I__9172\ : Odrv4
    port map (
            O => \N__41815\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9171\ : Odrv4
    port map (
            O => \N__41812\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9170\ : Odrv4
    port map (
            O => \N__41809\,
            I => \current_shift_inst.elapsed_time_ns_s1_5\
        );

    \I__9169\ : CascadeMux
    port map (
            O => \N__41802\,
            I => \N__41799\
        );

    \I__9168\ : InMux
    port map (
            O => \N__41799\,
            I => \N__41796\
        );

    \I__9167\ : LocalMux
    port map (
            O => \N__41796\,
            I => \N__41793\
        );

    \I__9166\ : Span4Mux_h
    port map (
            O => \N__41793\,
            I => \N__41790\
        );

    \I__9165\ : Odrv4
    port map (
            O => \N__41790\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41784\
        );

    \I__9163\ : LocalMux
    port map (
            O => \N__41784\,
            I => \N__41781\
        );

    \I__9162\ : Odrv4
    port map (
            O => \N__41781\,
            I => \current_shift_inst.un4_control_input_1_axb_2\
        );

    \I__9161\ : InMux
    port map (
            O => \N__41778\,
            I => \N__41775\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41775\,
            I => \N__41771\
        );

    \I__9159\ : InMux
    port map (
            O => \N__41774\,
            I => \N__41768\
        );

    \I__9158\ : Span4Mux_v
    port map (
            O => \N__41771\,
            I => \N__41762\
        );

    \I__9157\ : LocalMux
    port map (
            O => \N__41768\,
            I => \N__41762\
        );

    \I__9156\ : InMux
    port map (
            O => \N__41767\,
            I => \N__41759\
        );

    \I__9155\ : Odrv4
    port map (
            O => \N__41762\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__41759\,
            I => \current_shift_inst.un4_control_input1_3\
        );

    \I__9153\ : InMux
    port map (
            O => \N__41754\,
            I => \current_shift_inst.un4_control_input_1_cry_1\
        );

    \I__9152\ : InMux
    port map (
            O => \N__41751\,
            I => \N__41748\
        );

    \I__9151\ : LocalMux
    port map (
            O => \N__41748\,
            I => \N__41745\
        );

    \I__9150\ : Span4Mux_v
    port map (
            O => \N__41745\,
            I => \N__41740\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41737\
        );

    \I__9148\ : InMux
    port map (
            O => \N__41743\,
            I => \N__41734\
        );

    \I__9147\ : Odrv4
    port map (
            O => \N__41740\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__41737\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9145\ : LocalMux
    port map (
            O => \N__41734\,
            I => \current_shift_inst.un4_control_input1_4\
        );

    \I__9144\ : InMux
    port map (
            O => \N__41727\,
            I => \current_shift_inst.un4_control_input_1_cry_2\
        );

    \I__9143\ : InMux
    port map (
            O => \N__41724\,
            I => \N__41721\
        );

    \I__9142\ : LocalMux
    port map (
            O => \N__41721\,
            I => \current_shift_inst.un4_control_input_1_axb_4\
        );

    \I__9141\ : InMux
    port map (
            O => \N__41718\,
            I => \N__41713\
        );

    \I__9140\ : InMux
    port map (
            O => \N__41717\,
            I => \N__41708\
        );

    \I__9139\ : InMux
    port map (
            O => \N__41716\,
            I => \N__41708\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41713\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__41708\,
            I => \current_shift_inst.un4_control_input1_5\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41703\,
            I => \current_shift_inst.un4_control_input_1_cry_3\
        );

    \I__9135\ : CascadeMux
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__9134\ : InMux
    port map (
            O => \N__41697\,
            I => \N__41692\
        );

    \I__9133\ : InMux
    port map (
            O => \N__41696\,
            I => \N__41687\
        );

    \I__9132\ : InMux
    port map (
            O => \N__41695\,
            I => \N__41687\
        );

    \I__9131\ : LocalMux
    port map (
            O => \N__41692\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9130\ : LocalMux
    port map (
            O => \N__41687\,
            I => \current_shift_inst.un4_control_input1_6\
        );

    \I__9129\ : InMux
    port map (
            O => \N__41682\,
            I => \N__41679\
        );

    \I__9128\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41673\
        );

    \I__9127\ : InMux
    port map (
            O => \N__41678\,
            I => \N__41670\
        );

    \I__9126\ : InMux
    port map (
            O => \N__41677\,
            I => \N__41665\
        );

    \I__9125\ : InMux
    port map (
            O => \N__41676\,
            I => \N__41665\
        );

    \I__9124\ : Span4Mux_h
    port map (
            O => \N__41673\,
            I => \N__41662\
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__41670\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__41665\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9121\ : Odrv4
    port map (
            O => \N__41662\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\
        );

    \I__9120\ : InMux
    port map (
            O => \N__41655\,
            I => \N__41652\
        );

    \I__9119\ : LocalMux
    port map (
            O => \N__41652\,
            I => \N__41648\
        );

    \I__9118\ : InMux
    port map (
            O => \N__41651\,
            I => \N__41645\
        );

    \I__9117\ : Odrv4
    port map (
            O => \N__41648\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__9116\ : LocalMux
    port map (
            O => \N__41645\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22\
        );

    \I__9115\ : InMux
    port map (
            O => \N__41640\,
            I => \N__41634\
        );

    \I__9114\ : InMux
    port map (
            O => \N__41639\,
            I => \N__41634\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__41634\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\
        );

    \I__9112\ : InMux
    port map (
            O => \N__41631\,
            I => \N__41625\
        );

    \I__9111\ : InMux
    port map (
            O => \N__41630\,
            I => \N__41625\
        );

    \I__9110\ : LocalMux
    port map (
            O => \N__41625\,
            I => \N__41620\
        );

    \I__9109\ : InMux
    port map (
            O => \N__41624\,
            I => \N__41617\
        );

    \I__9108\ : InMux
    port map (
            O => \N__41623\,
            I => \N__41614\
        );

    \I__9107\ : Span4Mux_v
    port map (
            O => \N__41620\,
            I => \N__41609\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__41617\,
            I => \N__41609\
        );

    \I__9105\ : LocalMux
    port map (
            O => \N__41614\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9104\ : Odrv4
    port map (
            O => \N__41609\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\
        );

    \I__9103\ : InMux
    port map (
            O => \N__41604\,
            I => \N__41601\
        );

    \I__9102\ : LocalMux
    port map (
            O => \N__41601\,
            I => \N__41598\
        );

    \I__9101\ : Span4Mux_h
    port map (
            O => \N__41598\,
            I => \N__41594\
        );

    \I__9100\ : InMux
    port map (
            O => \N__41597\,
            I => \N__41591\
        );

    \I__9099\ : Odrv4
    port map (
            O => \N__41594\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9098\ : LocalMux
    port map (
            O => \N__41591\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26\
        );

    \I__9097\ : InMux
    port map (
            O => \N__41586\,
            I => \N__41582\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41579\
        );

    \I__9095\ : LocalMux
    port map (
            O => \N__41582\,
            I => \N__41576\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41579\,
            I => \N__41570\
        );

    \I__9093\ : Sp12to4
    port map (
            O => \N__41576\,
            I => \N__41570\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41567\
        );

    \I__9091\ : Span12Mux_s10_h
    port map (
            O => \N__41570\,
            I => \N__41564\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__41567\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__9089\ : Odrv12
    port map (
            O => \N__41564\,
            I => \elapsed_time_ns_1_RNI14DN9_0_23\
        );

    \I__9088\ : InMux
    port map (
            O => \N__41559\,
            I => \N__41555\
        );

    \I__9087\ : InMux
    port map (
            O => \N__41558\,
            I => \N__41552\
        );

    \I__9086\ : LocalMux
    port map (
            O => \N__41555\,
            I => \N__41547\
        );

    \I__9085\ : LocalMux
    port map (
            O => \N__41552\,
            I => \N__41544\
        );

    \I__9084\ : InMux
    port map (
            O => \N__41551\,
            I => \N__41541\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41550\,
            I => \N__41538\
        );

    \I__9082\ : Span4Mux_v
    port map (
            O => \N__41547\,
            I => \N__41533\
        );

    \I__9081\ : Span4Mux_h
    port map (
            O => \N__41544\,
            I => \N__41533\
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__41541\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__41538\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9078\ : Odrv4
    port map (
            O => \N__41533\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41522\
        );

    \I__9076\ : InMux
    port map (
            O => \N__41525\,
            I => \N__41519\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__41522\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41519\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\
        );

    \I__9073\ : InMux
    port map (
            O => \N__41514\,
            I => \N__41510\
        );

    \I__9072\ : InMux
    port map (
            O => \N__41513\,
            I => \N__41506\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__41510\,
            I => \N__41503\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41509\,
            I => \N__41500\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__41506\,
            I => \N__41497\
        );

    \I__9068\ : Span4Mux_v
    port map (
            O => \N__41503\,
            I => \N__41493\
        );

    \I__9067\ : LocalMux
    port map (
            O => \N__41500\,
            I => \N__41490\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__41497\,
            I => \N__41487\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41496\,
            I => \N__41484\
        );

    \I__9064\ : Odrv4
    port map (
            O => \N__41493\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9063\ : Odrv4
    port map (
            O => \N__41490\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9062\ : Odrv4
    port map (
            O => \N__41487\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__41484\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\
        );

    \I__9060\ : InMux
    port map (
            O => \N__41475\,
            I => \N__41471\
        );

    \I__9059\ : InMux
    port map (
            O => \N__41474\,
            I => \N__41468\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41471\,
            I => \N__41465\
        );

    \I__9057\ : LocalMux
    port map (
            O => \N__41468\,
            I => \N__41462\
        );

    \I__9056\ : Span4Mux_h
    port map (
            O => \N__41465\,
            I => \N__41456\
        );

    \I__9055\ : Span4Mux_v
    port map (
            O => \N__41462\,
            I => \N__41456\
        );

    \I__9054\ : InMux
    port map (
            O => \N__41461\,
            I => \N__41453\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__41456\,
            I => \N__41450\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41453\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__9051\ : Odrv4
    port map (
            O => \N__41450\,
            I => \elapsed_time_ns_1_RNIF13T9_0_3\
        );

    \I__9050\ : CascadeMux
    port map (
            O => \N__41445\,
            I => \N__41442\
        );

    \I__9049\ : InMux
    port map (
            O => \N__41442\,
            I => \N__41439\
        );

    \I__9048\ : LocalMux
    port map (
            O => \N__41439\,
            I => \N__41436\
        );

    \I__9047\ : Odrv12
    port map (
            O => \N__41436\,
            I => \current_shift_inst.un38_control_input_cry_0_s0_sf\
        );

    \I__9046\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41427\
        );

    \I__9045\ : InMux
    port map (
            O => \N__41432\,
            I => \N__41424\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41431\,
            I => \N__41421\
        );

    \I__9043\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41418\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41413\
        );

    \I__9041\ : LocalMux
    port map (
            O => \N__41424\,
            I => \N__41413\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__41421\,
            I => \N__41408\
        );

    \I__9039\ : LocalMux
    port map (
            O => \N__41418\,
            I => \N__41408\
        );

    \I__9038\ : Span4Mux_v
    port map (
            O => \N__41413\,
            I => \N__41405\
        );

    \I__9037\ : Odrv4
    port map (
            O => \N__41408\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9036\ : Odrv4
    port map (
            O => \N__41405\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\
        );

    \I__9035\ : InMux
    port map (
            O => \N__41400\,
            I => \N__41397\
        );

    \I__9034\ : LocalMux
    port map (
            O => \N__41397\,
            I => \N__41392\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41396\,
            I => \N__41389\
        );

    \I__9032\ : InMux
    port map (
            O => \N__41395\,
            I => \N__41386\
        );

    \I__9031\ : Span4Mux_h
    port map (
            O => \N__41392\,
            I => \N__41383\
        );

    \I__9030\ : LocalMux
    port map (
            O => \N__41389\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__9029\ : LocalMux
    port map (
            O => \N__41386\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__9028\ : Odrv4
    port map (
            O => \N__41383\,
            I => \elapsed_time_ns_1_RNIL73T9_0_9\
        );

    \I__9027\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41371\
        );

    \I__9026\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41368\
        );

    \I__9025\ : InMux
    port map (
            O => \N__41374\,
            I => \N__41364\
        );

    \I__9024\ : LocalMux
    port map (
            O => \N__41371\,
            I => \N__41359\
        );

    \I__9023\ : LocalMux
    port map (
            O => \N__41368\,
            I => \N__41359\
        );

    \I__9022\ : InMux
    port map (
            O => \N__41367\,
            I => \N__41356\
        );

    \I__9021\ : LocalMux
    port map (
            O => \N__41364\,
            I => \N__41353\
        );

    \I__9020\ : Span4Mux_v
    port map (
            O => \N__41359\,
            I => \N__41350\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__41356\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9018\ : Odrv4
    port map (
            O => \N__41353\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9017\ : Odrv4
    port map (
            O => \N__41350\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41343\,
            I => \N__41338\
        );

    \I__9015\ : InMux
    port map (
            O => \N__41342\,
            I => \N__41335\
        );

    \I__9014\ : InMux
    port map (
            O => \N__41341\,
            I => \N__41332\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41338\,
            I => \N__41329\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__41335\,
            I => \N__41326\
        );

    \I__9011\ : LocalMux
    port map (
            O => \N__41332\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__9010\ : Odrv12
    port map (
            O => \N__41329\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__9009\ : Odrv4
    port map (
            O => \N__41326\,
            I => \elapsed_time_ns_1_RNIV0CN9_0_12\
        );

    \I__9008\ : CascadeMux
    port map (
            O => \N__41319\,
            I => \N__41315\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41318\,
            I => \N__41312\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41315\,
            I => \N__41309\
        );

    \I__9005\ : LocalMux
    port map (
            O => \N__41312\,
            I => \N__41305\
        );

    \I__9004\ : LocalMux
    port map (
            O => \N__41309\,
            I => \N__41302\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41308\,
            I => \N__41299\
        );

    \I__9002\ : Span4Mux_v
    port map (
            O => \N__41305\,
            I => \N__41294\
        );

    \I__9001\ : Span4Mux_h
    port map (
            O => \N__41302\,
            I => \N__41294\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41299\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8999\ : Odrv4
    port map (
            O => \N__41294\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__8998\ : InMux
    port map (
            O => \N__41289\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__8997\ : IoInMux
    port map (
            O => \N__41286\,
            I => \N__41283\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__41283\,
            I => \N__41280\
        );

    \I__8995\ : IoSpan4Mux
    port map (
            O => \N__41280\,
            I => \N__41266\
        );

    \I__8994\ : InMux
    port map (
            O => \N__41279\,
            I => \N__41254\
        );

    \I__8993\ : InMux
    port map (
            O => \N__41278\,
            I => \N__41254\
        );

    \I__8992\ : InMux
    port map (
            O => \N__41277\,
            I => \N__41254\
        );

    \I__8991\ : InMux
    port map (
            O => \N__41276\,
            I => \N__41254\
        );

    \I__8990\ : InMux
    port map (
            O => \N__41275\,
            I => \N__41235\
        );

    \I__8989\ : InMux
    port map (
            O => \N__41274\,
            I => \N__41235\
        );

    \I__8988\ : InMux
    port map (
            O => \N__41273\,
            I => \N__41235\
        );

    \I__8987\ : InMux
    port map (
            O => \N__41272\,
            I => \N__41226\
        );

    \I__8986\ : InMux
    port map (
            O => \N__41271\,
            I => \N__41226\
        );

    \I__8985\ : InMux
    port map (
            O => \N__41270\,
            I => \N__41226\
        );

    \I__8984\ : InMux
    port map (
            O => \N__41269\,
            I => \N__41226\
        );

    \I__8983\ : Sp12to4
    port map (
            O => \N__41266\,
            I => \N__41223\
        );

    \I__8982\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41216\
        );

    \I__8981\ : InMux
    port map (
            O => \N__41264\,
            I => \N__41216\
        );

    \I__8980\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41216\
        );

    \I__8979\ : LocalMux
    port map (
            O => \N__41254\,
            I => \N__41208\
        );

    \I__8978\ : InMux
    port map (
            O => \N__41253\,
            I => \N__41199\
        );

    \I__8977\ : InMux
    port map (
            O => \N__41252\,
            I => \N__41199\
        );

    \I__8976\ : InMux
    port map (
            O => \N__41251\,
            I => \N__41199\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41250\,
            I => \N__41199\
        );

    \I__8974\ : InMux
    port map (
            O => \N__41249\,
            I => \N__41190\
        );

    \I__8973\ : InMux
    port map (
            O => \N__41248\,
            I => \N__41190\
        );

    \I__8972\ : InMux
    port map (
            O => \N__41247\,
            I => \N__41190\
        );

    \I__8971\ : InMux
    port map (
            O => \N__41246\,
            I => \N__41190\
        );

    \I__8970\ : InMux
    port map (
            O => \N__41245\,
            I => \N__41181\
        );

    \I__8969\ : InMux
    port map (
            O => \N__41244\,
            I => \N__41181\
        );

    \I__8968\ : InMux
    port map (
            O => \N__41243\,
            I => \N__41181\
        );

    \I__8967\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41181\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__41235\,
            I => \N__41178\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__41226\,
            I => \N__41175\
        );

    \I__8964\ : Span12Mux_v
    port map (
            O => \N__41223\,
            I => \N__41172\
        );

    \I__8963\ : LocalMux
    port map (
            O => \N__41216\,
            I => \N__41169\
        );

    \I__8962\ : InMux
    port map (
            O => \N__41215\,
            I => \N__41166\
        );

    \I__8961\ : InMux
    port map (
            O => \N__41214\,
            I => \N__41157\
        );

    \I__8960\ : InMux
    port map (
            O => \N__41213\,
            I => \N__41157\
        );

    \I__8959\ : InMux
    port map (
            O => \N__41212\,
            I => \N__41157\
        );

    \I__8958\ : InMux
    port map (
            O => \N__41211\,
            I => \N__41157\
        );

    \I__8957\ : Span4Mux_h
    port map (
            O => \N__41208\,
            I => \N__41144\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__41199\,
            I => \N__41144\
        );

    \I__8955\ : LocalMux
    port map (
            O => \N__41190\,
            I => \N__41144\
        );

    \I__8954\ : LocalMux
    port map (
            O => \N__41181\,
            I => \N__41144\
        );

    \I__8953\ : Span4Mux_v
    port map (
            O => \N__41178\,
            I => \N__41144\
        );

    \I__8952\ : Span4Mux_v
    port map (
            O => \N__41175\,
            I => \N__41144\
        );

    \I__8951\ : Span12Mux_v
    port map (
            O => \N__41172\,
            I => \N__41141\
        );

    \I__8950\ : Odrv4
    port map (
            O => \N__41169\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8949\ : LocalMux
    port map (
            O => \N__41166\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__41157\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__41144\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8946\ : Odrv12
    port map (
            O => \N__41141\,
            I => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41130\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__41127\,
            I => \N__41124\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41124\,
            I => \N__41121\
        );

    \I__8942\ : LocalMux
    port map (
            O => \N__41121\,
            I => \N__41116\
        );

    \I__8941\ : InMux
    port map (
            O => \N__41120\,
            I => \N__41113\
        );

    \I__8940\ : InMux
    port map (
            O => \N__41119\,
            I => \N__41110\
        );

    \I__8939\ : Span4Mux_h
    port map (
            O => \N__41116\,
            I => \N__41107\
        );

    \I__8938\ : LocalMux
    port map (
            O => \N__41113\,
            I => \N__41104\
        );

    \I__8937\ : LocalMux
    port map (
            O => \N__41110\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8936\ : Odrv4
    port map (
            O => \N__41107\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8935\ : Odrv12
    port map (
            O => \N__41104\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__8934\ : CascadeMux
    port map (
            O => \N__41097\,
            I => \N__41094\
        );

    \I__8933\ : InMux
    port map (
            O => \N__41094\,
            I => \N__41091\
        );

    \I__8932\ : LocalMux
    port map (
            O => \N__41091\,
            I => \N__41088\
        );

    \I__8931\ : Span4Mux_h
    port map (
            O => \N__41088\,
            I => \N__41085\
        );

    \I__8930\ : Odrv4
    port map (
            O => \N__41085\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt22\
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__41082\,
            I => \N__41078\
        );

    \I__8928\ : InMux
    port map (
            O => \N__41081\,
            I => \N__41072\
        );

    \I__8927\ : InMux
    port map (
            O => \N__41078\,
            I => \N__41072\
        );

    \I__8926\ : InMux
    port map (
            O => \N__41077\,
            I => \N__41069\
        );

    \I__8925\ : LocalMux
    port map (
            O => \N__41072\,
            I => \N__41066\
        );

    \I__8924\ : LocalMux
    port map (
            O => \N__41069\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8923\ : Odrv4
    port map (
            O => \N__41066\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__8922\ : CascadeMux
    port map (
            O => \N__41061\,
            I => \N__41058\
        );

    \I__8921\ : InMux
    port map (
            O => \N__41058\,
            I => \N__41053\
        );

    \I__8920\ : InMux
    port map (
            O => \N__41057\,
            I => \N__41050\
        );

    \I__8919\ : InMux
    port map (
            O => \N__41056\,
            I => \N__41047\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41053\,
            I => \N__41042\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__41050\,
            I => \N__41042\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__41047\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8915\ : Odrv4
    port map (
            O => \N__41042\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__8914\ : InMux
    port map (
            O => \N__41037\,
            I => \N__41034\
        );

    \I__8913\ : LocalMux
    port map (
            O => \N__41034\,
            I => \N__41031\
        );

    \I__8912\ : Odrv4
    port map (
            O => \N__41031\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\
        );

    \I__8911\ : InMux
    port map (
            O => \N__41028\,
            I => \N__41025\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__41025\,
            I => \N__41020\
        );

    \I__8909\ : InMux
    port map (
            O => \N__41024\,
            I => \N__41017\
        );

    \I__8908\ : InMux
    port map (
            O => \N__41023\,
            I => \N__41014\
        );

    \I__8907\ : Span4Mux_h
    port map (
            O => \N__41020\,
            I => \N__41011\
        );

    \I__8906\ : LocalMux
    port map (
            O => \N__41017\,
            I => \N__41008\
        );

    \I__8905\ : LocalMux
    port map (
            O => \N__41014\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__8904\ : Odrv4
    port map (
            O => \N__41011\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__8903\ : Odrv4
    port map (
            O => \N__41008\,
            I => \elapsed_time_ns_1_RNITUBN9_0_10\
        );

    \I__8902\ : InMux
    port map (
            O => \N__41001\,
            I => \N__40998\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__40998\,
            I => \N__40993\
        );

    \I__8900\ : InMux
    port map (
            O => \N__40997\,
            I => \N__40988\
        );

    \I__8899\ : InMux
    port map (
            O => \N__40996\,
            I => \N__40988\
        );

    \I__8898\ : Span4Mux_h
    port map (
            O => \N__40993\,
            I => \N__40982\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__40988\,
            I => \N__40982\
        );

    \I__8896\ : InMux
    port map (
            O => \N__40987\,
            I => \N__40979\
        );

    \I__8895\ : Span4Mux_v
    port map (
            O => \N__40982\,
            I => \N__40976\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__40979\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8893\ : Odrv4
    port map (
            O => \N__40976\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\
        );

    \I__8892\ : InMux
    port map (
            O => \N__40971\,
            I => \N__40968\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__40968\,
            I => \N__40965\
        );

    \I__8890\ : Odrv4
    port map (
            O => \N__40965\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\
        );

    \I__8889\ : CascadeMux
    port map (
            O => \N__40962\,
            I => \N__40957\
        );

    \I__8888\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40954\
        );

    \I__8887\ : InMux
    port map (
            O => \N__40960\,
            I => \N__40951\
        );

    \I__8886\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40948\
        );

    \I__8885\ : LocalMux
    port map (
            O => \N__40954\,
            I => \N__40940\
        );

    \I__8884\ : LocalMux
    port map (
            O => \N__40951\,
            I => \N__40940\
        );

    \I__8883\ : LocalMux
    port map (
            O => \N__40948\,
            I => \N__40940\
        );

    \I__8882\ : InMux
    port map (
            O => \N__40947\,
            I => \N__40937\
        );

    \I__8881\ : Span4Mux_v
    port map (
            O => \N__40940\,
            I => \N__40934\
        );

    \I__8880\ : LocalMux
    port map (
            O => \N__40937\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__8879\ : Odrv4
    port map (
            O => \N__40934\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\
        );

    \I__8878\ : InMux
    port map (
            O => \N__40929\,
            I => \N__40926\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__40926\,
            I => \N__40922\
        );

    \I__8876\ : InMux
    port map (
            O => \N__40925\,
            I => \N__40918\
        );

    \I__8875\ : Span4Mux_h
    port map (
            O => \N__40922\,
            I => \N__40915\
        );

    \I__8874\ : InMux
    port map (
            O => \N__40921\,
            I => \N__40912\
        );

    \I__8873\ : LocalMux
    port map (
            O => \N__40918\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__8872\ : Odrv4
    port map (
            O => \N__40915\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__40912\,
            I => \elapsed_time_ns_1_RNIUVBN9_0_11\
        );

    \I__8870\ : CascadeMux
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__8869\ : InMux
    port map (
            O => \N__40902\,
            I => \N__40899\
        );

    \I__8868\ : LocalMux
    port map (
            O => \N__40899\,
            I => \N__40896\
        );

    \I__8867\ : Odrv4
    port map (
            O => \N__40896\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\
        );

    \I__8866\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40890\
        );

    \I__8865\ : LocalMux
    port map (
            O => \N__40890\,
            I => \N__40887\
        );

    \I__8864\ : Span4Mux_h
    port map (
            O => \N__40887\,
            I => \N__40884\
        );

    \I__8863\ : Odrv4
    port map (
            O => \N__40884\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\
        );

    \I__8862\ : InMux
    port map (
            O => \N__40881\,
            I => \N__40878\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__40878\,
            I => \N__40875\
        );

    \I__8860\ : Span4Mux_h
    port map (
            O => \N__40875\,
            I => \N__40872\
        );

    \I__8859\ : Odrv4
    port map (
            O => \N__40872\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\
        );

    \I__8858\ : InMux
    port map (
            O => \N__40869\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__8857\ : InMux
    port map (
            O => \N__40866\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40863\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__8855\ : InMux
    port map (
            O => \N__40860\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__8854\ : InMux
    port map (
            O => \N__40857\,
            I => \bfn_17_10_0_\
        );

    \I__8853\ : InMux
    port map (
            O => \N__40854\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40851\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__8851\ : InMux
    port map (
            O => \N__40848\,
            I => \N__40841\
        );

    \I__8850\ : InMux
    port map (
            O => \N__40847\,
            I => \N__40841\
        );

    \I__8849\ : InMux
    port map (
            O => \N__40846\,
            I => \N__40838\
        );

    \I__8848\ : LocalMux
    port map (
            O => \N__40841\,
            I => \N__40835\
        );

    \I__8847\ : LocalMux
    port map (
            O => \N__40838\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8846\ : Odrv12
    port map (
            O => \N__40835\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__8845\ : InMux
    port map (
            O => \N__40830\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__8844\ : CascadeMux
    port map (
            O => \N__40827\,
            I => \N__40824\
        );

    \I__8843\ : InMux
    port map (
            O => \N__40824\,
            I => \N__40817\
        );

    \I__8842\ : InMux
    port map (
            O => \N__40823\,
            I => \N__40817\
        );

    \I__8841\ : InMux
    port map (
            O => \N__40822\,
            I => \N__40814\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40817\,
            I => \N__40811\
        );

    \I__8839\ : LocalMux
    port map (
            O => \N__40814\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__8838\ : Odrv12
    port map (
            O => \N__40811\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__8837\ : InMux
    port map (
            O => \N__40806\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__8836\ : InMux
    port map (
            O => \N__40803\,
            I => \N__40799\
        );

    \I__8835\ : InMux
    port map (
            O => \N__40802\,
            I => \N__40796\
        );

    \I__8834\ : LocalMux
    port map (
            O => \N__40799\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__8833\ : LocalMux
    port map (
            O => \N__40796\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__8832\ : InMux
    port map (
            O => \N__40791\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__8831\ : InMux
    port map (
            O => \N__40788\,
            I => \N__40784\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40787\,
            I => \N__40781\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40784\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__8828\ : LocalMux
    port map (
            O => \N__40781\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__8827\ : InMux
    port map (
            O => \N__40776\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__8826\ : InMux
    port map (
            O => \N__40773\,
            I => \N__40769\
        );

    \I__8825\ : InMux
    port map (
            O => \N__40772\,
            I => \N__40766\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__40769\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40766\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__8822\ : InMux
    port map (
            O => \N__40761\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__8821\ : InMux
    port map (
            O => \N__40758\,
            I => \N__40754\
        );

    \I__8820\ : InMux
    port map (
            O => \N__40757\,
            I => \N__40751\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__40754\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8818\ : LocalMux
    port map (
            O => \N__40751\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40746\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40743\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__8815\ : InMux
    port map (
            O => \N__40740\,
            I => \bfn_17_9_0_\
        );

    \I__8814\ : CascadeMux
    port map (
            O => \N__40737\,
            I => \N__40734\
        );

    \I__8813\ : InMux
    port map (
            O => \N__40734\,
            I => \N__40728\
        );

    \I__8812\ : InMux
    port map (
            O => \N__40733\,
            I => \N__40728\
        );

    \I__8811\ : LocalMux
    port map (
            O => \N__40728\,
            I => \N__40724\
        );

    \I__8810\ : InMux
    port map (
            O => \N__40727\,
            I => \N__40721\
        );

    \I__8809\ : Span4Mux_v
    port map (
            O => \N__40724\,
            I => \N__40718\
        );

    \I__8808\ : LocalMux
    port map (
            O => \N__40721\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__8807\ : Odrv4
    port map (
            O => \N__40718\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__8806\ : InMux
    port map (
            O => \N__40713\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__8805\ : InMux
    port map (
            O => \N__40710\,
            I => \N__40704\
        );

    \I__8804\ : InMux
    port map (
            O => \N__40709\,
            I => \N__40704\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__40704\,
            I => \N__40700\
        );

    \I__8802\ : InMux
    port map (
            O => \N__40703\,
            I => \N__40697\
        );

    \I__8801\ : Span4Mux_h
    port map (
            O => \N__40700\,
            I => \N__40694\
        );

    \I__8800\ : LocalMux
    port map (
            O => \N__40697\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8799\ : Odrv4
    port map (
            O => \N__40694\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__8798\ : InMux
    port map (
            O => \N__40689\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__8797\ : InMux
    port map (
            O => \N__40686\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__8796\ : InMux
    port map (
            O => \N__40683\,
            I => \N__40679\
        );

    \I__8795\ : InMux
    port map (
            O => \N__40682\,
            I => \N__40676\
        );

    \I__8794\ : LocalMux
    port map (
            O => \N__40679\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__40676\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40671\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__8791\ : InMux
    port map (
            O => \N__40668\,
            I => \N__40664\
        );

    \I__8790\ : InMux
    port map (
            O => \N__40667\,
            I => \N__40661\
        );

    \I__8789\ : LocalMux
    port map (
            O => \N__40664\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__40661\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__8787\ : InMux
    port map (
            O => \N__40656\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__8786\ : InMux
    port map (
            O => \N__40653\,
            I => \N__40649\
        );

    \I__8785\ : InMux
    port map (
            O => \N__40652\,
            I => \N__40646\
        );

    \I__8784\ : LocalMux
    port map (
            O => \N__40649\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__40646\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__8782\ : InMux
    port map (
            O => \N__40641\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__8781\ : InMux
    port map (
            O => \N__40638\,
            I => \N__40634\
        );

    \I__8780\ : InMux
    port map (
            O => \N__40637\,
            I => \N__40631\
        );

    \I__8779\ : LocalMux
    port map (
            O => \N__40634\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__8778\ : LocalMux
    port map (
            O => \N__40631\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__8777\ : InMux
    port map (
            O => \N__40626\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__8776\ : InMux
    port map (
            O => \N__40623\,
            I => \N__40619\
        );

    \I__8775\ : InMux
    port map (
            O => \N__40622\,
            I => \N__40616\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__40619\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__8773\ : LocalMux
    port map (
            O => \N__40616\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__8772\ : InMux
    port map (
            O => \N__40611\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__8771\ : InMux
    port map (
            O => \N__40608\,
            I => \N__40604\
        );

    \I__8770\ : InMux
    port map (
            O => \N__40607\,
            I => \N__40601\
        );

    \I__8769\ : LocalMux
    port map (
            O => \N__40604\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__40601\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__8767\ : InMux
    port map (
            O => \N__40596\,
            I => \bfn_17_8_0_\
        );

    \I__8766\ : InMux
    port map (
            O => \N__40593\,
            I => \N__40589\
        );

    \I__8765\ : InMux
    port map (
            O => \N__40592\,
            I => \N__40586\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__40589\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8763\ : LocalMux
    port map (
            O => \N__40586\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40581\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__8761\ : InMux
    port map (
            O => \N__40578\,
            I => \N__40574\
        );

    \I__8760\ : InMux
    port map (
            O => \N__40577\,
            I => \N__40571\
        );

    \I__8759\ : LocalMux
    port map (
            O => \N__40574\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__8758\ : LocalMux
    port map (
            O => \N__40571\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__8757\ : InMux
    port map (
            O => \N__40566\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__40563\,
            I => \N__40559\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__40562\,
            I => \N__40556\
        );

    \I__8754\ : InMux
    port map (
            O => \N__40559\,
            I => \N__40553\
        );

    \I__8753\ : InMux
    port map (
            O => \N__40556\,
            I => \N__40549\
        );

    \I__8752\ : LocalMux
    port map (
            O => \N__40553\,
            I => \N__40545\
        );

    \I__8751\ : InMux
    port map (
            O => \N__40552\,
            I => \N__40542\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__40549\,
            I => \N__40539\
        );

    \I__8749\ : InMux
    port map (
            O => \N__40548\,
            I => \N__40536\
        );

    \I__8748\ : Span4Mux_v
    port map (
            O => \N__40545\,
            I => \N__40533\
        );

    \I__8747\ : LocalMux
    port map (
            O => \N__40542\,
            I => \N__40530\
        );

    \I__8746\ : Span4Mux_h
    port map (
            O => \N__40539\,
            I => \N__40525\
        );

    \I__8745\ : LocalMux
    port map (
            O => \N__40536\,
            I => \N__40525\
        );

    \I__8744\ : Odrv4
    port map (
            O => \N__40533\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8743\ : Odrv4
    port map (
            O => \N__40530\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8742\ : Odrv4
    port map (
            O => \N__40525\,
            I => \current_shift_inst.elapsed_time_ns_s1_18\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__40518\,
            I => \N__40515\
        );

    \I__8740\ : InMux
    port map (
            O => \N__40515\,
            I => \N__40512\
        );

    \I__8739\ : LocalMux
    port map (
            O => \N__40512\,
            I => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\
        );

    \I__8738\ : CascadeMux
    port map (
            O => \N__40509\,
            I => \N__40506\
        );

    \I__8737\ : InMux
    port map (
            O => \N__40506\,
            I => \N__40503\
        );

    \I__8736\ : LocalMux
    port map (
            O => \N__40503\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\
        );

    \I__8735\ : InMux
    port map (
            O => \N__40500\,
            I => \N__40497\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40497\,
            I => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\
        );

    \I__8733\ : CascadeMux
    port map (
            O => \N__40494\,
            I => \N__40491\
        );

    \I__8732\ : InMux
    port map (
            O => \N__40491\,
            I => \N__40488\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__40488\,
            I => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\
        );

    \I__8730\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40482\
        );

    \I__8729\ : LocalMux
    port map (
            O => \N__40482\,
            I => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\
        );

    \I__8728\ : InMux
    port map (
            O => \N__40479\,
            I => \N__40474\
        );

    \I__8727\ : InMux
    port map (
            O => \N__40478\,
            I => \N__40469\
        );

    \I__8726\ : InMux
    port map (
            O => \N__40477\,
            I => \N__40469\
        );

    \I__8725\ : LocalMux
    port map (
            O => \N__40474\,
            I => \N__40465\
        );

    \I__8724\ : LocalMux
    port map (
            O => \N__40469\,
            I => \N__40462\
        );

    \I__8723\ : InMux
    port map (
            O => \N__40468\,
            I => \N__40459\
        );

    \I__8722\ : Span4Mux_h
    port map (
            O => \N__40465\,
            I => \N__40454\
        );

    \I__8721\ : Span4Mux_h
    port map (
            O => \N__40462\,
            I => \N__40454\
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__40459\,
            I => \N__40451\
        );

    \I__8719\ : Span4Mux_v
    port map (
            O => \N__40454\,
            I => \N__40448\
        );

    \I__8718\ : Span4Mux_h
    port map (
            O => \N__40451\,
            I => \N__40445\
        );

    \I__8717\ : Odrv4
    port map (
            O => \N__40448\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8716\ : Odrv4
    port map (
            O => \N__40445\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\
        );

    \I__8715\ : InMux
    port map (
            O => \N__40440\,
            I => \N__40437\
        );

    \I__8714\ : LocalMux
    port map (
            O => \N__40437\,
            I => \N__40433\
        );

    \I__8713\ : InMux
    port map (
            O => \N__40436\,
            I => \N__40430\
        );

    \I__8712\ : Odrv12
    port map (
            O => \N__40433\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__40430\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24\
        );

    \I__8710\ : InMux
    port map (
            O => \N__40425\,
            I => \N__40422\
        );

    \I__8709\ : LocalMux
    port map (
            O => \N__40422\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\
        );

    \I__8708\ : CascadeMux
    port map (
            O => \N__40419\,
            I => \N__40415\
        );

    \I__8707\ : InMux
    port map (
            O => \N__40418\,
            I => \N__40411\
        );

    \I__8706\ : InMux
    port map (
            O => \N__40415\,
            I => \N__40408\
        );

    \I__8705\ : InMux
    port map (
            O => \N__40414\,
            I => \N__40405\
        );

    \I__8704\ : LocalMux
    port map (
            O => \N__40411\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8703\ : LocalMux
    port map (
            O => \N__40408\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8702\ : LocalMux
    port map (
            O => \N__40405\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__8701\ : InMux
    port map (
            O => \N__40398\,
            I => \N__40394\
        );

    \I__8700\ : InMux
    port map (
            O => \N__40397\,
            I => \N__40391\
        );

    \I__8699\ : LocalMux
    port map (
            O => \N__40394\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__8698\ : LocalMux
    port map (
            O => \N__40391\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__8697\ : InMux
    port map (
            O => \N__40386\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__8696\ : CascadeMux
    port map (
            O => \N__40383\,
            I => \N__40380\
        );

    \I__8695\ : InMux
    port map (
            O => \N__40380\,
            I => \N__40377\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__40377\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\
        );

    \I__8693\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40370\
        );

    \I__8692\ : InMux
    port map (
            O => \N__40373\,
            I => \N__40367\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__40370\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__40367\,
            I => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__8689\ : InMux
    port map (
            O => \N__40362\,
            I => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__8688\ : InMux
    port map (
            O => \N__40359\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\
        );

    \I__8687\ : InMux
    port map (
            O => \N__40356\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\
        );

    \I__8686\ : InMux
    port map (
            O => \N__40353\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\
        );

    \I__8685\ : InMux
    port map (
            O => \N__40350\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\
        );

    \I__8684\ : CascadeMux
    port map (
            O => \N__40347\,
            I => \N__40344\
        );

    \I__8683\ : InMux
    port map (
            O => \N__40344\,
            I => \N__40341\
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__40341\,
            I => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40338\,
            I => \N__40335\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__40335\,
            I => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\
        );

    \I__8679\ : InMux
    port map (
            O => \N__40332\,
            I => \N__40329\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40329\,
            I => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\
        );

    \I__8677\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40321\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40325\,
            I => \N__40318\
        );

    \I__8675\ : InMux
    port map (
            O => \N__40324\,
            I => \N__40314\
        );

    \I__8674\ : LocalMux
    port map (
            O => \N__40321\,
            I => \N__40309\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__40318\,
            I => \N__40309\
        );

    \I__8672\ : InMux
    port map (
            O => \N__40317\,
            I => \N__40306\
        );

    \I__8671\ : LocalMux
    port map (
            O => \N__40314\,
            I => \N__40303\
        );

    \I__8670\ : Span4Mux_h
    port map (
            O => \N__40309\,
            I => \N__40298\
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__40306\,
            I => \N__40298\
        );

    \I__8668\ : Odrv12
    port map (
            O => \N__40303\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__40298\,
            I => \current_shift_inst.elapsed_time_ns_s1_22\
        );

    \I__8666\ : CascadeMux
    port map (
            O => \N__40293\,
            I => \N__40290\
        );

    \I__8665\ : InMux
    port map (
            O => \N__40290\,
            I => \N__40287\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__40287\,
            I => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\
        );

    \I__8663\ : CascadeMux
    port map (
            O => \N__40284\,
            I => \N__40281\
        );

    \I__8662\ : InMux
    port map (
            O => \N__40281\,
            I => \N__40278\
        );

    \I__8661\ : LocalMux
    port map (
            O => \N__40278\,
            I => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\
        );

    \I__8660\ : InMux
    port map (
            O => \N__40275\,
            I => \bfn_16_21_0_\
        );

    \I__8659\ : InMux
    port map (
            O => \N__40272\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\
        );

    \I__8658\ : InMux
    port map (
            O => \N__40269\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\
        );

    \I__8657\ : InMux
    port map (
            O => \N__40266\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\
        );

    \I__8656\ : CascadeMux
    port map (
            O => \N__40263\,
            I => \N__40260\
        );

    \I__8655\ : InMux
    port map (
            O => \N__40260\,
            I => \N__40257\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40257\,
            I => \N__40253\
        );

    \I__8653\ : InMux
    port map (
            O => \N__40256\,
            I => \N__40250\
        );

    \I__8652\ : Sp12to4
    port map (
            O => \N__40253\,
            I => \N__40245\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__40250\,
            I => \N__40242\
        );

    \I__8650\ : InMux
    port map (
            O => \N__40249\,
            I => \N__40237\
        );

    \I__8649\ : InMux
    port map (
            O => \N__40248\,
            I => \N__40237\
        );

    \I__8648\ : Span12Mux_v
    port map (
            O => \N__40245\,
            I => \N__40234\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__40242\,
            I => \N__40229\
        );

    \I__8646\ : LocalMux
    port map (
            O => \N__40237\,
            I => \N__40229\
        );

    \I__8645\ : Odrv12
    port map (
            O => \N__40234\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8644\ : Odrv4
    port map (
            O => \N__40229\,
            I => \current_shift_inst.elapsed_time_ns_s1_23\
        );

    \I__8643\ : InMux
    port map (
            O => \N__40224\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\
        );

    \I__8642\ : InMux
    port map (
            O => \N__40221\,
            I => \N__40217\
        );

    \I__8641\ : InMux
    port map (
            O => \N__40220\,
            I => \N__40214\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__40217\,
            I => \N__40210\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__40214\,
            I => \N__40207\
        );

    \I__8638\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40204\
        );

    \I__8637\ : Span4Mux_v
    port map (
            O => \N__40210\,
            I => \N__40200\
        );

    \I__8636\ : Span4Mux_h
    port map (
            O => \N__40207\,
            I => \N__40197\
        );

    \I__8635\ : LocalMux
    port map (
            O => \N__40204\,
            I => \N__40194\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40191\
        );

    \I__8633\ : Odrv4
    port map (
            O => \N__40200\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8632\ : Odrv4
    port map (
            O => \N__40197\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8631\ : Odrv4
    port map (
            O => \N__40194\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8630\ : LocalMux
    port map (
            O => \N__40191\,
            I => \current_shift_inst.elapsed_time_ns_s1_24\
        );

    \I__8629\ : InMux
    port map (
            O => \N__40182\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\
        );

    \I__8628\ : InMux
    port map (
            O => \N__40179\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40176\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\
        );

    \I__8626\ : InMux
    port map (
            O => \N__40173\,
            I => \bfn_16_22_0_\
        );

    \I__8625\ : CascadeMux
    port map (
            O => \N__40170\,
            I => \N__40167\
        );

    \I__8624\ : InMux
    port map (
            O => \N__40167\,
            I => \N__40163\
        );

    \I__8623\ : CascadeMux
    port map (
            O => \N__40166\,
            I => \N__40160\
        );

    \I__8622\ : LocalMux
    port map (
            O => \N__40163\,
            I => \N__40155\
        );

    \I__8621\ : InMux
    port map (
            O => \N__40160\,
            I => \N__40152\
        );

    \I__8620\ : InMux
    port map (
            O => \N__40159\,
            I => \N__40147\
        );

    \I__8619\ : InMux
    port map (
            O => \N__40158\,
            I => \N__40147\
        );

    \I__8618\ : Sp12to4
    port map (
            O => \N__40155\,
            I => \N__40142\
        );

    \I__8617\ : LocalMux
    port map (
            O => \N__40152\,
            I => \N__40142\
        );

    \I__8616\ : LocalMux
    port map (
            O => \N__40147\,
            I => \N__40139\
        );

    \I__8615\ : Odrv12
    port map (
            O => \N__40142\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8614\ : Odrv4
    port map (
            O => \N__40139\,
            I => \current_shift_inst.elapsed_time_ns_s1_10\
        );

    \I__8613\ : InMux
    port map (
            O => \N__40134\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\
        );

    \I__8612\ : InMux
    port map (
            O => \N__40131\,
            I => \bfn_16_20_0_\
        );

    \I__8611\ : InMux
    port map (
            O => \N__40128\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\
        );

    \I__8610\ : InMux
    port map (
            O => \N__40125\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\
        );

    \I__8609\ : InMux
    port map (
            O => \N__40122\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\
        );

    \I__8608\ : InMux
    port map (
            O => \N__40119\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\
        );

    \I__8607\ : InMux
    port map (
            O => \N__40116\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\
        );

    \I__8606\ : InMux
    port map (
            O => \N__40113\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\
        );

    \I__8605\ : InMux
    port map (
            O => \N__40110\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\
        );

    \I__8604\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40104\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__40104\,
            I => \N__40101\
        );

    \I__8602\ : Span4Mux_v
    port map (
            O => \N__40101\,
            I => \N__40098\
        );

    \I__8601\ : Odrv4
    port map (
            O => \N__40098\,
            I => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\
        );

    \I__8600\ : CascadeMux
    port map (
            O => \N__40095\,
            I => \N__40091\
        );

    \I__8599\ : CascadeMux
    port map (
            O => \N__40094\,
            I => \N__40088\
        );

    \I__8598\ : InMux
    port map (
            O => \N__40091\,
            I => \N__40085\
        );

    \I__8597\ : InMux
    port map (
            O => \N__40088\,
            I => \N__40082\
        );

    \I__8596\ : LocalMux
    port map (
            O => \N__40085\,
            I => \N__40075\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__40082\,
            I => \N__40075\
        );

    \I__8594\ : InMux
    port map (
            O => \N__40081\,
            I => \N__40072\
        );

    \I__8593\ : InMux
    port map (
            O => \N__40080\,
            I => \N__40069\
        );

    \I__8592\ : Span4Mux_v
    port map (
            O => \N__40075\,
            I => \N__40066\
        );

    \I__8591\ : LocalMux
    port map (
            O => \N__40072\,
            I => \N__40063\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__40069\,
            I => \N__40060\
        );

    \I__8589\ : Odrv4
    port map (
            O => \N__40066\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8588\ : Odrv12
    port map (
            O => \N__40063\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__40060\,
            I => \current_shift_inst.elapsed_time_ns_s1_3\
        );

    \I__8586\ : InMux
    port map (
            O => \N__40053\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\
        );

    \I__8585\ : InMux
    port map (
            O => \N__40050\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40047\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\
        );

    \I__8583\ : InMux
    port map (
            O => \N__40044\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\
        );

    \I__8582\ : CascadeMux
    port map (
            O => \N__40041\,
            I => \N__40038\
        );

    \I__8581\ : InMux
    port map (
            O => \N__40038\,
            I => \N__40034\
        );

    \I__8580\ : CascadeMux
    port map (
            O => \N__40037\,
            I => \N__40031\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__40034\,
            I => \N__40028\
        );

    \I__8578\ : InMux
    port map (
            O => \N__40031\,
            I => \N__40024\
        );

    \I__8577\ : Span4Mux_h
    port map (
            O => \N__40028\,
            I => \N__40021\
        );

    \I__8576\ : InMux
    port map (
            O => \N__40027\,
            I => \N__40018\
        );

    \I__8575\ : LocalMux
    port map (
            O => \N__40024\,
            I => \N__40015\
        );

    \I__8574\ : Span4Mux_v
    port map (
            O => \N__40021\,
            I => \N__40012\
        );

    \I__8573\ : LocalMux
    port map (
            O => \N__40018\,
            I => \N__40009\
        );

    \I__8572\ : Span4Mux_v
    port map (
            O => \N__40015\,
            I => \N__40005\
        );

    \I__8571\ : Span4Mux_h
    port map (
            O => \N__40012\,
            I => \N__40002\
        );

    \I__8570\ : Span4Mux_v
    port map (
            O => \N__40009\,
            I => \N__39999\
        );

    \I__8569\ : InMux
    port map (
            O => \N__40008\,
            I => \N__39996\
        );

    \I__8568\ : Odrv4
    port map (
            O => \N__40005\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8567\ : Odrv4
    port map (
            O => \N__40002\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8566\ : Odrv4
    port map (
            O => \N__39999\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__39996\,
            I => \current_shift_inst.elapsed_time_ns_s1_8\
        );

    \I__8564\ : InMux
    port map (
            O => \N__39987\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\
        );

    \I__8563\ : InMux
    port map (
            O => \N__39984\,
            I => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__39981\,
            I => \N__39978\
        );

    \I__8561\ : InMux
    port map (
            O => \N__39978\,
            I => \N__39975\
        );

    \I__8560\ : LocalMux
    port map (
            O => \N__39975\,
            I => \N__39972\
        );

    \I__8559\ : Span4Mux_v
    port map (
            O => \N__39972\,
            I => \N__39969\
        );

    \I__8558\ : Odrv4
    port map (
            O => \N__39969\,
            I => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\
        );

    \I__8557\ : CascadeMux
    port map (
            O => \N__39966\,
            I => \N__39963\
        );

    \I__8556\ : InMux
    port map (
            O => \N__39963\,
            I => \N__39960\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39960\,
            I => \N__39957\
        );

    \I__8554\ : Odrv12
    port map (
            O => \N__39957\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\
        );

    \I__8553\ : CascadeMux
    port map (
            O => \N__39954\,
            I => \N__39951\
        );

    \I__8552\ : InMux
    port map (
            O => \N__39951\,
            I => \N__39948\
        );

    \I__8551\ : LocalMux
    port map (
            O => \N__39948\,
            I => \N__39945\
        );

    \I__8550\ : Span4Mux_v
    port map (
            O => \N__39945\,
            I => \N__39942\
        );

    \I__8549\ : Odrv4
    port map (
            O => \N__39942\,
            I => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\
        );

    \I__8548\ : CascadeMux
    port map (
            O => \N__39939\,
            I => \N__39936\
        );

    \I__8547\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39933\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__39933\,
            I => \N__39930\
        );

    \I__8545\ : Span4Mux_h
    port map (
            O => \N__39930\,
            I => \N__39927\
        );

    \I__8544\ : Odrv4
    port map (
            O => \N__39927\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\
        );

    \I__8543\ : CascadeMux
    port map (
            O => \N__39924\,
            I => \N__39921\
        );

    \I__8542\ : InMux
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__8541\ : LocalMux
    port map (
            O => \N__39918\,
            I => \N__39915\
        );

    \I__8540\ : Span4Mux_v
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__8539\ : Odrv4
    port map (
            O => \N__39912\,
            I => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\
        );

    \I__8538\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39906\
        );

    \I__8537\ : LocalMux
    port map (
            O => \N__39906\,
            I => \N__39903\
        );

    \I__8536\ : Span4Mux_v
    port map (
            O => \N__39903\,
            I => \N__39900\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__39900\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\
        );

    \I__8534\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39894\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39891\
        );

    \I__8532\ : Odrv4
    port map (
            O => \N__39891\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\
        );

    \I__8531\ : CascadeMux
    port map (
            O => \N__39888\,
            I => \N__39885\
        );

    \I__8530\ : InMux
    port map (
            O => \N__39885\,
            I => \N__39882\
        );

    \I__8529\ : LocalMux
    port map (
            O => \N__39882\,
            I => \N__39879\
        );

    \I__8528\ : Span4Mux_v
    port map (
            O => \N__39879\,
            I => \N__39876\
        );

    \I__8527\ : Span4Mux_v
    port map (
            O => \N__39876\,
            I => \N__39873\
        );

    \I__8526\ : Odrv4
    port map (
            O => \N__39873\,
            I => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\
        );

    \I__8525\ : InMux
    port map (
            O => \N__39870\,
            I => \N__39867\
        );

    \I__8524\ : LocalMux
    port map (
            O => \N__39867\,
            I => \N__39864\
        );

    \I__8523\ : Span4Mux_v
    port map (
            O => \N__39864\,
            I => \N__39861\
        );

    \I__8522\ : Odrv4
    port map (
            O => \N__39861\,
            I => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\
        );

    \I__8521\ : InMux
    port map (
            O => \N__39858\,
            I => \N__39855\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__39855\,
            I => \N__39852\
        );

    \I__8519\ : Span4Mux_v
    port map (
            O => \N__39852\,
            I => \N__39849\
        );

    \I__8518\ : Span4Mux_v
    port map (
            O => \N__39849\,
            I => \N__39846\
        );

    \I__8517\ : Odrv4
    port map (
            O => \N__39846\,
            I => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\
        );

    \I__8516\ : CascadeMux
    port map (
            O => \N__39843\,
            I => \N__39840\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39840\,
            I => \N__39837\
        );

    \I__8514\ : LocalMux
    port map (
            O => \N__39837\,
            I => \N__39834\
        );

    \I__8513\ : Span4Mux_v
    port map (
            O => \N__39834\,
            I => \N__39831\
        );

    \I__8512\ : Odrv4
    port map (
            O => \N__39831\,
            I => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\
        );

    \I__8511\ : InMux
    port map (
            O => \N__39828\,
            I => \N__39825\
        );

    \I__8510\ : LocalMux
    port map (
            O => \N__39825\,
            I => \N__39822\
        );

    \I__8509\ : Span4Mux_v
    port map (
            O => \N__39822\,
            I => \N__39819\
        );

    \I__8508\ : Odrv4
    port map (
            O => \N__39819\,
            I => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\
        );

    \I__8507\ : CascadeMux
    port map (
            O => \N__39816\,
            I => \N__39813\
        );

    \I__8506\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39810\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__39810\,
            I => \N__39807\
        );

    \I__8504\ : Span4Mux_v
    port map (
            O => \N__39807\,
            I => \N__39804\
        );

    \I__8503\ : Odrv4
    port map (
            O => \N__39804\,
            I => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\
        );

    \I__8502\ : InMux
    port map (
            O => \N__39801\,
            I => \N__39798\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__39798\,
            I => \N__39795\
        );

    \I__8500\ : Span4Mux_v
    port map (
            O => \N__39795\,
            I => \N__39792\
        );

    \I__8499\ : Odrv4
    port map (
            O => \N__39792\,
            I => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\
        );

    \I__8498\ : InMux
    port map (
            O => \N__39789\,
            I => \N__39786\
        );

    \I__8497\ : LocalMux
    port map (
            O => \N__39786\,
            I => \N__39783\
        );

    \I__8496\ : Span4Mux_h
    port map (
            O => \N__39783\,
            I => \N__39780\
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__39780\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\
        );

    \I__8494\ : CascadeMux
    port map (
            O => \N__39777\,
            I => \N__39774\
        );

    \I__8493\ : InMux
    port map (
            O => \N__39774\,
            I => \N__39771\
        );

    \I__8492\ : LocalMux
    port map (
            O => \N__39771\,
            I => \N__39768\
        );

    \I__8491\ : Span4Mux_v
    port map (
            O => \N__39768\,
            I => \N__39765\
        );

    \I__8490\ : Odrv4
    port map (
            O => \N__39765\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\
        );

    \I__8489\ : InMux
    port map (
            O => \N__39762\,
            I => \N__39759\
        );

    \I__8488\ : LocalMux
    port map (
            O => \N__39759\,
            I => \N__39756\
        );

    \I__8487\ : Span4Mux_v
    port map (
            O => \N__39756\,
            I => \N__39753\
        );

    \I__8486\ : Odrv4
    port map (
            O => \N__39753\,
            I => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\
        );

    \I__8485\ : InMux
    port map (
            O => \N__39750\,
            I => \N__39747\
        );

    \I__8484\ : LocalMux
    port map (
            O => \N__39747\,
            I => \N__39744\
        );

    \I__8483\ : Span4Mux_h
    port map (
            O => \N__39744\,
            I => \N__39741\
        );

    \I__8482\ : Odrv4
    port map (
            O => \N__39741\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39738\,
            I => \N__39735\
        );

    \I__8480\ : LocalMux
    port map (
            O => \N__39735\,
            I => \N__39732\
        );

    \I__8479\ : Span4Mux_v
    port map (
            O => \N__39732\,
            I => \N__39729\
        );

    \I__8478\ : Odrv4
    port map (
            O => \N__39729\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\
        );

    \I__8477\ : InMux
    port map (
            O => \N__39726\,
            I => \N__39723\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__39723\,
            I => \N__39720\
        );

    \I__8475\ : Span4Mux_v
    port map (
            O => \N__39720\,
            I => \N__39717\
        );

    \I__8474\ : Span4Mux_v
    port map (
            O => \N__39717\,
            I => \N__39714\
        );

    \I__8473\ : Odrv4
    port map (
            O => \N__39714\,
            I => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__39711\,
            I => \N__39708\
        );

    \I__8471\ : InMux
    port map (
            O => \N__39708\,
            I => \N__39705\
        );

    \I__8470\ : LocalMux
    port map (
            O => \N__39705\,
            I => \N__39702\
        );

    \I__8469\ : Span4Mux_v
    port map (
            O => \N__39702\,
            I => \N__39699\
        );

    \I__8468\ : Odrv4
    port map (
            O => \N__39699\,
            I => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\
        );

    \I__8467\ : InMux
    port map (
            O => \N__39696\,
            I => \N__39690\
        );

    \I__8466\ : InMux
    port map (
            O => \N__39695\,
            I => \N__39685\
        );

    \I__8465\ : InMux
    port map (
            O => \N__39694\,
            I => \N__39685\
        );

    \I__8464\ : InMux
    port map (
            O => \N__39693\,
            I => \N__39682\
        );

    \I__8463\ : LocalMux
    port map (
            O => \N__39690\,
            I => \N__39679\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__39685\,
            I => \N__39676\
        );

    \I__8461\ : LocalMux
    port map (
            O => \N__39682\,
            I => \N__39673\
        );

    \I__8460\ : Span4Mux_h
    port map (
            O => \N__39679\,
            I => \N__39670\
        );

    \I__8459\ : Span4Mux_v
    port map (
            O => \N__39676\,
            I => \N__39667\
        );

    \I__8458\ : Span4Mux_v
    port map (
            O => \N__39673\,
            I => \N__39664\
        );

    \I__8457\ : Odrv4
    port map (
            O => \N__39670\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__8456\ : Odrv4
    port map (
            O => \N__39667\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__8455\ : Odrv4
    port map (
            O => \N__39664\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\
        );

    \I__8454\ : InMux
    port map (
            O => \N__39657\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__8453\ : InMux
    port map (
            O => \N__39654\,
            I => \N__39650\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39645\
        );

    \I__8451\ : LocalMux
    port map (
            O => \N__39650\,
            I => \N__39642\
        );

    \I__8450\ : InMux
    port map (
            O => \N__39649\,
            I => \N__39639\
        );

    \I__8449\ : InMux
    port map (
            O => \N__39648\,
            I => \N__39636\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__39645\,
            I => \N__39633\
        );

    \I__8447\ : Span4Mux_v
    port map (
            O => \N__39642\,
            I => \N__39626\
        );

    \I__8446\ : LocalMux
    port map (
            O => \N__39639\,
            I => \N__39626\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__39636\,
            I => \N__39626\
        );

    \I__8444\ : Span4Mux_v
    port map (
            O => \N__39633\,
            I => \N__39623\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__39626\,
            I => \N__39620\
        );

    \I__8442\ : Odrv4
    port map (
            O => \N__39623\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__8441\ : Odrv4
    port map (
            O => \N__39620\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\
        );

    \I__8440\ : InMux
    port map (
            O => \N__39615\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__8439\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39607\
        );

    \I__8438\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39604\
        );

    \I__8437\ : CascadeMux
    port map (
            O => \N__39610\,
            I => \N__39601\
        );

    \I__8436\ : LocalMux
    port map (
            O => \N__39607\,
            I => \N__39595\
        );

    \I__8435\ : LocalMux
    port map (
            O => \N__39604\,
            I => \N__39595\
        );

    \I__8434\ : InMux
    port map (
            O => \N__39601\,
            I => \N__39592\
        );

    \I__8433\ : InMux
    port map (
            O => \N__39600\,
            I => \N__39589\
        );

    \I__8432\ : Span4Mux_v
    port map (
            O => \N__39595\,
            I => \N__39584\
        );

    \I__8431\ : LocalMux
    port map (
            O => \N__39592\,
            I => \N__39584\
        );

    \I__8430\ : LocalMux
    port map (
            O => \N__39589\,
            I => \N__39581\
        );

    \I__8429\ : Span4Mux_h
    port map (
            O => \N__39584\,
            I => \N__39578\
        );

    \I__8428\ : Odrv12
    port map (
            O => \N__39581\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8427\ : Odrv4
    port map (
            O => \N__39578\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\
        );

    \I__8426\ : InMux
    port map (
            O => \N__39573\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__8425\ : InMux
    port map (
            O => \N__39570\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__8424\ : InMux
    port map (
            O => \N__39567\,
            I => \N__39564\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__39564\,
            I => \N__39558\
        );

    \I__8422\ : InMux
    port map (
            O => \N__39563\,
            I => \N__39555\
        );

    \I__8421\ : InMux
    port map (
            O => \N__39562\,
            I => \N__39550\
        );

    \I__8420\ : InMux
    port map (
            O => \N__39561\,
            I => \N__39550\
        );

    \I__8419\ : Span4Mux_v
    port map (
            O => \N__39558\,
            I => \N__39543\
        );

    \I__8418\ : LocalMux
    port map (
            O => \N__39555\,
            I => \N__39543\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__39550\,
            I => \N__39543\
        );

    \I__8416\ : Span4Mux_h
    port map (
            O => \N__39543\,
            I => \N__39540\
        );

    \I__8415\ : Odrv4
    port map (
            O => \N__39540\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\
        );

    \I__8414\ : CascadeMux
    port map (
            O => \N__39537\,
            I => \N__39534\
        );

    \I__8413\ : InMux
    port map (
            O => \N__39534\,
            I => \N__39529\
        );

    \I__8412\ : InMux
    port map (
            O => \N__39533\,
            I => \N__39526\
        );

    \I__8411\ : CascadeMux
    port map (
            O => \N__39532\,
            I => \N__39522\
        );

    \I__8410\ : LocalMux
    port map (
            O => \N__39529\,
            I => \N__39517\
        );

    \I__8409\ : LocalMux
    port map (
            O => \N__39526\,
            I => \N__39517\
        );

    \I__8408\ : InMux
    port map (
            O => \N__39525\,
            I => \N__39512\
        );

    \I__8407\ : InMux
    port map (
            O => \N__39522\,
            I => \N__39512\
        );

    \I__8406\ : Span4Mux_v
    port map (
            O => \N__39517\,
            I => \N__39507\
        );

    \I__8405\ : LocalMux
    port map (
            O => \N__39512\,
            I => \N__39507\
        );

    \I__8404\ : Odrv4
    port map (
            O => \N__39507\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\
        );

    \I__8403\ : InMux
    port map (
            O => \N__39504\,
            I => \N__39501\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__39501\,
            I => \N__39498\
        );

    \I__8401\ : Span4Mux_h
    port map (
            O => \N__39498\,
            I => \N__39495\
        );

    \I__8400\ : Odrv4
    port map (
            O => \N__39495\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\
        );

    \I__8399\ : CascadeMux
    port map (
            O => \N__39492\,
            I => \N__39489\
        );

    \I__8398\ : InMux
    port map (
            O => \N__39489\,
            I => \N__39486\
        );

    \I__8397\ : LocalMux
    port map (
            O => \N__39486\,
            I => \N__39483\
        );

    \I__8396\ : Span4Mux_v
    port map (
            O => \N__39483\,
            I => \N__39480\
        );

    \I__8395\ : Odrv4
    port map (
            O => \N__39480\,
            I => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\
        );

    \I__8394\ : InMux
    port map (
            O => \N__39477\,
            I => \N__39474\
        );

    \I__8393\ : LocalMux
    port map (
            O => \N__39474\,
            I => \N__39471\
        );

    \I__8392\ : Span4Mux_v
    port map (
            O => \N__39471\,
            I => \N__39468\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__39468\,
            I => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\
        );

    \I__8390\ : InMux
    port map (
            O => \N__39465\,
            I => \N__39461\
        );

    \I__8389\ : InMux
    port map (
            O => \N__39464\,
            I => \N__39457\
        );

    \I__8388\ : LocalMux
    port map (
            O => \N__39461\,
            I => \N__39454\
        );

    \I__8387\ : InMux
    port map (
            O => \N__39460\,
            I => \N__39451\
        );

    \I__8386\ : LocalMux
    port map (
            O => \N__39457\,
            I => \N__39447\
        );

    \I__8385\ : Span4Mux_h
    port map (
            O => \N__39454\,
            I => \N__39442\
        );

    \I__8384\ : LocalMux
    port map (
            O => \N__39451\,
            I => \N__39442\
        );

    \I__8383\ : InMux
    port map (
            O => \N__39450\,
            I => \N__39439\
        );

    \I__8382\ : Span4Mux_v
    port map (
            O => \N__39447\,
            I => \N__39436\
        );

    \I__8381\ : Odrv4
    port map (
            O => \N__39442\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__39439\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__8379\ : Odrv4
    port map (
            O => \N__39436\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\
        );

    \I__8378\ : InMux
    port map (
            O => \N__39429\,
            I => \bfn_16_12_0_\
        );

    \I__8377\ : InMux
    port map (
            O => \N__39426\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__8376\ : InMux
    port map (
            O => \N__39423\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__8375\ : InMux
    port map (
            O => \N__39420\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__8374\ : InMux
    port map (
            O => \N__39417\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__8373\ : InMux
    port map (
            O => \N__39414\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__8372\ : InMux
    port map (
            O => \N__39411\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__8371\ : InMux
    port map (
            O => \N__39408\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__8370\ : InMux
    port map (
            O => \N__39405\,
            I => \bfn_16_13_0_\
        );

    \I__8369\ : InMux
    port map (
            O => \N__39402\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__8368\ : InMux
    port map (
            O => \N__39399\,
            I => \bfn_16_11_0_\
        );

    \I__8367\ : InMux
    port map (
            O => \N__39396\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__8366\ : InMux
    port map (
            O => \N__39393\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__8365\ : InMux
    port map (
            O => \N__39390\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__8364\ : InMux
    port map (
            O => \N__39387\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__8363\ : InMux
    port map (
            O => \N__39384\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__8362\ : InMux
    port map (
            O => \N__39381\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__8361\ : InMux
    port map (
            O => \N__39378\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__8360\ : InMux
    port map (
            O => \N__39375\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30\
        );

    \I__8359\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39365\
        );

    \I__8358\ : InMux
    port map (
            O => \N__39371\,
            I => \N__39365\
        );

    \I__8357\ : InMux
    port map (
            O => \N__39370\,
            I => \N__39362\
        );

    \I__8356\ : LocalMux
    port map (
            O => \N__39365\,
            I => \N__39357\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__39362\,
            I => \N__39357\
        );

    \I__8354\ : Odrv12
    port map (
            O => \N__39357\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__8353\ : InMux
    port map (
            O => \N__39354\,
            I => \N__39349\
        );

    \I__8352\ : InMux
    port map (
            O => \N__39353\,
            I => \N__39346\
        );

    \I__8351\ : InMux
    port map (
            O => \N__39352\,
            I => \N__39343\
        );

    \I__8350\ : LocalMux
    port map (
            O => \N__39349\,
            I => \N__39338\
        );

    \I__8349\ : LocalMux
    port map (
            O => \N__39346\,
            I => \N__39338\
        );

    \I__8348\ : LocalMux
    port map (
            O => \N__39343\,
            I => \N__39334\
        );

    \I__8347\ : Span4Mux_v
    port map (
            O => \N__39338\,
            I => \N__39331\
        );

    \I__8346\ : InMux
    port map (
            O => \N__39337\,
            I => \N__39328\
        );

    \I__8345\ : Odrv4
    port map (
            O => \N__39334\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8344\ : Odrv4
    port map (
            O => \N__39331\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8343\ : LocalMux
    port map (
            O => \N__39328\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\
        );

    \I__8342\ : InMux
    port map (
            O => \N__39321\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__8341\ : InMux
    port map (
            O => \N__39318\,
            I => \N__39310\
        );

    \I__8340\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39310\
        );

    \I__8339\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39307\
        );

    \I__8338\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39304\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__39310\,
            I => \N__39301\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__39307\,
            I => \N__39298\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__39304\,
            I => \N__39295\
        );

    \I__8334\ : Span4Mux_h
    port map (
            O => \N__39301\,
            I => \N__39292\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__39298\,
            I => \N__39289\
        );

    \I__8332\ : Odrv4
    port map (
            O => \N__39295\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8331\ : Odrv4
    port map (
            O => \N__39292\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8330\ : Odrv4
    port map (
            O => \N__39289\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39282\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__8328\ : InMux
    port map (
            O => \N__39279\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39276\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__8326\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39269\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39272\,
            I => \N__39265\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__39269\,
            I => \N__39261\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39268\,
            I => \N__39258\
        );

    \I__8322\ : LocalMux
    port map (
            O => \N__39265\,
            I => \N__39255\
        );

    \I__8321\ : InMux
    port map (
            O => \N__39264\,
            I => \N__39252\
        );

    \I__8320\ : Span4Mux_v
    port map (
            O => \N__39261\,
            I => \N__39247\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39258\,
            I => \N__39247\
        );

    \I__8318\ : Span4Mux_h
    port map (
            O => \N__39255\,
            I => \N__39240\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39252\,
            I => \N__39240\
        );

    \I__8316\ : Span4Mux_h
    port map (
            O => \N__39247\,
            I => \N__39240\
        );

    \I__8315\ : Span4Mux_v
    port map (
            O => \N__39240\,
            I => \N__39237\
        );

    \I__8314\ : Odrv4
    port map (
            O => \N__39237\,
            I => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\
        );

    \I__8313\ : InMux
    port map (
            O => \N__39234\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__8312\ : InMux
    port map (
            O => \N__39231\,
            I => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__8311\ : InMux
    port map (
            O => \N__39228\,
            I => \N__39225\
        );

    \I__8310\ : LocalMux
    port map (
            O => \N__39225\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\
        );

    \I__8309\ : InMux
    port map (
            O => \N__39222\,
            I => \N__39219\
        );

    \I__8308\ : LocalMux
    port map (
            O => \N__39219\,
            I => \N__39216\
        );

    \I__8307\ : Span4Mux_v
    port map (
            O => \N__39216\,
            I => \N__39213\
        );

    \I__8306\ : Odrv4
    port map (
            O => \N__39213\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\
        );

    \I__8305\ : CascadeMux
    port map (
            O => \N__39210\,
            I => \N__39207\
        );

    \I__8304\ : InMux
    port map (
            O => \N__39207\,
            I => \N__39204\
        );

    \I__8303\ : LocalMux
    port map (
            O => \N__39204\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt18\
        );

    \I__8302\ : InMux
    port map (
            O => \N__39201\,
            I => \N__39198\
        );

    \I__8301\ : LocalMux
    port map (
            O => \N__39198\,
            I => \N__39195\
        );

    \I__8300\ : Span4Mux_v
    port map (
            O => \N__39195\,
            I => \N__39192\
        );

    \I__8299\ : Span4Mux_h
    port map (
            O => \N__39192\,
            I => \N__39189\
        );

    \I__8298\ : Odrv4
    port map (
            O => \N__39189\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\
        );

    \I__8297\ : CascadeMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__8296\ : InMux
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__39180\,
            I => \N__39177\
        );

    \I__8294\ : Span4Mux_v
    port map (
            O => \N__39177\,
            I => \N__39174\
        );

    \I__8293\ : Odrv4
    port map (
            O => \N__39174\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt28\
        );

    \I__8292\ : InMux
    port map (
            O => \N__39171\,
            I => \N__39168\
        );

    \I__8291\ : LocalMux
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__39165\,
            I => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\
        );

    \I__8289\ : CascadeMux
    port map (
            O => \N__39162\,
            I => \N__39159\
        );

    \I__8288\ : InMux
    port map (
            O => \N__39159\,
            I => \N__39156\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__39156\,
            I => \N__39153\
        );

    \I__8286\ : Span4Mux_h
    port map (
            O => \N__39153\,
            I => \N__39150\
        );

    \I__8285\ : Odrv4
    port map (
            O => \N__39150\,
            I => \phase_controller_inst2.stoper_hc.un4_running_lt30\
        );

    \I__8284\ : CascadeMux
    port map (
            O => \N__39147\,
            I => \N__39144\
        );

    \I__8283\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39141\
        );

    \I__8282\ : LocalMux
    port map (
            O => \N__39141\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39135\
        );

    \I__8280\ : LocalMux
    port map (
            O => \N__39135\,
            I => \N__39132\
        );

    \I__8279\ : Span4Mux_v
    port map (
            O => \N__39132\,
            I => \N__39129\
        );

    \I__8278\ : Span4Mux_h
    port map (
            O => \N__39129\,
            I => \N__39126\
        );

    \I__8277\ : Odrv4
    port map (
            O => \N__39126\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\
        );

    \I__8276\ : CascadeMux
    port map (
            O => \N__39123\,
            I => \N__39120\
        );

    \I__8275\ : InMux
    port map (
            O => \N__39120\,
            I => \N__39117\
        );

    \I__8274\ : LocalMux
    port map (
            O => \N__39117\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\
        );

    \I__8273\ : CascadeMux
    port map (
            O => \N__39114\,
            I => \N__39111\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39111\,
            I => \N__39108\
        );

    \I__8271\ : LocalMux
    port map (
            O => \N__39108\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\
        );

    \I__8270\ : CascadeMux
    port map (
            O => \N__39105\,
            I => \N__39102\
        );

    \I__8269\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39099\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__39099\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39096\,
            I => \N__39093\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__39093\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__39090\,
            I => \N__39087\
        );

    \I__8264\ : InMux
    port map (
            O => \N__39087\,
            I => \N__39084\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__39084\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\
        );

    \I__8262\ : CascadeMux
    port map (
            O => \N__39081\,
            I => \N__39078\
        );

    \I__8261\ : InMux
    port map (
            O => \N__39078\,
            I => \N__39075\
        );

    \I__8260\ : LocalMux
    port map (
            O => \N__39075\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__39072\,
            I => \N__39069\
        );

    \I__8258\ : InMux
    port map (
            O => \N__39069\,
            I => \N__39066\
        );

    \I__8257\ : LocalMux
    port map (
            O => \N__39066\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39052\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39062\,
            I => \N__39052\
        );

    \I__8254\ : InMux
    port map (
            O => \N__39061\,
            I => \N__39052\
        );

    \I__8253\ : InMux
    port map (
            O => \N__39060\,
            I => \N__39047\
        );

    \I__8252\ : InMux
    port map (
            O => \N__39059\,
            I => \N__39047\
        );

    \I__8251\ : LocalMux
    port map (
            O => \N__39052\,
            I => \N__39044\
        );

    \I__8250\ : LocalMux
    port map (
            O => \N__39047\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__8249\ : Odrv4
    port map (
            O => \N__39044\,
            I => \phase_controller_inst2.stoper_hc.un2_start_0\
        );

    \I__8248\ : CascadeMux
    port map (
            O => \N__39039\,
            I => \N__39036\
        );

    \I__8247\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39030\
        );

    \I__8246\ : InMux
    port map (
            O => \N__39035\,
            I => \N__39030\
        );

    \I__8245\ : LocalMux
    port map (
            O => \N__39030\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\
        );

    \I__8244\ : CascadeMux
    port map (
            O => \N__39027\,
            I => \N__39023\
        );

    \I__8243\ : CascadeMux
    port map (
            O => \N__39026\,
            I => \N__39020\
        );

    \I__8242\ : InMux
    port map (
            O => \N__39023\,
            I => \N__39013\
        );

    \I__8241\ : InMux
    port map (
            O => \N__39020\,
            I => \N__39013\
        );

    \I__8240\ : InMux
    port map (
            O => \N__39019\,
            I => \N__39008\
        );

    \I__8239\ : InMux
    port map (
            O => \N__39018\,
            I => \N__39008\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__39013\,
            I => \N__39005\
        );

    \I__8237\ : LocalMux
    port map (
            O => \N__39008\,
            I => \N__39002\
        );

    \I__8236\ : Span4Mux_h
    port map (
            O => \N__39005\,
            I => \N__38998\
        );

    \I__8235\ : Span4Mux_h
    port map (
            O => \N__39002\,
            I => \N__38995\
        );

    \I__8234\ : InMux
    port map (
            O => \N__39001\,
            I => \N__38992\
        );

    \I__8233\ : Odrv4
    port map (
            O => \N__38998\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8232\ : Odrv4
    port map (
            O => \N__38995\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8231\ : LocalMux
    port map (
            O => \N__38992\,
            I => \phase_controller_inst2.stoper_hc.start_latchedZ0\
        );

    \I__8230\ : InMux
    port map (
            O => \N__38985\,
            I => \N__38981\
        );

    \I__8229\ : InMux
    port map (
            O => \N__38984\,
            I => \N__38976\
        );

    \I__8228\ : LocalMux
    port map (
            O => \N__38981\,
            I => \N__38973\
        );

    \I__8227\ : InMux
    port map (
            O => \N__38980\,
            I => \N__38970\
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__38979\,
            I => \N__38967\
        );

    \I__8225\ : LocalMux
    port map (
            O => \N__38976\,
            I => \N__38960\
        );

    \I__8224\ : Span4Mux_v
    port map (
            O => \N__38973\,
            I => \N__38960\
        );

    \I__8223\ : LocalMux
    port map (
            O => \N__38970\,
            I => \N__38960\
        );

    \I__8222\ : InMux
    port map (
            O => \N__38967\,
            I => \N__38957\
        );

    \I__8221\ : Span4Mux_h
    port map (
            O => \N__38960\,
            I => \N__38954\
        );

    \I__8220\ : LocalMux
    port map (
            O => \N__38957\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__38954\,
            I => \phase_controller_inst2.start_timer_hcZ0\
        );

    \I__8218\ : CascadeMux
    port map (
            O => \N__38949\,
            I => \N__38946\
        );

    \I__8217\ : InMux
    port map (
            O => \N__38946\,
            I => \N__38943\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__8215\ : Odrv4
    port map (
            O => \N__38940\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\
        );

    \I__8214\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__8213\ : LocalMux
    port map (
            O => \N__38934\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__38931\,
            I => \N__38928\
        );

    \I__8211\ : InMux
    port map (
            O => \N__38928\,
            I => \N__38925\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__38925\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\
        );

    \I__8209\ : InMux
    port map (
            O => \N__38922\,
            I => \N__38919\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__38919\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\
        );

    \I__8207\ : CascadeMux
    port map (
            O => \N__38916\,
            I => \N__38913\
        );

    \I__8206\ : InMux
    port map (
            O => \N__38913\,
            I => \N__38910\
        );

    \I__8205\ : LocalMux
    port map (
            O => \N__38910\,
            I => \N__38907\
        );

    \I__8204\ : Odrv4
    port map (
            O => \N__38907\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\
        );

    \I__8203\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38901\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__38901\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\
        );

    \I__8201\ : CascadeMux
    port map (
            O => \N__38898\,
            I => \N__38895\
        );

    \I__8200\ : InMux
    port map (
            O => \N__38895\,
            I => \N__38892\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__38892\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\
        );

    \I__8198\ : InMux
    port map (
            O => \N__38889\,
            I => \N__38886\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38886\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\
        );

    \I__8196\ : CascadeMux
    port map (
            O => \N__38883\,
            I => \N__38880\
        );

    \I__8195\ : InMux
    port map (
            O => \N__38880\,
            I => \N__38877\
        );

    \I__8194\ : LocalMux
    port map (
            O => \N__38877\,
            I => \N__38874\
        );

    \I__8193\ : Odrv4
    port map (
            O => \N__38874\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\
        );

    \I__8192\ : CascadeMux
    port map (
            O => \N__38871\,
            I => \N__38868\
        );

    \I__8191\ : InMux
    port map (
            O => \N__38868\,
            I => \N__38865\
        );

    \I__8190\ : LocalMux
    port map (
            O => \N__38865\,
            I => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38862\,
            I => \N__38845\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38861\,
            I => \N__38838\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38860\,
            I => \N__38838\
        );

    \I__8186\ : InMux
    port map (
            O => \N__38859\,
            I => \N__38838\
        );

    \I__8185\ : InMux
    port map (
            O => \N__38858\,
            I => \N__38829\
        );

    \I__8184\ : InMux
    port map (
            O => \N__38857\,
            I => \N__38829\
        );

    \I__8183\ : InMux
    port map (
            O => \N__38856\,
            I => \N__38829\
        );

    \I__8182\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38829\
        );

    \I__8181\ : CascadeMux
    port map (
            O => \N__38854\,
            I => \N__38825\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__38853\,
            I => \N__38821\
        );

    \I__8179\ : CascadeMux
    port map (
            O => \N__38852\,
            I => \N__38817\
        );

    \I__8178\ : CascadeMux
    port map (
            O => \N__38851\,
            I => \N__38812\
        );

    \I__8177\ : CascadeMux
    port map (
            O => \N__38850\,
            I => \N__38808\
        );

    \I__8176\ : CascadeMux
    port map (
            O => \N__38849\,
            I => \N__38804\
        );

    \I__8175\ : InMux
    port map (
            O => \N__38848\,
            I => \N__38800\
        );

    \I__8174\ : LocalMux
    port map (
            O => \N__38845\,
            I => \N__38793\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__38838\,
            I => \N__38793\
        );

    \I__8172\ : LocalMux
    port map (
            O => \N__38829\,
            I => \N__38793\
        );

    \I__8171\ : InMux
    port map (
            O => \N__38828\,
            I => \N__38778\
        );

    \I__8170\ : InMux
    port map (
            O => \N__38825\,
            I => \N__38778\
        );

    \I__8169\ : InMux
    port map (
            O => \N__38824\,
            I => \N__38778\
        );

    \I__8168\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38778\
        );

    \I__8167\ : InMux
    port map (
            O => \N__38820\,
            I => \N__38778\
        );

    \I__8166\ : InMux
    port map (
            O => \N__38817\,
            I => \N__38778\
        );

    \I__8165\ : InMux
    port map (
            O => \N__38816\,
            I => \N__38778\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38815\,
            I => \N__38763\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38763\
        );

    \I__8162\ : InMux
    port map (
            O => \N__38811\,
            I => \N__38763\
        );

    \I__8161\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38763\
        );

    \I__8160\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38763\
        );

    \I__8159\ : InMux
    port map (
            O => \N__38804\,
            I => \N__38763\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38803\,
            I => \N__38763\
        );

    \I__8157\ : LocalMux
    port map (
            O => \N__38800\,
            I => \N__38750\
        );

    \I__8156\ : Span4Mux_v
    port map (
            O => \N__38793\,
            I => \N__38743\
        );

    \I__8155\ : LocalMux
    port map (
            O => \N__38778\,
            I => \N__38740\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__38763\,
            I => \N__38737\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__38762\,
            I => \N__38733\
        );

    \I__8152\ : CascadeMux
    port map (
            O => \N__38761\,
            I => \N__38729\
        );

    \I__8151\ : CascadeMux
    port map (
            O => \N__38760\,
            I => \N__38725\
        );

    \I__8150\ : CascadeMux
    port map (
            O => \N__38759\,
            I => \N__38721\
        );

    \I__8149\ : InMux
    port map (
            O => \N__38758\,
            I => \N__38718\
        );

    \I__8148\ : InMux
    port map (
            O => \N__38757\,
            I => \N__38713\
        );

    \I__8147\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38713\
        );

    \I__8146\ : InMux
    port map (
            O => \N__38755\,
            I => \N__38710\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38754\,
            I => \N__38703\
        );

    \I__8144\ : InMux
    port map (
            O => \N__38753\,
            I => \N__38700\
        );

    \I__8143\ : Span4Mux_s1_h
    port map (
            O => \N__38750\,
            I => \N__38697\
        );

    \I__8142\ : CascadeMux
    port map (
            O => \N__38749\,
            I => \N__38694\
        );

    \I__8141\ : CascadeMux
    port map (
            O => \N__38748\,
            I => \N__38690\
        );

    \I__8140\ : CascadeMux
    port map (
            O => \N__38747\,
            I => \N__38686\
        );

    \I__8139\ : CascadeMux
    port map (
            O => \N__38746\,
            I => \N__38682\
        );

    \I__8138\ : Sp12to4
    port map (
            O => \N__38743\,
            I => \N__38667\
        );

    \I__8137\ : Span4Mux_v
    port map (
            O => \N__38740\,
            I => \N__38662\
        );

    \I__8136\ : Span4Mux_v
    port map (
            O => \N__38737\,
            I => \N__38662\
        );

    \I__8135\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38645\
        );

    \I__8134\ : InMux
    port map (
            O => \N__38733\,
            I => \N__38645\
        );

    \I__8133\ : InMux
    port map (
            O => \N__38732\,
            I => \N__38645\
        );

    \I__8132\ : InMux
    port map (
            O => \N__38729\,
            I => \N__38645\
        );

    \I__8131\ : InMux
    port map (
            O => \N__38728\,
            I => \N__38645\
        );

    \I__8130\ : InMux
    port map (
            O => \N__38725\,
            I => \N__38645\
        );

    \I__8129\ : InMux
    port map (
            O => \N__38724\,
            I => \N__38645\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38721\,
            I => \N__38645\
        );

    \I__8127\ : LocalMux
    port map (
            O => \N__38718\,
            I => \N__38638\
        );

    \I__8126\ : LocalMux
    port map (
            O => \N__38713\,
            I => \N__38638\
        );

    \I__8125\ : LocalMux
    port map (
            O => \N__38710\,
            I => \N__38638\
        );

    \I__8124\ : InMux
    port map (
            O => \N__38709\,
            I => \N__38635\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38708\,
            I => \N__38630\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38707\,
            I => \N__38630\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38706\,
            I => \N__38627\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38622\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38622\
        );

    \I__8118\ : Sp12to4
    port map (
            O => \N__38697\,
            I => \N__38619\
        );

    \I__8117\ : InMux
    port map (
            O => \N__38694\,
            I => \N__38602\
        );

    \I__8116\ : InMux
    port map (
            O => \N__38693\,
            I => \N__38602\
        );

    \I__8115\ : InMux
    port map (
            O => \N__38690\,
            I => \N__38602\
        );

    \I__8114\ : InMux
    port map (
            O => \N__38689\,
            I => \N__38602\
        );

    \I__8113\ : InMux
    port map (
            O => \N__38686\,
            I => \N__38602\
        );

    \I__8112\ : InMux
    port map (
            O => \N__38685\,
            I => \N__38602\
        );

    \I__8111\ : InMux
    port map (
            O => \N__38682\,
            I => \N__38602\
        );

    \I__8110\ : InMux
    port map (
            O => \N__38681\,
            I => \N__38602\
        );

    \I__8109\ : InMux
    port map (
            O => \N__38680\,
            I => \N__38599\
        );

    \I__8108\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38596\
        );

    \I__8107\ : InMux
    port map (
            O => \N__38678\,
            I => \N__38593\
        );

    \I__8106\ : InMux
    port map (
            O => \N__38677\,
            I => \N__38590\
        );

    \I__8105\ : InMux
    port map (
            O => \N__38676\,
            I => \N__38583\
        );

    \I__8104\ : InMux
    port map (
            O => \N__38675\,
            I => \N__38583\
        );

    \I__8103\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38583\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38574\
        );

    \I__8101\ : InMux
    port map (
            O => \N__38672\,
            I => \N__38574\
        );

    \I__8100\ : InMux
    port map (
            O => \N__38671\,
            I => \N__38574\
        );

    \I__8099\ : InMux
    port map (
            O => \N__38670\,
            I => \N__38574\
        );

    \I__8098\ : Span12Mux_s8_h
    port map (
            O => \N__38667\,
            I => \N__38565\
        );

    \I__8097\ : Sp12to4
    port map (
            O => \N__38662\,
            I => \N__38565\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38645\,
            I => \N__38565\
        );

    \I__8095\ : Span12Mux_s9_v
    port map (
            O => \N__38638\,
            I => \N__38556\
        );

    \I__8094\ : LocalMux
    port map (
            O => \N__38635\,
            I => \N__38556\
        );

    \I__8093\ : LocalMux
    port map (
            O => \N__38630\,
            I => \N__38556\
        );

    \I__8092\ : LocalMux
    port map (
            O => \N__38627\,
            I => \N__38556\
        );

    \I__8091\ : Span4Mux_v
    port map (
            O => \N__38622\,
            I => \N__38553\
        );

    \I__8090\ : Span12Mux_s8_v
    port map (
            O => \N__38619\,
            I => \N__38548\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__38602\,
            I => \N__38548\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__38599\,
            I => \N__38535\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__38596\,
            I => \N__38535\
        );

    \I__8086\ : LocalMux
    port map (
            O => \N__38593\,
            I => \N__38535\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38590\,
            I => \N__38535\
        );

    \I__8084\ : LocalMux
    port map (
            O => \N__38583\,
            I => \N__38535\
        );

    \I__8083\ : LocalMux
    port map (
            O => \N__38574\,
            I => \N__38535\
        );

    \I__8082\ : CascadeMux
    port map (
            O => \N__38573\,
            I => \N__38532\
        );

    \I__8081\ : CascadeMux
    port map (
            O => \N__38572\,
            I => \N__38528\
        );

    \I__8080\ : Span12Mux_h
    port map (
            O => \N__38565\,
            I => \N__38525\
        );

    \I__8079\ : Span12Mux_v
    port map (
            O => \N__38556\,
            I => \N__38516\
        );

    \I__8078\ : Sp12to4
    port map (
            O => \N__38553\,
            I => \N__38516\
        );

    \I__8077\ : Span12Mux_h
    port map (
            O => \N__38548\,
            I => \N__38516\
        );

    \I__8076\ : Span12Mux_s8_v
    port map (
            O => \N__38535\,
            I => \N__38516\
        );

    \I__8075\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38509\
        );

    \I__8074\ : InMux
    port map (
            O => \N__38531\,
            I => \N__38509\
        );

    \I__8073\ : InMux
    port map (
            O => \N__38528\,
            I => \N__38509\
        );

    \I__8072\ : Odrv12
    port map (
            O => \N__38525\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8071\ : Odrv12
    port map (
            O => \N__38516\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8070\ : LocalMux
    port map (
            O => \N__38509\,
            I => \CONSTANT_ONE_NET\
        );

    \I__8069\ : InMux
    port map (
            O => \N__38502\,
            I => \current_shift_inst.un10_control_input_cry_30\
        );

    \I__8068\ : CascadeMux
    port map (
            O => \N__38499\,
            I => \N__38486\
        );

    \I__8067\ : InMux
    port map (
            O => \N__38498\,
            I => \N__38480\
        );

    \I__8066\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38480\
        );

    \I__8065\ : InMux
    port map (
            O => \N__38496\,
            I => \N__38476\
        );

    \I__8064\ : InMux
    port map (
            O => \N__38495\,
            I => \N__38471\
        );

    \I__8063\ : InMux
    port map (
            O => \N__38494\,
            I => \N__38471\
        );

    \I__8062\ : InMux
    port map (
            O => \N__38493\,
            I => \N__38468\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__38492\,
            I => \N__38464\
        );

    \I__8060\ : InMux
    port map (
            O => \N__38491\,
            I => \N__38449\
        );

    \I__8059\ : InMux
    port map (
            O => \N__38490\,
            I => \N__38449\
        );

    \I__8058\ : InMux
    port map (
            O => \N__38489\,
            I => \N__38446\
        );

    \I__8057\ : InMux
    port map (
            O => \N__38486\,
            I => \N__38443\
        );

    \I__8056\ : InMux
    port map (
            O => \N__38485\,
            I => \N__38439\
        );

    \I__8055\ : LocalMux
    port map (
            O => \N__38480\,
            I => \N__38436\
        );

    \I__8054\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38433\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__38476\,
            I => \N__38419\
        );

    \I__8052\ : LocalMux
    port map (
            O => \N__38471\,
            I => \N__38419\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__38468\,
            I => \N__38419\
        );

    \I__8050\ : InMux
    port map (
            O => \N__38467\,
            I => \N__38406\
        );

    \I__8049\ : InMux
    port map (
            O => \N__38464\,
            I => \N__38406\
        );

    \I__8048\ : InMux
    port map (
            O => \N__38463\,
            I => \N__38406\
        );

    \I__8047\ : InMux
    port map (
            O => \N__38462\,
            I => \N__38406\
        );

    \I__8046\ : InMux
    port map (
            O => \N__38461\,
            I => \N__38406\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38460\,
            I => \N__38406\
        );

    \I__8044\ : InMux
    port map (
            O => \N__38459\,
            I => \N__38393\
        );

    \I__8043\ : InMux
    port map (
            O => \N__38458\,
            I => \N__38393\
        );

    \I__8042\ : InMux
    port map (
            O => \N__38457\,
            I => \N__38393\
        );

    \I__8041\ : InMux
    port map (
            O => \N__38456\,
            I => \N__38393\
        );

    \I__8040\ : InMux
    port map (
            O => \N__38455\,
            I => \N__38393\
        );

    \I__8039\ : InMux
    port map (
            O => \N__38454\,
            I => \N__38393\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__38449\,
            I => \N__38388\
        );

    \I__8037\ : LocalMux
    port map (
            O => \N__38446\,
            I => \N__38388\
        );

    \I__8036\ : LocalMux
    port map (
            O => \N__38443\,
            I => \N__38385\
        );

    \I__8035\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38382\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__38439\,
            I => \N__38379\
        );

    \I__8033\ : Span4Mux_v
    port map (
            O => \N__38436\,
            I => \N__38374\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__38433\,
            I => \N__38374\
        );

    \I__8031\ : InMux
    port map (
            O => \N__38432\,
            I => \N__38365\
        );

    \I__8030\ : InMux
    port map (
            O => \N__38431\,
            I => \N__38365\
        );

    \I__8029\ : InMux
    port map (
            O => \N__38430\,
            I => \N__38365\
        );

    \I__8028\ : InMux
    port map (
            O => \N__38429\,
            I => \N__38365\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38428\,
            I => \N__38358\
        );

    \I__8026\ : InMux
    port map (
            O => \N__38427\,
            I => \N__38358\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38426\,
            I => \N__38358\
        );

    \I__8024\ : Sp12to4
    port map (
            O => \N__38419\,
            I => \N__38349\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__38406\,
            I => \N__38349\
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38393\,
            I => \N__38349\
        );

    \I__8021\ : Sp12to4
    port map (
            O => \N__38388\,
            I => \N__38349\
        );

    \I__8020\ : Span4Mux_v
    port map (
            O => \N__38385\,
            I => \N__38340\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__38382\,
            I => \N__38340\
        );

    \I__8018\ : Span4Mux_h
    port map (
            O => \N__38379\,
            I => \N__38340\
        );

    \I__8017\ : Span4Mux_h
    port map (
            O => \N__38374\,
            I => \N__38340\
        );

    \I__8016\ : LocalMux
    port map (
            O => \N__38365\,
            I => \N__38335\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38358\,
            I => \N__38335\
        );

    \I__8014\ : Span12Mux_v
    port map (
            O => \N__38349\,
            I => \N__38332\
        );

    \I__8013\ : Sp12to4
    port map (
            O => \N__38340\,
            I => \N__38327\
        );

    \I__8012\ : Span12Mux_v
    port map (
            O => \N__38335\,
            I => \N__38327\
        );

    \I__8011\ : Odrv12
    port map (
            O => \N__38332\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__8010\ : Odrv12
    port map (
            O => \N__38327\,
            I => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\
        );

    \I__8009\ : CascadeMux
    port map (
            O => \N__38322\,
            I => \N__38317\
        );

    \I__8008\ : InMux
    port map (
            O => \N__38321\,
            I => \N__38313\
        );

    \I__8007\ : InMux
    port map (
            O => \N__38320\,
            I => \N__38310\
        );

    \I__8006\ : InMux
    port map (
            O => \N__38317\,
            I => \N__38307\
        );

    \I__8005\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38304\
        );

    \I__8004\ : LocalMux
    port map (
            O => \N__38313\,
            I => \N__38297\
        );

    \I__8003\ : LocalMux
    port map (
            O => \N__38310\,
            I => \N__38297\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38307\,
            I => \N__38297\
        );

    \I__8001\ : LocalMux
    port map (
            O => \N__38304\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__8000\ : Odrv12
    port map (
            O => \N__38297\,
            I => \phase_controller_inst2.hc_time_passed\
        );

    \I__7999\ : InMux
    port map (
            O => \N__38292\,
            I => \N__38288\
        );

    \I__7998\ : InMux
    port map (
            O => \N__38291\,
            I => \N__38285\
        );

    \I__7997\ : LocalMux
    port map (
            O => \N__38288\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__7996\ : LocalMux
    port map (
            O => \N__38285\,
            I => \phase_controller_inst2.stoper_hc.runningZ0\
        );

    \I__7995\ : CascadeMux
    port map (
            O => \N__38280\,
            I => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__7994\ : CascadeMux
    port map (
            O => \N__38277\,
            I => \N__38273\
        );

    \I__7993\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38268\
        );

    \I__7992\ : InMux
    port map (
            O => \N__38273\,
            I => \N__38265\
        );

    \I__7991\ : InMux
    port map (
            O => \N__38272\,
            I => \N__38260\
        );

    \I__7990\ : InMux
    port map (
            O => \N__38271\,
            I => \N__38260\
        );

    \I__7989\ : LocalMux
    port map (
            O => \N__38268\,
            I => \N__38257\
        );

    \I__7988\ : LocalMux
    port map (
            O => \N__38265\,
            I => \N__38254\
        );

    \I__7987\ : LocalMux
    port map (
            O => \N__38260\,
            I => \N__38250\
        );

    \I__7986\ : Span4Mux_v
    port map (
            O => \N__38257\,
            I => \N__38244\
        );

    \I__7985\ : Span4Mux_h
    port map (
            O => \N__38254\,
            I => \N__38244\
        );

    \I__7984\ : InMux
    port map (
            O => \N__38253\,
            I => \N__38241\
        );

    \I__7983\ : Span12Mux_v
    port map (
            O => \N__38250\,
            I => \N__38238\
        );

    \I__7982\ : InMux
    port map (
            O => \N__38249\,
            I => \N__38235\
        );

    \I__7981\ : Odrv4
    port map (
            O => \N__38244\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38241\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7979\ : Odrv12
    port map (
            O => \N__38238\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__38235\,
            I => \current_shift_inst.elapsed_time_ns_s1_i_31\
        );

    \I__7977\ : InMux
    port map (
            O => \N__38226\,
            I => \N__38223\
        );

    \I__7976\ : LocalMux
    port map (
            O => \N__38223\,
            I => \N__38220\
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__38220\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\
        );

    \I__7974\ : CascadeMux
    port map (
            O => \N__38217\,
            I => \N__38214\
        );

    \I__7973\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38211\
        );

    \I__7972\ : LocalMux
    port map (
            O => \N__38211\,
            I => \N__38208\
        );

    \I__7971\ : Odrv4
    port map (
            O => \N__38208\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\
        );

    \I__7970\ : InMux
    port map (
            O => \N__38205\,
            I => \N__38202\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__38202\,
            I => \N__38199\
        );

    \I__7968\ : Odrv4
    port map (
            O => \N__38199\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\
        );

    \I__7967\ : CascadeMux
    port map (
            O => \N__38196\,
            I => \N__38193\
        );

    \I__7966\ : InMux
    port map (
            O => \N__38193\,
            I => \N__38190\
        );

    \I__7965\ : LocalMux
    port map (
            O => \N__38190\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__38187\,
            I => \N__38184\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38184\,
            I => \N__38181\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__38181\,
            I => \N__38178\
        );

    \I__7961\ : Odrv4
    port map (
            O => \N__38178\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\
        );

    \I__7960\ : CascadeMux
    port map (
            O => \N__38175\,
            I => \N__38172\
        );

    \I__7959\ : InMux
    port map (
            O => \N__38172\,
            I => \N__38169\
        );

    \I__7958\ : LocalMux
    port map (
            O => \N__38169\,
            I => \N__38166\
        );

    \I__7957\ : Odrv4
    port map (
            O => \N__38166\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38163\,
            I => \N__38160\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__38160\,
            I => \N__38157\
        );

    \I__7954\ : Odrv12
    port map (
            O => \N__38157\,
            I => \current_shift_inst.un38_control_input_0_s1_7\
        );

    \I__7953\ : InMux
    port map (
            O => \N__38154\,
            I => \N__38151\
        );

    \I__7952\ : LocalMux
    port map (
            O => \N__38151\,
            I => \N__38148\
        );

    \I__7951\ : Odrv4
    port map (
            O => \N__38148\,
            I => \current_shift_inst.un38_control_input_0_s0_7\
        );

    \I__7950\ : InMux
    port map (
            O => \N__38145\,
            I => \N__38142\
        );

    \I__7949\ : LocalMux
    port map (
            O => \N__38142\,
            I => \N__38139\
        );

    \I__7948\ : Span4Mux_h
    port map (
            O => \N__38139\,
            I => \N__38136\
        );

    \I__7947\ : Odrv4
    port map (
            O => \N__38136\,
            I => \current_shift_inst.control_input_axb_4\
        );

    \I__7946\ : CascadeMux
    port map (
            O => \N__38133\,
            I => \N__38130\
        );

    \I__7945\ : InMux
    port map (
            O => \N__38130\,
            I => \N__38127\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__38127\,
            I => \N__38124\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__38124\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\
        );

    \I__7942\ : InMux
    port map (
            O => \N__38121\,
            I => \N__38118\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__38118\,
            I => \N__38115\
        );

    \I__7940\ : Odrv4
    port map (
            O => \N__38115\,
            I => \current_shift_inst.un38_control_input_0_s0_10\
        );

    \I__7939\ : InMux
    port map (
            O => \N__38112\,
            I => \N__38109\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__38109\,
            I => \N__38106\
        );

    \I__7937\ : Span4Mux_h
    port map (
            O => \N__38106\,
            I => \N__38103\
        );

    \I__7936\ : Odrv4
    port map (
            O => \N__38103\,
            I => \current_shift_inst.un38_control_input_0_s1_10\
        );

    \I__7935\ : InMux
    port map (
            O => \N__38100\,
            I => \N__38097\
        );

    \I__7934\ : LocalMux
    port map (
            O => \N__38097\,
            I => \N__38094\
        );

    \I__7933\ : Span4Mux_h
    port map (
            O => \N__38094\,
            I => \N__38091\
        );

    \I__7932\ : Odrv4
    port map (
            O => \N__38091\,
            I => \current_shift_inst.control_input_axb_7\
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38085\,
            I => \N__38082\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__38082\,
            I => \N__38079\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__38079\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\
        );

    \I__7927\ : InMux
    port map (
            O => \N__38076\,
            I => \N__38073\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__38073\,
            I => \N__38070\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__38070\,
            I => \current_shift_inst.un38_control_input_0_s0_11\
        );

    \I__7924\ : CascadeMux
    port map (
            O => \N__38067\,
            I => \N__38064\
        );

    \I__7923\ : InMux
    port map (
            O => \N__38064\,
            I => \N__38061\
        );

    \I__7922\ : LocalMux
    port map (
            O => \N__38061\,
            I => \N__38058\
        );

    \I__7921\ : Span4Mux_h
    port map (
            O => \N__38058\,
            I => \N__38055\
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__38055\,
            I => \current_shift_inst.un38_control_input_0_s1_11\
        );

    \I__7919\ : InMux
    port map (
            O => \N__38052\,
            I => \N__38049\
        );

    \I__7918\ : LocalMux
    port map (
            O => \N__38049\,
            I => \N__38046\
        );

    \I__7917\ : Span4Mux_v
    port map (
            O => \N__38046\,
            I => \N__38043\
        );

    \I__7916\ : Odrv4
    port map (
            O => \N__38043\,
            I => \current_shift_inst.control_input_axb_8\
        );

    \I__7915\ : InMux
    port map (
            O => \N__38040\,
            I => \N__38037\
        );

    \I__7914\ : LocalMux
    port map (
            O => \N__38037\,
            I => \N__38034\
        );

    \I__7913\ : Odrv4
    port map (
            O => \N__38034\,
            I => \current_shift_inst.un38_control_input_0_s0_6\
        );

    \I__7912\ : InMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__7911\ : LocalMux
    port map (
            O => \N__38028\,
            I => \N__38025\
        );

    \I__7910\ : Odrv4
    port map (
            O => \N__38025\,
            I => \current_shift_inst.un38_control_input_0_s1_6\
        );

    \I__7909\ : InMux
    port map (
            O => \N__38022\,
            I => \N__38019\
        );

    \I__7908\ : LocalMux
    port map (
            O => \N__38019\,
            I => \N__38016\
        );

    \I__7907\ : Span4Mux_h
    port map (
            O => \N__38016\,
            I => \N__38013\
        );

    \I__7906\ : Odrv4
    port map (
            O => \N__38013\,
            I => \current_shift_inst.control_input_axb_3\
        );

    \I__7905\ : CascadeMux
    port map (
            O => \N__38010\,
            I => \N__38007\
        );

    \I__7904\ : InMux
    port map (
            O => \N__38007\,
            I => \N__38004\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__38004\,
            I => \N__38001\
        );

    \I__7902\ : Odrv4
    port map (
            O => \N__38001\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\
        );

    \I__7901\ : InMux
    port map (
            O => \N__37998\,
            I => \N__37995\
        );

    \I__7900\ : LocalMux
    port map (
            O => \N__37995\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\
        );

    \I__7899\ : InMux
    port map (
            O => \N__37992\,
            I => \N__37989\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__37989\,
            I => \N__37986\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__37986\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\
        );

    \I__7896\ : CascadeMux
    port map (
            O => \N__37983\,
            I => \N__37980\
        );

    \I__7895\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__37977\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\
        );

    \I__7893\ : CascadeMux
    port map (
            O => \N__37974\,
            I => \N__37971\
        );

    \I__7892\ : InMux
    port map (
            O => \N__37971\,
            I => \N__37968\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__37968\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\
        );

    \I__7890\ : InMux
    port map (
            O => \N__37965\,
            I => \N__37962\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__37962\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\
        );

    \I__7888\ : CascadeMux
    port map (
            O => \N__37959\,
            I => \N__37956\
        );

    \I__7887\ : InMux
    port map (
            O => \N__37956\,
            I => \N__37953\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__37953\,
            I => \N__37950\
        );

    \I__7885\ : Span4Mux_h
    port map (
            O => \N__37950\,
            I => \N__37947\
        );

    \I__7884\ : Odrv4
    port map (
            O => \N__37947\,
            I => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\
        );

    \I__7883\ : CascadeMux
    port map (
            O => \N__37944\,
            I => \N__37941\
        );

    \I__7882\ : InMux
    port map (
            O => \N__37941\,
            I => \N__37938\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37938\,
            I => \N__37935\
        );

    \I__7880\ : Odrv4
    port map (
            O => \N__37935\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\
        );

    \I__7879\ : CascadeMux
    port map (
            O => \N__37932\,
            I => \N__37929\
        );

    \I__7878\ : InMux
    port map (
            O => \N__37929\,
            I => \N__37926\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__37926\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\
        );

    \I__7876\ : InMux
    port map (
            O => \N__37923\,
            I => \N__37920\
        );

    \I__7875\ : LocalMux
    port map (
            O => \N__37920\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\
        );

    \I__7874\ : InMux
    port map (
            O => \N__37917\,
            I => \N__37914\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__37914\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\
        );

    \I__7872\ : InMux
    port map (
            O => \N__37911\,
            I => \N__37908\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__37908\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\
        );

    \I__7870\ : InMux
    port map (
            O => \N__37905\,
            I => \N__37902\
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__37902\,
            I => \N__37897\
        );

    \I__7868\ : InMux
    port map (
            O => \N__37901\,
            I => \N__37894\
        );

    \I__7867\ : InMux
    port map (
            O => \N__37900\,
            I => \N__37891\
        );

    \I__7866\ : Span4Mux_v
    port map (
            O => \N__37897\,
            I => \N__37886\
        );

    \I__7865\ : LocalMux
    port map (
            O => \N__37894\,
            I => \N__37886\
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__37891\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7863\ : Odrv4
    port map (
            O => \N__37886\,
            I => \elapsed_time_ns_1_RNIK63T9_0_8\
        );

    \I__7862\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37878\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37878\,
            I => \N__37875\
        );

    \I__7860\ : Span4Mux_h
    port map (
            O => \N__37875\,
            I => \N__37872\
        );

    \I__7859\ : Span4Mux_v
    port map (
            O => \N__37872\,
            I => \N__37869\
        );

    \I__7858\ : Odrv4
    port map (
            O => \N__37869\,
            I => \current_shift_inst.un38_control_input_0_s1_8\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37863\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37863\,
            I => \current_shift_inst.un38_control_input_0_s0_8\
        );

    \I__7855\ : InMux
    port map (
            O => \N__37860\,
            I => \N__37857\
        );

    \I__7854\ : LocalMux
    port map (
            O => \N__37857\,
            I => \N__37854\
        );

    \I__7853\ : Span4Mux_h
    port map (
            O => \N__37854\,
            I => \N__37851\
        );

    \I__7852\ : Odrv4
    port map (
            O => \N__37851\,
            I => \current_shift_inst.control_input_axb_5\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37848\,
            I => \N__37845\
        );

    \I__7850\ : LocalMux
    port map (
            O => \N__37845\,
            I => \current_shift_inst.un38_control_input_0_s0_3\
        );

    \I__7849\ : InMux
    port map (
            O => \N__37842\,
            I => \N__37839\
        );

    \I__7848\ : LocalMux
    port map (
            O => \N__37839\,
            I => \N__37836\
        );

    \I__7847\ : Span4Mux_h
    port map (
            O => \N__37836\,
            I => \N__37833\
        );

    \I__7846\ : Odrv4
    port map (
            O => \N__37833\,
            I => \current_shift_inst.un38_control_input_0_s1_3\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37830\,
            I => \N__37826\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37829\,
            I => \N__37823\
        );

    \I__7843\ : LocalMux
    port map (
            O => \N__37826\,
            I => \N__37818\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__37823\,
            I => \N__37818\
        );

    \I__7841\ : Odrv12
    port map (
            O => \N__37818\,
            I => \current_shift_inst.control_input_axb_0\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37815\,
            I => \N__37812\
        );

    \I__7839\ : LocalMux
    port map (
            O => \N__37812\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\
        );

    \I__7838\ : CascadeMux
    port map (
            O => \N__37809\,
            I => \N__37806\
        );

    \I__7837\ : InMux
    port map (
            O => \N__37806\,
            I => \N__37803\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37803\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\
        );

    \I__7835\ : InMux
    port map (
            O => \N__37800\,
            I => \N__37797\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37797\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__37794\,
            I => \N__37791\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37791\,
            I => \N__37788\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37788\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37782\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__37782\,
            I => \N__37779\
        );

    \I__7828\ : Odrv12
    port map (
            O => \N__37779\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\
        );

    \I__7827\ : CascadeMux
    port map (
            O => \N__37776\,
            I => \N__37773\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37773\,
            I => \N__37770\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__37770\,
            I => \N__37767\
        );

    \I__7824\ : Span4Mux_v
    port map (
            O => \N__37767\,
            I => \N__37764\
        );

    \I__7823\ : Span4Mux_h
    port map (
            O => \N__37764\,
            I => \N__37761\
        );

    \I__7822\ : Odrv4
    port map (
            O => \N__37761\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt22\
        );

    \I__7821\ : CascadeMux
    port map (
            O => \N__37758\,
            I => \N__37754\
        );

    \I__7820\ : InMux
    port map (
            O => \N__37757\,
            I => \N__37748\
        );

    \I__7819\ : InMux
    port map (
            O => \N__37754\,
            I => \N__37748\
        );

    \I__7818\ : InMux
    port map (
            O => \N__37753\,
            I => \N__37745\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37748\,
            I => \N__37742\
        );

    \I__7816\ : LocalMux
    port map (
            O => \N__37745\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__7815\ : Odrv4
    port map (
            O => \N__37742\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\
        );

    \I__7814\ : CascadeMux
    port map (
            O => \N__37737\,
            I => \N__37733\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37736\,
            I => \N__37727\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37733\,
            I => \N__37727\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37732\,
            I => \N__37724\
        );

    \I__7810\ : LocalMux
    port map (
            O => \N__37727\,
            I => \N__37721\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__37724\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__7808\ : Odrv4
    port map (
            O => \N__37721\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37716\,
            I => \N__37713\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__37713\,
            I => \N__37710\
        );

    \I__7805\ : Span4Mux_h
    port map (
            O => \N__37710\,
            I => \N__37707\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__37707\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\
        );

    \I__7803\ : InMux
    port map (
            O => \N__37704\,
            I => \N__37698\
        );

    \I__7802\ : InMux
    port map (
            O => \N__37703\,
            I => \N__37698\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__37698\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\
        );

    \I__7800\ : CascadeMux
    port map (
            O => \N__37695\,
            I => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\
        );

    \I__7799\ : InMux
    port map (
            O => \N__37692\,
            I => \N__37686\
        );

    \I__7798\ : InMux
    port map (
            O => \N__37691\,
            I => \N__37686\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37686\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\
        );

    \I__7796\ : InMux
    port map (
            O => \N__37683\,
            I => \N__37680\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__37680\,
            I => \N__37676\
        );

    \I__7794\ : InMux
    port map (
            O => \N__37679\,
            I => \N__37672\
        );

    \I__7793\ : Span4Mux_h
    port map (
            O => \N__37676\,
            I => \N__37669\
        );

    \I__7792\ : InMux
    port map (
            O => \N__37675\,
            I => \N__37666\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37672\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__7790\ : Odrv4
    port map (
            O => \N__37669\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37666\,
            I => \elapsed_time_ns_1_RNIG23T9_0_4\
        );

    \I__7788\ : InMux
    port map (
            O => \N__37659\,
            I => \N__37656\
        );

    \I__7787\ : LocalMux
    port map (
            O => \N__37656\,
            I => \N__37653\
        );

    \I__7786\ : Span4Mux_h
    port map (
            O => \N__37653\,
            I => \N__37650\
        );

    \I__7785\ : Span4Mux_v
    port map (
            O => \N__37650\,
            I => \N__37647\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__37647\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\
        );

    \I__7783\ : CEMux
    port map (
            O => \N__37644\,
            I => \N__37635\
        );

    \I__7782\ : CEMux
    port map (
            O => \N__37643\,
            I => \N__37631\
        );

    \I__7781\ : CEMux
    port map (
            O => \N__37642\,
            I => \N__37616\
        );

    \I__7780\ : CEMux
    port map (
            O => \N__37641\,
            I => \N__37613\
        );

    \I__7779\ : CEMux
    port map (
            O => \N__37640\,
            I => \N__37604\
        );

    \I__7778\ : CEMux
    port map (
            O => \N__37639\,
            I => \N__37601\
        );

    \I__7777\ : CEMux
    port map (
            O => \N__37638\,
            I => \N__37598\
        );

    \I__7776\ : LocalMux
    port map (
            O => \N__37635\,
            I => \N__37594\
        );

    \I__7775\ : CEMux
    port map (
            O => \N__37634\,
            I => \N__37591\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37631\,
            I => \N__37580\
        );

    \I__7773\ : CEMux
    port map (
            O => \N__37630\,
            I => \N__37577\
        );

    \I__7772\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37568\
        );

    \I__7771\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37568\
        );

    \I__7770\ : InMux
    port map (
            O => \N__37627\,
            I => \N__37568\
        );

    \I__7769\ : InMux
    port map (
            O => \N__37626\,
            I => \N__37568\
        );

    \I__7768\ : InMux
    port map (
            O => \N__37625\,
            I => \N__37559\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37624\,
            I => \N__37559\
        );

    \I__7766\ : InMux
    port map (
            O => \N__37623\,
            I => \N__37559\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37622\,
            I => \N__37559\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37621\,
            I => \N__37548\
        );

    \I__7763\ : InMux
    port map (
            O => \N__37620\,
            I => \N__37548\
        );

    \I__7762\ : InMux
    port map (
            O => \N__37619\,
            I => \N__37548\
        );

    \I__7761\ : LocalMux
    port map (
            O => \N__37616\,
            I => \N__37543\
        );

    \I__7760\ : LocalMux
    port map (
            O => \N__37613\,
            I => \N__37543\
        );

    \I__7759\ : InMux
    port map (
            O => \N__37612\,
            I => \N__37534\
        );

    \I__7758\ : InMux
    port map (
            O => \N__37611\,
            I => \N__37534\
        );

    \I__7757\ : InMux
    port map (
            O => \N__37610\,
            I => \N__37534\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37609\,
            I => \N__37534\
        );

    \I__7755\ : CEMux
    port map (
            O => \N__37608\,
            I => \N__37531\
        );

    \I__7754\ : CEMux
    port map (
            O => \N__37607\,
            I => \N__37528\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__37604\,
            I => \N__37525\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__37601\,
            I => \N__37520\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__37598\,
            I => \N__37520\
        );

    \I__7750\ : CEMux
    port map (
            O => \N__37597\,
            I => \N__37515\
        );

    \I__7749\ : Span4Mux_v
    port map (
            O => \N__37594\,
            I => \N__37510\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__37591\,
            I => \N__37510\
        );

    \I__7747\ : InMux
    port map (
            O => \N__37590\,
            I => \N__37503\
        );

    \I__7746\ : InMux
    port map (
            O => \N__37589\,
            I => \N__37496\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37588\,
            I => \N__37496\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37587\,
            I => \N__37496\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37586\,
            I => \N__37487\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37585\,
            I => \N__37487\
        );

    \I__7741\ : InMux
    port map (
            O => \N__37584\,
            I => \N__37487\
        );

    \I__7740\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37487\
        );

    \I__7739\ : Span4Mux_v
    port map (
            O => \N__37580\,
            I => \N__37478\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37577\,
            I => \N__37478\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__37568\,
            I => \N__37478\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37559\,
            I => \N__37478\
        );

    \I__7735\ : InMux
    port map (
            O => \N__37558\,
            I => \N__37469\
        );

    \I__7734\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37469\
        );

    \I__7733\ : InMux
    port map (
            O => \N__37556\,
            I => \N__37469\
        );

    \I__7732\ : InMux
    port map (
            O => \N__37555\,
            I => \N__37469\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__37548\,
            I => \N__37460\
        );

    \I__7730\ : Span4Mux_v
    port map (
            O => \N__37543\,
            I => \N__37460\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__37534\,
            I => \N__37460\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__37531\,
            I => \N__37460\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__37528\,
            I => \N__37457\
        );

    \I__7726\ : Span4Mux_h
    port map (
            O => \N__37525\,
            I => \N__37454\
        );

    \I__7725\ : Span4Mux_v
    port map (
            O => \N__37520\,
            I => \N__37451\
        );

    \I__7724\ : CEMux
    port map (
            O => \N__37519\,
            I => \N__37448\
        );

    \I__7723\ : CEMux
    port map (
            O => \N__37518\,
            I => \N__37445\
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__37515\,
            I => \N__37442\
        );

    \I__7721\ : Span4Mux_v
    port map (
            O => \N__37510\,
            I => \N__37439\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37509\,
            I => \N__37430\
        );

    \I__7719\ : InMux
    port map (
            O => \N__37508\,
            I => \N__37430\
        );

    \I__7718\ : InMux
    port map (
            O => \N__37507\,
            I => \N__37430\
        );

    \I__7717\ : InMux
    port map (
            O => \N__37506\,
            I => \N__37430\
        );

    \I__7716\ : LocalMux
    port map (
            O => \N__37503\,
            I => \N__37427\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__37496\,
            I => \N__37416\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37487\,
            I => \N__37416\
        );

    \I__7713\ : Span4Mux_v
    port map (
            O => \N__37478\,
            I => \N__37416\
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__37469\,
            I => \N__37416\
        );

    \I__7711\ : Span4Mux_v
    port map (
            O => \N__37460\,
            I => \N__37416\
        );

    \I__7710\ : Span4Mux_v
    port map (
            O => \N__37457\,
            I => \N__37409\
        );

    \I__7709\ : Span4Mux_v
    port map (
            O => \N__37454\,
            I => \N__37409\
        );

    \I__7708\ : Span4Mux_v
    port map (
            O => \N__37451\,
            I => \N__37409\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__37448\,
            I => \N__37404\
        );

    \I__7706\ : LocalMux
    port map (
            O => \N__37445\,
            I => \N__37404\
        );

    \I__7705\ : Span4Mux_h
    port map (
            O => \N__37442\,
            I => \N__37397\
        );

    \I__7704\ : Span4Mux_h
    port map (
            O => \N__37439\,
            I => \N__37397\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__37430\,
            I => \N__37397\
        );

    \I__7702\ : Span4Mux_v
    port map (
            O => \N__37427\,
            I => \N__37392\
        );

    \I__7701\ : Span4Mux_v
    port map (
            O => \N__37416\,
            I => \N__37392\
        );

    \I__7700\ : Span4Mux_v
    port map (
            O => \N__37409\,
            I => \N__37389\
        );

    \I__7699\ : Odrv12
    port map (
            O => \N__37404\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7698\ : Odrv4
    port map (
            O => \N__37397\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7697\ : Odrv4
    port map (
            O => \N__37392\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7696\ : Odrv4
    port map (
            O => \N__37389\,
            I => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\
        );

    \I__7695\ : CascadeMux
    port map (
            O => \N__37380\,
            I => \N__37377\
        );

    \I__7694\ : InMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__37374\,
            I => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\
        );

    \I__7692\ : InMux
    port map (
            O => \N__37371\,
            I => \N__37368\
        );

    \I__7691\ : LocalMux
    port map (
            O => \N__37368\,
            I => \current_shift_inst.un38_control_input_0_s0_4\
        );

    \I__7690\ : InMux
    port map (
            O => \N__37365\,
            I => \N__37362\
        );

    \I__7689\ : LocalMux
    port map (
            O => \N__37362\,
            I => \N__37359\
        );

    \I__7688\ : Span4Mux_v
    port map (
            O => \N__37359\,
            I => \N__37356\
        );

    \I__7687\ : Odrv4
    port map (
            O => \N__37356\,
            I => \current_shift_inst.un38_control_input_0_s1_4\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__7685\ : LocalMux
    port map (
            O => \N__37350\,
            I => \N__37347\
        );

    \I__7684\ : Span4Mux_h
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__7683\ : Odrv4
    port map (
            O => \N__37344\,
            I => \current_shift_inst.control_input_axb_1\
        );

    \I__7682\ : CascadeMux
    port map (
            O => \N__37341\,
            I => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37338\,
            I => \N__37332\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37337\,
            I => \N__37332\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37332\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\
        );

    \I__7678\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37324\
        );

    \I__7677\ : InMux
    port map (
            O => \N__37328\,
            I => \N__37319\
        );

    \I__7676\ : InMux
    port map (
            O => \N__37327\,
            I => \N__37319\
        );

    \I__7675\ : LocalMux
    port map (
            O => \N__37324\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__37319\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\
        );

    \I__7673\ : CascadeMux
    port map (
            O => \N__37314\,
            I => \N__37310\
        );

    \I__7672\ : CascadeMux
    port map (
            O => \N__37313\,
            I => \N__37307\
        );

    \I__7671\ : InMux
    port map (
            O => \N__37310\,
            I => \N__37302\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37307\,
            I => \N__37302\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__37302\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\
        );

    \I__7668\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37294\
        );

    \I__7667\ : InMux
    port map (
            O => \N__37298\,
            I => \N__37289\
        );

    \I__7666\ : InMux
    port map (
            O => \N__37297\,
            I => \N__37289\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__37294\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37289\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\
        );

    \I__7663\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37281\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__37281\,
            I => \N__37278\
        );

    \I__7661\ : Odrv4
    port map (
            O => \N__37278\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\
        );

    \I__7660\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37272\
        );

    \I__7659\ : LocalMux
    port map (
            O => \N__37272\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\
        );

    \I__7658\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37266\
        );

    \I__7657\ : LocalMux
    port map (
            O => \N__37266\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\
        );

    \I__7656\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37259\
        );

    \I__7655\ : InMux
    port map (
            O => \N__37262\,
            I => \N__37255\
        );

    \I__7654\ : LocalMux
    port map (
            O => \N__37259\,
            I => \N__37252\
        );

    \I__7653\ : InMux
    port map (
            O => \N__37258\,
            I => \N__37249\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__37255\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7651\ : Odrv4
    port map (
            O => \N__37252\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7650\ : LocalMux
    port map (
            O => \N__37249\,
            I => \elapsed_time_ns_1_RNI68CN9_0_19\
        );

    \I__7649\ : InMux
    port map (
            O => \N__37242\,
            I => \N__37238\
        );

    \I__7648\ : InMux
    port map (
            O => \N__37241\,
            I => \N__37235\
        );

    \I__7647\ : LocalMux
    port map (
            O => \N__37238\,
            I => \N__37232\
        );

    \I__7646\ : LocalMux
    port map (
            O => \N__37235\,
            I => \N__37229\
        );

    \I__7645\ : Span4Mux_h
    port map (
            O => \N__37232\,
            I => \N__37226\
        );

    \I__7644\ : Odrv4
    port map (
            O => \N__37229\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__7643\ : Odrv4
    port map (
            O => \N__37226\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37217\
        );

    \I__7641\ : InMux
    port map (
            O => \N__37220\,
            I => \N__37214\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__37217\,
            I => \N__37211\
        );

    \I__7639\ : LocalMux
    port map (
            O => \N__37214\,
            I => \N__37208\
        );

    \I__7638\ : Span4Mux_v
    port map (
            O => \N__37211\,
            I => \N__37205\
        );

    \I__7637\ : Odrv4
    port map (
            O => \N__37208\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__7636\ : Odrv4
    port map (
            O => \N__37205\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37195\
        );

    \I__7634\ : InMux
    port map (
            O => \N__37199\,
            I => \N__37192\
        );

    \I__7633\ : InMux
    port map (
            O => \N__37198\,
            I => \N__37189\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__37195\,
            I => \N__37184\
        );

    \I__7631\ : LocalMux
    port map (
            O => \N__37192\,
            I => \N__37184\
        );

    \I__7630\ : LocalMux
    port map (
            O => \N__37189\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__7629\ : Odrv4
    port map (
            O => \N__37184\,
            I => \elapsed_time_ns_1_RNIE03T9_0_2\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37179\,
            I => \N__37174\
        );

    \I__7627\ : InMux
    port map (
            O => \N__37178\,
            I => \N__37169\
        );

    \I__7626\ : InMux
    port map (
            O => \N__37177\,
            I => \N__37169\
        );

    \I__7625\ : LocalMux
    port map (
            O => \N__37174\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7624\ : LocalMux
    port map (
            O => \N__37169\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\
        );

    \I__7623\ : CascadeMux
    port map (
            O => \N__37164\,
            I => \N__37160\
        );

    \I__7622\ : InMux
    port map (
            O => \N__37163\,
            I => \N__37156\
        );

    \I__7621\ : InMux
    port map (
            O => \N__37160\,
            I => \N__37151\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37151\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__37156\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7618\ : LocalMux
    port map (
            O => \N__37151\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\
        );

    \I__7617\ : InMux
    port map (
            O => \N__37146\,
            I => \N__37143\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37143\,
            I => \N__37140\
        );

    \I__7615\ : Span4Mux_h
    port map (
            O => \N__37140\,
            I => \N__37137\
        );

    \I__7614\ : Odrv4
    port map (
            O => \N__37137\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\
        );

    \I__7613\ : CascadeMux
    port map (
            O => \N__37134\,
            I => \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\
        );

    \I__7612\ : CascadeMux
    port map (
            O => \N__37131\,
            I => \N__37127\
        );

    \I__7611\ : InMux
    port map (
            O => \N__37130\,
            I => \N__37122\
        );

    \I__7610\ : InMux
    port map (
            O => \N__37127\,
            I => \N__37122\
        );

    \I__7609\ : LocalMux
    port map (
            O => \N__37122\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__37119\,
            I => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\
        );

    \I__7607\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37110\
        );

    \I__7606\ : InMux
    port map (
            O => \N__37115\,
            I => \N__37110\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__37110\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\
        );

    \I__7604\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37104\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__37104\,
            I => \N__37101\
        );

    \I__7602\ : Span4Mux_h
    port map (
            O => \N__37101\,
            I => \N__37098\
        );

    \I__7601\ : Odrv4
    port map (
            O => \N__37098\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\
        );

    \I__7600\ : InMux
    port map (
            O => \N__37095\,
            I => \N__37092\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__37092\,
            I => \N__37089\
        );

    \I__7598\ : Span4Mux_v
    port map (
            O => \N__37089\,
            I => \N__37086\
        );

    \I__7597\ : Odrv4
    port map (
            O => \N__37086\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\
        );

    \I__7596\ : CascadeMux
    port map (
            O => \N__37083\,
            I => \N__37080\
        );

    \I__7595\ : InMux
    port map (
            O => \N__37080\,
            I => \N__37077\
        );

    \I__7594\ : LocalMux
    port map (
            O => \N__37077\,
            I => \N__37074\
        );

    \I__7593\ : Odrv12
    port map (
            O => \N__37074\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt18\
        );

    \I__7592\ : CascadeMux
    port map (
            O => \N__37071\,
            I => \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\
        );

    \I__7591\ : CascadeMux
    port map (
            O => \N__37068\,
            I => \N__37064\
        );

    \I__7590\ : InMux
    port map (
            O => \N__37067\,
            I => \N__37059\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37059\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__37059\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\
        );

    \I__7587\ : CascadeMux
    port map (
            O => \N__37056\,
            I => \N__37053\
        );

    \I__7586\ : InMux
    port map (
            O => \N__37053\,
            I => \N__37047\
        );

    \I__7585\ : InMux
    port map (
            O => \N__37052\,
            I => \N__37047\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37047\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\
        );

    \I__7583\ : InMux
    port map (
            O => \N__37044\,
            I => \N__37041\
        );

    \I__7582\ : LocalMux
    port map (
            O => \N__37041\,
            I => \N__37037\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37040\,
            I => \N__37034\
        );

    \I__7580\ : Odrv4
    port map (
            O => \N__37037\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__37034\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5\
        );

    \I__7578\ : CascadeMux
    port map (
            O => \N__37029\,
            I => \N__37026\
        );

    \I__7577\ : InMux
    port map (
            O => \N__37026\,
            I => \N__37023\
        );

    \I__7576\ : LocalMux
    port map (
            O => \N__37023\,
            I => \N__37020\
        );

    \I__7575\ : Span4Mux_h
    port map (
            O => \N__37020\,
            I => \N__37017\
        );

    \I__7574\ : Odrv4
    port map (
            O => \N__37017\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt20\
        );

    \I__7573\ : CascadeMux
    port map (
            O => \N__37014\,
            I => \N__37007\
        );

    \I__7572\ : InMux
    port map (
            O => \N__37013\,
            I => \N__37004\
        );

    \I__7571\ : InMux
    port map (
            O => \N__37012\,
            I => \N__36997\
        );

    \I__7570\ : InMux
    port map (
            O => \N__37011\,
            I => \N__36997\
        );

    \I__7569\ : InMux
    port map (
            O => \N__37010\,
            I => \N__36997\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37007\,
            I => \N__36994\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__37004\,
            I => \N__36991\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__36997\,
            I => \N__36988\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__36994\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7564\ : Odrv4
    port map (
            O => \N__36991\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7563\ : Odrv4
    port map (
            O => \N__36988\,
            I => \phase_controller_inst1.stoper_hc.start_latchedZ0\
        );

    \I__7562\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36975\
        );

    \I__7561\ : InMux
    port map (
            O => \N__36980\,
            I => \N__36972\
        );

    \I__7560\ : InMux
    port map (
            O => \N__36979\,
            I => \N__36967\
        );

    \I__7559\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36967\
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__36975\,
            I => \N__36964\
        );

    \I__7557\ : LocalMux
    port map (
            O => \N__36972\,
            I => \N__36961\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__36967\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7555\ : Odrv12
    port map (
            O => \N__36964\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7554\ : Odrv4
    port map (
            O => \N__36961\,
            I => \phase_controller_inst1.start_timer_hcZ0\
        );

    \I__7553\ : CascadeMux
    port map (
            O => \N__36954\,
            I => \N__36950\
        );

    \I__7552\ : InMux
    port map (
            O => \N__36953\,
            I => \N__36945\
        );

    \I__7551\ : InMux
    port map (
            O => \N__36950\,
            I => \N__36945\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__36945\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\
        );

    \I__7549\ : CascadeMux
    port map (
            O => \N__36942\,
            I => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\
        );

    \I__7548\ : InMux
    port map (
            O => \N__36939\,
            I => \N__36936\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__36936\,
            I => \N__36933\
        );

    \I__7546\ : Span4Mux_h
    port map (
            O => \N__36933\,
            I => \N__36930\
        );

    \I__7545\ : Odrv4
    port map (
            O => \N__36930\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\
        );

    \I__7544\ : CascadeMux
    port map (
            O => \N__36927\,
            I => \N__36924\
        );

    \I__7543\ : InMux
    port map (
            O => \N__36924\,
            I => \N__36921\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__36921\,
            I => \N__36918\
        );

    \I__7541\ : Span4Mux_h
    port map (
            O => \N__36918\,
            I => \N__36915\
        );

    \I__7540\ : Odrv4
    port map (
            O => \N__36915\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36912\,
            I => \N__36907\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36911\,
            I => \N__36902\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36910\,
            I => \N__36902\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36907\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__36902\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\
        );

    \I__7534\ : CascadeMux
    port map (
            O => \N__36897\,
            I => \N__36894\
        );

    \I__7533\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36888\
        );

    \I__7532\ : InMux
    port map (
            O => \N__36893\,
            I => \N__36888\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__36888\,
            I => \N__36885\
        );

    \I__7530\ : Odrv4
    port map (
            O => \N__36885\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\
        );

    \I__7529\ : InMux
    port map (
            O => \N__36882\,
            I => \N__36875\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36875\
        );

    \I__7527\ : InMux
    port map (
            O => \N__36880\,
            I => \N__36872\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__36875\,
            I => \N__36869\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__36872\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7524\ : Odrv4
    port map (
            O => \N__36869\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\
        );

    \I__7523\ : InMux
    port map (
            O => \N__36864\,
            I => \N__36861\
        );

    \I__7522\ : LocalMux
    port map (
            O => \N__36861\,
            I => \N__36858\
        );

    \I__7521\ : Span4Mux_v
    port map (
            O => \N__36858\,
            I => \N__36855\
        );

    \I__7520\ : Odrv4
    port map (
            O => \N__36855\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt16\
        );

    \I__7519\ : CascadeMux
    port map (
            O => \N__36852\,
            I => \N__36849\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36849\,
            I => \N__36846\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__36846\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\
        );

    \I__7516\ : CascadeMux
    port map (
            O => \N__36843\,
            I => \N__36840\
        );

    \I__7515\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36837\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36837\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\
        );

    \I__7513\ : CascadeMux
    port map (
            O => \N__36834\,
            I => \N__36831\
        );

    \I__7512\ : InMux
    port map (
            O => \N__36831\,
            I => \N__36828\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36825\
        );

    \I__7510\ : Odrv4
    port map (
            O => \N__36825\,
            I => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\
        );

    \I__7509\ : InMux
    port map (
            O => \N__36822\,
            I => \N__36819\
        );

    \I__7508\ : LocalMux
    port map (
            O => \N__36819\,
            I => \current_shift_inst.un38_control_input_0_s1_24\
        );

    \I__7507\ : InMux
    port map (
            O => \N__36816\,
            I => \N__36813\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36813\,
            I => \N__36810\
        );

    \I__7505\ : Odrv12
    port map (
            O => \N__36810\,
            I => \current_shift_inst.un38_control_input_0_s0_24\
        );

    \I__7504\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36804\
        );

    \I__7503\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36801\
        );

    \I__7502\ : Span4Mux_h
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__7501\ : Odrv4
    port map (
            O => \N__36798\,
            I => \current_shift_inst.control_input_axb_21\
        );

    \I__7500\ : InMux
    port map (
            O => \N__36795\,
            I => \N__36791\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36794\,
            I => \N__36788\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__36791\,
            I => \N__36785\
        );

    \I__7497\ : LocalMux
    port map (
            O => \N__36788\,
            I => \N__36782\
        );

    \I__7496\ : Span4Mux_h
    port map (
            O => \N__36785\,
            I => \N__36779\
        );

    \I__7495\ : Odrv12
    port map (
            O => \N__36782\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7494\ : Odrv4
    port map (
            O => \N__36779\,
            I => \current_shift_inst.un38_control_input_5_0\
        );

    \I__7493\ : InMux
    port map (
            O => \N__36774\,
            I => \N__36770\
        );

    \I__7492\ : InMux
    port map (
            O => \N__36773\,
            I => \N__36767\
        );

    \I__7491\ : LocalMux
    port map (
            O => \N__36770\,
            I => \N__36764\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36759\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__36764\,
            I => \N__36756\
        );

    \I__7488\ : InMux
    port map (
            O => \N__36763\,
            I => \N__36753\
        );

    \I__7487\ : InMux
    port map (
            O => \N__36762\,
            I => \N__36750\
        );

    \I__7486\ : Span4Mux_v
    port map (
            O => \N__36759\,
            I => \N__36747\
        );

    \I__7485\ : Span4Mux_v
    port map (
            O => \N__36756\,
            I => \N__36744\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36753\,
            I => \N__36741\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36738\
        );

    \I__7482\ : Span4Mux_v
    port map (
            O => \N__36747\,
            I => \N__36733\
        );

    \I__7481\ : Span4Mux_v
    port map (
            O => \N__36744\,
            I => \N__36733\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__36741\,
            I => \N__36728\
        );

    \I__7479\ : Span4Mux_v
    port map (
            O => \N__36738\,
            I => \N__36728\
        );

    \I__7478\ : Odrv4
    port map (
            O => \N__36733\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7477\ : Odrv4
    port map (
            O => \N__36728\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\
        );

    \I__7476\ : InMux
    port map (
            O => \N__36723\,
            I => \N__36715\
        );

    \I__7475\ : CascadeMux
    port map (
            O => \N__36722\,
            I => \N__36708\
        );

    \I__7474\ : CascadeMux
    port map (
            O => \N__36721\,
            I => \N__36705\
        );

    \I__7473\ : InMux
    port map (
            O => \N__36720\,
            I => \N__36695\
        );

    \I__7472\ : InMux
    port map (
            O => \N__36719\,
            I => \N__36695\
        );

    \I__7471\ : InMux
    port map (
            O => \N__36718\,
            I => \N__36692\
        );

    \I__7470\ : LocalMux
    port map (
            O => \N__36715\,
            I => \N__36683\
        );

    \I__7469\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36667\
        );

    \I__7468\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36664\
        );

    \I__7467\ : InMux
    port map (
            O => \N__36712\,
            I => \N__36659\
        );

    \I__7466\ : InMux
    port map (
            O => \N__36711\,
            I => \N__36659\
        );

    \I__7465\ : InMux
    port map (
            O => \N__36708\,
            I => \N__36652\
        );

    \I__7464\ : InMux
    port map (
            O => \N__36705\,
            I => \N__36652\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36704\,
            I => \N__36652\
        );

    \I__7462\ : CascadeMux
    port map (
            O => \N__36703\,
            I => \N__36646\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36702\,
            I => \N__36642\
        );

    \I__7460\ : InMux
    port map (
            O => \N__36701\,
            I => \N__36625\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36700\,
            I => \N__36625\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36695\,
            I => \N__36620\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__36692\,
            I => \N__36620\
        );

    \I__7456\ : InMux
    port map (
            O => \N__36691\,
            I => \N__36613\
        );

    \I__7455\ : InMux
    port map (
            O => \N__36690\,
            I => \N__36613\
        );

    \I__7454\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36613\
        );

    \I__7453\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36610\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36687\,
            I => \N__36607\
        );

    \I__7451\ : InMux
    port map (
            O => \N__36686\,
            I => \N__36604\
        );

    \I__7450\ : Span4Mux_h
    port map (
            O => \N__36683\,
            I => \N__36599\
        );

    \I__7449\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36594\
        );

    \I__7448\ : InMux
    port map (
            O => \N__36681\,
            I => \N__36591\
        );

    \I__7447\ : InMux
    port map (
            O => \N__36680\,
            I => \N__36586\
        );

    \I__7446\ : InMux
    port map (
            O => \N__36679\,
            I => \N__36586\
        );

    \I__7445\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36573\
        );

    \I__7444\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36573\
        );

    \I__7443\ : InMux
    port map (
            O => \N__36676\,
            I => \N__36573\
        );

    \I__7442\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36573\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36674\,
            I => \N__36573\
        );

    \I__7440\ : InMux
    port map (
            O => \N__36673\,
            I => \N__36573\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36672\,
            I => \N__36570\
        );

    \I__7438\ : InMux
    port map (
            O => \N__36671\,
            I => \N__36565\
        );

    \I__7437\ : InMux
    port map (
            O => \N__36670\,
            I => \N__36565\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36667\,
            I => \N__36562\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__36664\,
            I => \N__36550\
        );

    \I__7434\ : LocalMux
    port map (
            O => \N__36659\,
            I => \N__36550\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__36652\,
            I => \N__36547\
        );

    \I__7432\ : InMux
    port map (
            O => \N__36651\,
            I => \N__36539\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36650\,
            I => \N__36530\
        );

    \I__7430\ : InMux
    port map (
            O => \N__36649\,
            I => \N__36530\
        );

    \I__7429\ : InMux
    port map (
            O => \N__36646\,
            I => \N__36530\
        );

    \I__7428\ : InMux
    port map (
            O => \N__36645\,
            I => \N__36530\
        );

    \I__7427\ : LocalMux
    port map (
            O => \N__36642\,
            I => \N__36527\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36641\,
            I => \N__36518\
        );

    \I__7425\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36518\
        );

    \I__7424\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36518\
        );

    \I__7423\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36518\
        );

    \I__7422\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36513\
        );

    \I__7421\ : InMux
    port map (
            O => \N__36636\,
            I => \N__36513\
        );

    \I__7420\ : InMux
    port map (
            O => \N__36635\,
            I => \N__36506\
        );

    \I__7419\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36506\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36633\,
            I => \N__36506\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36632\,
            I => \N__36503\
        );

    \I__7416\ : InMux
    port map (
            O => \N__36631\,
            I => \N__36498\
        );

    \I__7415\ : InMux
    port map (
            O => \N__36630\,
            I => \N__36498\
        );

    \I__7414\ : LocalMux
    port map (
            O => \N__36625\,
            I => \N__36491\
        );

    \I__7413\ : Span4Mux_v
    port map (
            O => \N__36620\,
            I => \N__36491\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__36613\,
            I => \N__36491\
        );

    \I__7411\ : LocalMux
    port map (
            O => \N__36610\,
            I => \N__36484\
        );

    \I__7410\ : LocalMux
    port map (
            O => \N__36607\,
            I => \N__36484\
        );

    \I__7409\ : LocalMux
    port map (
            O => \N__36604\,
            I => \N__36484\
        );

    \I__7408\ : InMux
    port map (
            O => \N__36603\,
            I => \N__36479\
        );

    \I__7407\ : InMux
    port map (
            O => \N__36602\,
            I => \N__36479\
        );

    \I__7406\ : Span4Mux_h
    port map (
            O => \N__36599\,
            I => \N__36474\
        );

    \I__7405\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36457\
        );

    \I__7404\ : InMux
    port map (
            O => \N__36597\,
            I => \N__36457\
        );

    \I__7403\ : LocalMux
    port map (
            O => \N__36594\,
            I => \N__36454\
        );

    \I__7402\ : LocalMux
    port map (
            O => \N__36591\,
            I => \N__36451\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__36586\,
            I => \N__36446\
        );

    \I__7400\ : LocalMux
    port map (
            O => \N__36573\,
            I => \N__36446\
        );

    \I__7399\ : LocalMux
    port map (
            O => \N__36570\,
            I => \N__36439\
        );

    \I__7398\ : LocalMux
    port map (
            O => \N__36565\,
            I => \N__36439\
        );

    \I__7397\ : Span4Mux_v
    port map (
            O => \N__36562\,
            I => \N__36439\
        );

    \I__7396\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36432\
        );

    \I__7395\ : InMux
    port map (
            O => \N__36560\,
            I => \N__36432\
        );

    \I__7394\ : InMux
    port map (
            O => \N__36559\,
            I => \N__36432\
        );

    \I__7393\ : InMux
    port map (
            O => \N__36558\,
            I => \N__36423\
        );

    \I__7392\ : InMux
    port map (
            O => \N__36557\,
            I => \N__36423\
        );

    \I__7391\ : InMux
    port map (
            O => \N__36556\,
            I => \N__36423\
        );

    \I__7390\ : InMux
    port map (
            O => \N__36555\,
            I => \N__36423\
        );

    \I__7389\ : Span4Mux_h
    port map (
            O => \N__36550\,
            I => \N__36418\
        );

    \I__7388\ : Span4Mux_s3_v
    port map (
            O => \N__36547\,
            I => \N__36418\
        );

    \I__7387\ : InMux
    port map (
            O => \N__36546\,
            I => \N__36401\
        );

    \I__7386\ : InMux
    port map (
            O => \N__36545\,
            I => \N__36401\
        );

    \I__7385\ : InMux
    port map (
            O => \N__36544\,
            I => \N__36394\
        );

    \I__7384\ : InMux
    port map (
            O => \N__36543\,
            I => \N__36394\
        );

    \I__7383\ : InMux
    port map (
            O => \N__36542\,
            I => \N__36394\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__36539\,
            I => \N__36391\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__36530\,
            I => \N__36378\
        );

    \I__7380\ : Span4Mux_h
    port map (
            O => \N__36527\,
            I => \N__36378\
        );

    \I__7379\ : LocalMux
    port map (
            O => \N__36518\,
            I => \N__36378\
        );

    \I__7378\ : LocalMux
    port map (
            O => \N__36513\,
            I => \N__36378\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__36506\,
            I => \N__36378\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__36503\,
            I => \N__36378\
        );

    \I__7375\ : LocalMux
    port map (
            O => \N__36498\,
            I => \N__36371\
        );

    \I__7374\ : Span4Mux_v
    port map (
            O => \N__36491\,
            I => \N__36371\
        );

    \I__7373\ : Span4Mux_v
    port map (
            O => \N__36484\,
            I => \N__36371\
        );

    \I__7372\ : LocalMux
    port map (
            O => \N__36479\,
            I => \N__36368\
        );

    \I__7371\ : InMux
    port map (
            O => \N__36478\,
            I => \N__36365\
        );

    \I__7370\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36362\
        );

    \I__7369\ : Span4Mux_v
    port map (
            O => \N__36474\,
            I => \N__36359\
        );

    \I__7368\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36356\
        );

    \I__7367\ : InMux
    port map (
            O => \N__36472\,
            I => \N__36353\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36471\,
            I => \N__36346\
        );

    \I__7365\ : InMux
    port map (
            O => \N__36470\,
            I => \N__36346\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36469\,
            I => \N__36346\
        );

    \I__7363\ : InMux
    port map (
            O => \N__36468\,
            I => \N__36341\
        );

    \I__7362\ : InMux
    port map (
            O => \N__36467\,
            I => \N__36341\
        );

    \I__7361\ : InMux
    port map (
            O => \N__36466\,
            I => \N__36330\
        );

    \I__7360\ : InMux
    port map (
            O => \N__36465\,
            I => \N__36330\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36464\,
            I => \N__36330\
        );

    \I__7358\ : InMux
    port map (
            O => \N__36463\,
            I => \N__36330\
        );

    \I__7357\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36330\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__36457\,
            I => \N__36327\
        );

    \I__7355\ : Span4Mux_v
    port map (
            O => \N__36454\,
            I => \N__36318\
        );

    \I__7354\ : Span4Mux_v
    port map (
            O => \N__36451\,
            I => \N__36318\
        );

    \I__7353\ : Span4Mux_v
    port map (
            O => \N__36446\,
            I => \N__36318\
        );

    \I__7352\ : Span4Mux_v
    port map (
            O => \N__36439\,
            I => \N__36318\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__36432\,
            I => \N__36311\
        );

    \I__7350\ : LocalMux
    port map (
            O => \N__36423\,
            I => \N__36311\
        );

    \I__7349\ : Span4Mux_v
    port map (
            O => \N__36418\,
            I => \N__36311\
        );

    \I__7348\ : InMux
    port map (
            O => \N__36417\,
            I => \N__36302\
        );

    \I__7347\ : InMux
    port map (
            O => \N__36416\,
            I => \N__36302\
        );

    \I__7346\ : InMux
    port map (
            O => \N__36415\,
            I => \N__36302\
        );

    \I__7345\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36302\
        );

    \I__7344\ : InMux
    port map (
            O => \N__36413\,
            I => \N__36291\
        );

    \I__7343\ : InMux
    port map (
            O => \N__36412\,
            I => \N__36291\
        );

    \I__7342\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36291\
        );

    \I__7341\ : InMux
    port map (
            O => \N__36410\,
            I => \N__36291\
        );

    \I__7340\ : InMux
    port map (
            O => \N__36409\,
            I => \N__36291\
        );

    \I__7339\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36284\
        );

    \I__7338\ : InMux
    port map (
            O => \N__36407\,
            I => \N__36284\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36406\,
            I => \N__36284\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__36401\,
            I => \N__36273\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__36394\,
            I => \N__36273\
        );

    \I__7334\ : Span4Mux_h
    port map (
            O => \N__36391\,
            I => \N__36273\
        );

    \I__7333\ : Span4Mux_v
    port map (
            O => \N__36378\,
            I => \N__36273\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__36371\,
            I => \N__36273\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__36368\,
            I => \N__36264\
        );

    \I__7330\ : LocalMux
    port map (
            O => \N__36365\,
            I => \N__36264\
        );

    \I__7329\ : LocalMux
    port map (
            O => \N__36362\,
            I => \N__36264\
        );

    \I__7328\ : Span4Mux_v
    port map (
            O => \N__36359\,
            I => \N__36264\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__36356\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__36353\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__36346\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7324\ : LocalMux
    port map (
            O => \N__36341\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__36330\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7322\ : Odrv12
    port map (
            O => \N__36327\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__36318\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7320\ : Odrv4
    port map (
            O => \N__36311\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__36302\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7318\ : LocalMux
    port map (
            O => \N__36291\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36284\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7316\ : Odrv4
    port map (
            O => \N__36273\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7315\ : Odrv4
    port map (
            O => \N__36264\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3\
        );

    \I__7314\ : InMux
    port map (
            O => \N__36237\,
            I => \N__36234\
        );

    \I__7313\ : LocalMux
    port map (
            O => \N__36234\,
            I => \N__36231\
        );

    \I__7312\ : Span4Mux_h
    port map (
            O => \N__36231\,
            I => \N__36227\
        );

    \I__7311\ : InMux
    port map (
            O => \N__36230\,
            I => \N__36224\
        );

    \I__7310\ : Span4Mux_v
    port map (
            O => \N__36227\,
            I => \N__36220\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__36224\,
            I => \N__36217\
        );

    \I__7308\ : InMux
    port map (
            O => \N__36223\,
            I => \N__36214\
        );

    \I__7307\ : Sp12to4
    port map (
            O => \N__36220\,
            I => \N__36209\
        );

    \I__7306\ : Span12Mux_h
    port map (
            O => \N__36217\,
            I => \N__36209\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__36214\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__7304\ : Odrv12
    port map (
            O => \N__36209\,
            I => \elapsed_time_ns_1_RNI4EOBB_0_17\
        );

    \I__7303\ : InMux
    port map (
            O => \N__36204\,
            I => \N__36201\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__36201\,
            I => \current_shift_inst.elapsed_time_ns_s1_fast_31\
        );

    \I__7301\ : InMux
    port map (
            O => \N__36198\,
            I => \N__36192\
        );

    \I__7300\ : InMux
    port map (
            O => \N__36197\,
            I => \N__36189\
        );

    \I__7299\ : InMux
    port map (
            O => \N__36196\,
            I => \N__36184\
        );

    \I__7298\ : InMux
    port map (
            O => \N__36195\,
            I => \N__36184\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__36192\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36189\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__36184\,
            I => \current_shift_inst.timer_s1.runningZ0\
        );

    \I__7294\ : InMux
    port map (
            O => \N__36177\,
            I => \N__36174\
        );

    \I__7293\ : LocalMux
    port map (
            O => \N__36174\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\
        );

    \I__7292\ : CascadeMux
    port map (
            O => \N__36171\,
            I => \N__36168\
        );

    \I__7291\ : InMux
    port map (
            O => \N__36168\,
            I => \N__36165\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__36165\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\
        );

    \I__7289\ : InMux
    port map (
            O => \N__36162\,
            I => \N__36159\
        );

    \I__7288\ : LocalMux
    port map (
            O => \N__36159\,
            I => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\
        );

    \I__7287\ : CascadeMux
    port map (
            O => \N__36156\,
            I => \N__36153\
        );

    \I__7286\ : InMux
    port map (
            O => \N__36153\,
            I => \N__36150\
        );

    \I__7285\ : LocalMux
    port map (
            O => \N__36150\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\
        );

    \I__7284\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36144\
        );

    \I__7283\ : LocalMux
    port map (
            O => \N__36144\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\
        );

    \I__7282\ : CascadeMux
    port map (
            O => \N__36141\,
            I => \N__36138\
        );

    \I__7281\ : InMux
    port map (
            O => \N__36138\,
            I => \N__36135\
        );

    \I__7280\ : LocalMux
    port map (
            O => \N__36135\,
            I => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\
        );

    \I__7279\ : InMux
    port map (
            O => \N__36132\,
            I => \N__36129\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__36129\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\
        );

    \I__7277\ : InMux
    port map (
            O => \N__36126\,
            I => \N__36123\
        );

    \I__7276\ : LocalMux
    port map (
            O => \N__36123\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\
        );

    \I__7275\ : InMux
    port map (
            O => \N__36120\,
            I => \N__36117\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__36117\,
            I => \N__36114\
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__36114\,
            I => \current_shift_inst.un38_control_input_0_s0_25\
        );

    \I__7272\ : InMux
    port map (
            O => \N__36111\,
            I => \N__36108\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__36108\,
            I => \current_shift_inst.un38_control_input_0_s1_25\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36105\,
            I => \N__36102\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__36102\,
            I => \N__36099\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__36099\,
            I => \N__36096\
        );

    \I__7267\ : Odrv4
    port map (
            O => \N__36096\,
            I => \current_shift_inst.control_input_axb_22\
        );

    \I__7266\ : InMux
    port map (
            O => \N__36093\,
            I => \N__36090\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__36090\,
            I => \N__36087\
        );

    \I__7264\ : Span4Mux_v
    port map (
            O => \N__36087\,
            I => \N__36084\
        );

    \I__7263\ : Odrv4
    port map (
            O => \N__36084\,
            I => \current_shift_inst.un38_control_input_0_s0_29\
        );

    \I__7262\ : InMux
    port map (
            O => \N__36081\,
            I => \current_shift_inst.un38_control_input_cry_28_s0\
        );

    \I__7261\ : InMux
    port map (
            O => \N__36078\,
            I => \N__36075\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__36075\,
            I => \N__36072\
        );

    \I__7259\ : Span4Mux_v
    port map (
            O => \N__36072\,
            I => \N__36069\
        );

    \I__7258\ : Odrv4
    port map (
            O => \N__36069\,
            I => \current_shift_inst.un38_control_input_0_s0_30\
        );

    \I__7257\ : InMux
    port map (
            O => \N__36066\,
            I => \current_shift_inst.un38_control_input_cry_29_s0\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36063\,
            I => \N__36060\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36060\,
            I => \N__36057\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__36057\,
            I => \N__36054\
        );

    \I__7253\ : Odrv4
    port map (
            O => \N__36054\,
            I => \current_shift_inst.un38_control_input_0_s1_31\
        );

    \I__7252\ : InMux
    port map (
            O => \N__36051\,
            I => \current_shift_inst.un38_control_input_cry_30_s0\
        );

    \I__7251\ : InMux
    port map (
            O => \N__36048\,
            I => \N__36045\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__36045\,
            I => \N__36042\
        );

    \I__7249\ : Odrv4
    port map (
            O => \N__36042\,
            I => \current_shift_inst.control_input_axb_28\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36039\,
            I => \N__36036\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36036\,
            I => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\
        );

    \I__7246\ : CascadeMux
    port map (
            O => \N__36033\,
            I => \N__36030\
        );

    \I__7245\ : InMux
    port map (
            O => \N__36030\,
            I => \N__36027\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__36027\,
            I => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\
        );

    \I__7243\ : InMux
    port map (
            O => \N__36024\,
            I => \N__36021\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__36021\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\
        );

    \I__7241\ : InMux
    port map (
            O => \N__36018\,
            I => \N__36015\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__36015\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\
        );

    \I__7239\ : InMux
    port map (
            O => \N__36012\,
            I => \N__36009\
        );

    \I__7238\ : LocalMux
    port map (
            O => \N__36009\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\
        );

    \I__7237\ : InMux
    port map (
            O => \N__36006\,
            I => \N__36003\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__36003\,
            I => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\
        );

    \I__7235\ : InMux
    port map (
            O => \N__36000\,
            I => \N__35997\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__35997\,
            I => \N__35994\
        );

    \I__7233\ : Span4Mux_v
    port map (
            O => \N__35994\,
            I => \N__35991\
        );

    \I__7232\ : Odrv4
    port map (
            O => \N__35991\,
            I => \current_shift_inst.un38_control_input_0_s0_21\
        );

    \I__7231\ : InMux
    port map (
            O => \N__35988\,
            I => \current_shift_inst.un38_control_input_cry_20_s0\
        );

    \I__7230\ : InMux
    port map (
            O => \N__35985\,
            I => \N__35982\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__35982\,
            I => \N__35979\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__35979\,
            I => \N__35976\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__35976\,
            I => \current_shift_inst.un38_control_input_0_s0_22\
        );

    \I__7226\ : InMux
    port map (
            O => \N__35973\,
            I => \current_shift_inst.un38_control_input_cry_21_s0\
        );

    \I__7225\ : InMux
    port map (
            O => \N__35970\,
            I => \N__35967\
        );

    \I__7224\ : LocalMux
    port map (
            O => \N__35967\,
            I => \N__35964\
        );

    \I__7223\ : Span4Mux_h
    port map (
            O => \N__35964\,
            I => \N__35961\
        );

    \I__7222\ : Odrv4
    port map (
            O => \N__35961\,
            I => \current_shift_inst.un38_control_input_0_s0_23\
        );

    \I__7221\ : InMux
    port map (
            O => \N__35958\,
            I => \current_shift_inst.un38_control_input_cry_22_s0\
        );

    \I__7220\ : InMux
    port map (
            O => \N__35955\,
            I => \bfn_14_16_0_\
        );

    \I__7219\ : InMux
    port map (
            O => \N__35952\,
            I => \current_shift_inst.un38_control_input_cry_24_s0\
        );

    \I__7218\ : InMux
    port map (
            O => \N__35949\,
            I => \N__35946\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__35946\,
            I => \N__35943\
        );

    \I__7216\ : Odrv4
    port map (
            O => \N__35943\,
            I => \current_shift_inst.un38_control_input_0_s0_26\
        );

    \I__7215\ : InMux
    port map (
            O => \N__35940\,
            I => \current_shift_inst.un38_control_input_cry_25_s0\
        );

    \I__7214\ : InMux
    port map (
            O => \N__35937\,
            I => \N__35934\
        );

    \I__7213\ : LocalMux
    port map (
            O => \N__35934\,
            I => \N__35931\
        );

    \I__7212\ : Odrv4
    port map (
            O => \N__35931\,
            I => \current_shift_inst.un38_control_input_0_s0_27\
        );

    \I__7211\ : InMux
    port map (
            O => \N__35928\,
            I => \current_shift_inst.un38_control_input_cry_26_s0\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35925\,
            I => \N__35922\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__7208\ : Span4Mux_v
    port map (
            O => \N__35919\,
            I => \N__35916\
        );

    \I__7207\ : Odrv4
    port map (
            O => \N__35916\,
            I => \current_shift_inst.un38_control_input_0_s0_28\
        );

    \I__7206\ : InMux
    port map (
            O => \N__35913\,
            I => \current_shift_inst.un38_control_input_cry_27_s0\
        );

    \I__7205\ : InMux
    port map (
            O => \N__35910\,
            I => \N__35907\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__35907\,
            I => \N__35904\
        );

    \I__7203\ : Span4Mux_v
    port map (
            O => \N__35904\,
            I => \N__35901\
        );

    \I__7202\ : Odrv4
    port map (
            O => \N__35901\,
            I => \current_shift_inst.un38_control_input_0_s0_12\
        );

    \I__7201\ : InMux
    port map (
            O => \N__35898\,
            I => \current_shift_inst.un38_control_input_cry_11_s0\
        );

    \I__7200\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35892\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__35892\,
            I => \N__35889\
        );

    \I__7198\ : Span4Mux_h
    port map (
            O => \N__35889\,
            I => \N__35886\
        );

    \I__7197\ : Odrv4
    port map (
            O => \N__35886\,
            I => \current_shift_inst.un38_control_input_0_s0_13\
        );

    \I__7196\ : InMux
    port map (
            O => \N__35883\,
            I => \current_shift_inst.un38_control_input_cry_12_s0\
        );

    \I__7195\ : InMux
    port map (
            O => \N__35880\,
            I => \N__35877\
        );

    \I__7194\ : LocalMux
    port map (
            O => \N__35877\,
            I => \N__35874\
        );

    \I__7193\ : Span4Mux_h
    port map (
            O => \N__35874\,
            I => \N__35871\
        );

    \I__7192\ : Odrv4
    port map (
            O => \N__35871\,
            I => \current_shift_inst.un38_control_input_0_s0_14\
        );

    \I__7191\ : InMux
    port map (
            O => \N__35868\,
            I => \current_shift_inst.un38_control_input_cry_13_s0\
        );

    \I__7190\ : InMux
    port map (
            O => \N__35865\,
            I => \N__35862\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__35862\,
            I => \N__35859\
        );

    \I__7188\ : Span4Mux_h
    port map (
            O => \N__35859\,
            I => \N__35856\
        );

    \I__7187\ : Odrv4
    port map (
            O => \N__35856\,
            I => \current_shift_inst.un38_control_input_0_s0_15\
        );

    \I__7186\ : InMux
    port map (
            O => \N__35853\,
            I => \current_shift_inst.un38_control_input_cry_14_s0\
        );

    \I__7185\ : InMux
    port map (
            O => \N__35850\,
            I => \N__35847\
        );

    \I__7184\ : LocalMux
    port map (
            O => \N__35847\,
            I => \N__35844\
        );

    \I__7183\ : Odrv4
    port map (
            O => \N__35844\,
            I => \current_shift_inst.un38_control_input_0_s0_16\
        );

    \I__7182\ : InMux
    port map (
            O => \N__35841\,
            I => \bfn_14_15_0_\
        );

    \I__7181\ : InMux
    port map (
            O => \N__35838\,
            I => \N__35835\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__35835\,
            I => \N__35832\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__35832\,
            I => \current_shift_inst.un38_control_input_0_s0_17\
        );

    \I__7178\ : InMux
    port map (
            O => \N__35829\,
            I => \current_shift_inst.un38_control_input_cry_16_s0\
        );

    \I__7177\ : InMux
    port map (
            O => \N__35826\,
            I => \N__35823\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__35823\,
            I => \N__35820\
        );

    \I__7175\ : Odrv4
    port map (
            O => \N__35820\,
            I => \current_shift_inst.un38_control_input_0_s0_18\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35817\,
            I => \current_shift_inst.un38_control_input_cry_17_s0\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35814\,
            I => \N__35811\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__35811\,
            I => \N__35808\
        );

    \I__7171\ : Span4Mux_h
    port map (
            O => \N__35808\,
            I => \N__35805\
        );

    \I__7170\ : Odrv4
    port map (
            O => \N__35805\,
            I => \current_shift_inst.un38_control_input_0_s0_19\
        );

    \I__7169\ : InMux
    port map (
            O => \N__35802\,
            I => \current_shift_inst.un38_control_input_cry_18_s0\
        );

    \I__7168\ : InMux
    port map (
            O => \N__35799\,
            I => \N__35796\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__35796\,
            I => \N__35793\
        );

    \I__7166\ : Span4Mux_h
    port map (
            O => \N__35793\,
            I => \N__35790\
        );

    \I__7165\ : Odrv4
    port map (
            O => \N__35790\,
            I => \current_shift_inst.un38_control_input_0_s0_20\
        );

    \I__7164\ : InMux
    port map (
            O => \N__35787\,
            I => \current_shift_inst.un38_control_input_cry_19_s0\
        );

    \I__7163\ : InMux
    port map (
            O => \N__35784\,
            I => \current_shift_inst.un38_control_input_cry_2_s0\
        );

    \I__7162\ : InMux
    port map (
            O => \N__35781\,
            I => \current_shift_inst.un38_control_input_cry_3_s0\
        );

    \I__7161\ : InMux
    port map (
            O => \N__35778\,
            I => \N__35775\
        );

    \I__7160\ : LocalMux
    port map (
            O => \N__35775\,
            I => \N__35772\
        );

    \I__7159\ : Span4Mux_h
    port map (
            O => \N__35772\,
            I => \N__35769\
        );

    \I__7158\ : Odrv4
    port map (
            O => \N__35769\,
            I => \current_shift_inst.un38_control_input_0_s0_5\
        );

    \I__7157\ : InMux
    port map (
            O => \N__35766\,
            I => \current_shift_inst.un38_control_input_cry_4_s0\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35763\,
            I => \current_shift_inst.un38_control_input_cry_5_s0\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35760\,
            I => \current_shift_inst.un38_control_input_cry_6_s0\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35757\,
            I => \bfn_14_14_0_\
        );

    \I__7153\ : InMux
    port map (
            O => \N__35754\,
            I => \N__35751\
        );

    \I__7152\ : LocalMux
    port map (
            O => \N__35751\,
            I => \N__35748\
        );

    \I__7151\ : Span4Mux_h
    port map (
            O => \N__35748\,
            I => \N__35745\
        );

    \I__7150\ : Odrv4
    port map (
            O => \N__35745\,
            I => \current_shift_inst.un38_control_input_0_s0_9\
        );

    \I__7149\ : InMux
    port map (
            O => \N__35742\,
            I => \current_shift_inst.un38_control_input_cry_8_s0\
        );

    \I__7148\ : InMux
    port map (
            O => \N__35739\,
            I => \current_shift_inst.un38_control_input_cry_9_s0\
        );

    \I__7147\ : InMux
    port map (
            O => \N__35736\,
            I => \current_shift_inst.un38_control_input_cry_10_s0\
        );

    \I__7146\ : CascadeMux
    port map (
            O => \N__35733\,
            I => \N__35730\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35730\,
            I => \N__35727\
        );

    \I__7144\ : LocalMux
    port map (
            O => \N__35727\,
            I => \N__35724\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__35724\,
            I => \N__35721\
        );

    \I__7142\ : Odrv4
    port map (
            O => \N__35721\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\
        );

    \I__7141\ : InMux
    port map (
            O => \N__35718\,
            I => \N__35714\
        );

    \I__7140\ : InMux
    port map (
            O => \N__35717\,
            I => \N__35711\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__35714\,
            I => \N__35707\
        );

    \I__7138\ : LocalMux
    port map (
            O => \N__35711\,
            I => \N__35702\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35710\,
            I => \N__35699\
        );

    \I__7136\ : Span4Mux_h
    port map (
            O => \N__35707\,
            I => \N__35696\
        );

    \I__7135\ : InMux
    port map (
            O => \N__35706\,
            I => \N__35691\
        );

    \I__7134\ : InMux
    port map (
            O => \N__35705\,
            I => \N__35691\
        );

    \I__7133\ : Span4Mux_v
    port map (
            O => \N__35702\,
            I => \N__35688\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__35699\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7131\ : Odrv4
    port map (
            O => \N__35696\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35691\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7129\ : Odrv4
    port map (
            O => \N__35688\,
            I => \phase_controller_inst2.stoper_tr.start_latchedZ0\
        );

    \I__7128\ : InMux
    port map (
            O => \N__35679\,
            I => \N__35675\
        );

    \I__7127\ : InMux
    port map (
            O => \N__35678\,
            I => \N__35672\
        );

    \I__7126\ : LocalMux
    port map (
            O => \N__35675\,
            I => \N__35669\
        );

    \I__7125\ : LocalMux
    port map (
            O => \N__35672\,
            I => \N__35664\
        );

    \I__7124\ : Span4Mux_v
    port map (
            O => \N__35669\,
            I => \N__35664\
        );

    \I__7123\ : Odrv4
    port map (
            O => \N__35664\,
            I => \phase_controller_inst2.stoper_tr.runningZ0\
        );

    \I__7122\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35657\
        );

    \I__7121\ : InMux
    port map (
            O => \N__35660\,
            I => \N__35652\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__35657\,
            I => \N__35649\
        );

    \I__7119\ : CascadeMux
    port map (
            O => \N__35656\,
            I => \N__35646\
        );

    \I__7118\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35643\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__35652\,
            I => \N__35638\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__35649\,
            I => \N__35638\
        );

    \I__7115\ : InMux
    port map (
            O => \N__35646\,
            I => \N__35635\
        );

    \I__7114\ : LocalMux
    port map (
            O => \N__35643\,
            I => \N__35632\
        );

    \I__7113\ : Span4Mux_v
    port map (
            O => \N__35638\,
            I => \N__35629\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__35635\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7111\ : Odrv4
    port map (
            O => \N__35632\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7110\ : Odrv4
    port map (
            O => \N__35629\,
            I => \phase_controller_inst2.start_timer_trZ0\
        );

    \I__7109\ : InMux
    port map (
            O => \N__35622\,
            I => \N__35613\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35621\,
            I => \N__35613\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35620\,
            I => \N__35606\
        );

    \I__7106\ : InMux
    port map (
            O => \N__35619\,
            I => \N__35606\
        );

    \I__7105\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35606\
        );

    \I__7104\ : LocalMux
    port map (
            O => \N__35613\,
            I => \N__35603\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__35606\,
            I => \N__35600\
        );

    \I__7102\ : Span12Mux_s11_v
    port map (
            O => \N__35603\,
            I => \N__35597\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__35600\,
            I => \N__35594\
        );

    \I__7100\ : Odrv12
    port map (
            O => \N__35597\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7099\ : Odrv4
    port map (
            O => \N__35594\,
            I => \phase_controller_inst2.stoper_tr.un2_start_0\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35589\,
            I => \N__35586\
        );

    \I__7097\ : LocalMux
    port map (
            O => \N__35586\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\
        );

    \I__7096\ : CascadeMux
    port map (
            O => \N__35583\,
            I => \N__35578\
        );

    \I__7095\ : InMux
    port map (
            O => \N__35582\,
            I => \N__35575\
        );

    \I__7094\ : InMux
    port map (
            O => \N__35581\,
            I => \N__35570\
        );

    \I__7093\ : InMux
    port map (
            O => \N__35578\,
            I => \N__35570\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__35575\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7091\ : LocalMux
    port map (
            O => \N__35570\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\
        );

    \I__7090\ : InMux
    port map (
            O => \N__35565\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\
        );

    \I__7089\ : InMux
    port map (
            O => \N__35562\,
            I => \N__35555\
        );

    \I__7088\ : InMux
    port map (
            O => \N__35561\,
            I => \N__35555\
        );

    \I__7087\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35552\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35555\,
            I => \N__35549\
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35552\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__7084\ : Odrv4
    port map (
            O => \N__35549\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\
        );

    \I__7083\ : InMux
    port map (
            O => \N__35544\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\
        );

    \I__7082\ : InMux
    port map (
            O => \N__35541\,
            I => \N__35534\
        );

    \I__7081\ : InMux
    port map (
            O => \N__35540\,
            I => \N__35534\
        );

    \I__7080\ : InMux
    port map (
            O => \N__35539\,
            I => \N__35531\
        );

    \I__7079\ : LocalMux
    port map (
            O => \N__35534\,
            I => \N__35528\
        );

    \I__7078\ : LocalMux
    port map (
            O => \N__35531\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__7077\ : Odrv4
    port map (
            O => \N__35528\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\
        );

    \I__7076\ : InMux
    port map (
            O => \N__35523\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\
        );

    \I__7075\ : CascadeMux
    port map (
            O => \N__35520\,
            I => \N__35516\
        );

    \I__7074\ : CascadeMux
    port map (
            O => \N__35519\,
            I => \N__35513\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35516\,
            I => \N__35510\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35513\,
            I => \N__35507\
        );

    \I__7071\ : LocalMux
    port map (
            O => \N__35510\,
            I => \N__35503\
        );

    \I__7070\ : LocalMux
    port map (
            O => \N__35507\,
            I => \N__35500\
        );

    \I__7069\ : InMux
    port map (
            O => \N__35506\,
            I => \N__35497\
        );

    \I__7068\ : Span4Mux_v
    port map (
            O => \N__35503\,
            I => \N__35494\
        );

    \I__7067\ : Span4Mux_v
    port map (
            O => \N__35500\,
            I => \N__35491\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35497\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7065\ : Odrv4
    port map (
            O => \N__35494\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7064\ : Odrv4
    port map (
            O => \N__35491\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\
        );

    \I__7063\ : InMux
    port map (
            O => \N__35484\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35481\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\
        );

    \I__7061\ : InMux
    port map (
            O => \N__35478\,
            I => \N__35474\
        );

    \I__7060\ : InMux
    port map (
            O => \N__35477\,
            I => \N__35471\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__35474\,
            I => \N__35467\
        );

    \I__7058\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35464\
        );

    \I__7057\ : InMux
    port map (
            O => \N__35470\,
            I => \N__35461\
        );

    \I__7056\ : Span4Mux_v
    port map (
            O => \N__35467\,
            I => \N__35458\
        );

    \I__7055\ : Span4Mux_v
    port map (
            O => \N__35464\,
            I => \N__35455\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__35461\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__35458\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__7052\ : Odrv4
    port map (
            O => \N__35455\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\
        );

    \I__7051\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35445\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__35445\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\
        );

    \I__7049\ : CascadeMux
    port map (
            O => \N__35442\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\
        );

    \I__7048\ : InMux
    port map (
            O => \N__35439\,
            I => \N__35436\
        );

    \I__7047\ : LocalMux
    port map (
            O => \N__35436\,
            I => \N__35433\
        );

    \I__7046\ : Span4Mux_v
    port map (
            O => \N__35433\,
            I => \N__35430\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__35430\,
            I => \N__35427\
        );

    \I__7044\ : Odrv4
    port map (
            O => \N__35427\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\
        );

    \I__7043\ : CascadeMux
    port map (
            O => \N__35424\,
            I => \N__35421\
        );

    \I__7042\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35418\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__35418\,
            I => \N__35415\
        );

    \I__7040\ : Odrv4
    port map (
            O => \N__35415\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35412\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35409\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35406\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35403\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\
        );

    \I__7035\ : InMux
    port map (
            O => \N__35400\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\
        );

    \I__7034\ : InMux
    port map (
            O => \N__35397\,
            I => \N__35390\
        );

    \I__7033\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35390\
        );

    \I__7032\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35387\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__35390\,
            I => \N__35384\
        );

    \I__7030\ : LocalMux
    port map (
            O => \N__35387\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7029\ : Odrv12
    port map (
            O => \N__35384\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\
        );

    \I__7028\ : InMux
    port map (
            O => \N__35379\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\
        );

    \I__7027\ : CascadeMux
    port map (
            O => \N__35376\,
            I => \N__35372\
        );

    \I__7026\ : InMux
    port map (
            O => \N__35375\,
            I => \N__35366\
        );

    \I__7025\ : InMux
    port map (
            O => \N__35372\,
            I => \N__35366\
        );

    \I__7024\ : InMux
    port map (
            O => \N__35371\,
            I => \N__35363\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__35366\,
            I => \N__35360\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__35363\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7021\ : Odrv12
    port map (
            O => \N__35360\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35355\,
            I => \bfn_14_10_0_\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35352\,
            I => \N__35347\
        );

    \I__7018\ : InMux
    port map (
            O => \N__35351\,
            I => \N__35342\
        );

    \I__7017\ : InMux
    port map (
            O => \N__35350\,
            I => \N__35342\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__35347\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7015\ : LocalMux
    port map (
            O => \N__35342\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\
        );

    \I__7014\ : InMux
    port map (
            O => \N__35337\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\
        );

    \I__7013\ : InMux
    port map (
            O => \N__35334\,
            I => \N__35330\
        );

    \I__7012\ : InMux
    port map (
            O => \N__35333\,
            I => \N__35327\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35330\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__35327\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\
        );

    \I__7009\ : InMux
    port map (
            O => \N__35322\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\
        );

    \I__7008\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35315\
        );

    \I__7007\ : InMux
    port map (
            O => \N__35318\,
            I => \N__35312\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__35315\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__35312\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\
        );

    \I__7004\ : InMux
    port map (
            O => \N__35307\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\
        );

    \I__7003\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35300\
        );

    \I__7002\ : InMux
    port map (
            O => \N__35303\,
            I => \N__35297\
        );

    \I__7001\ : LocalMux
    port map (
            O => \N__35300\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__35297\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\
        );

    \I__6999\ : InMux
    port map (
            O => \N__35292\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\
        );

    \I__6998\ : InMux
    port map (
            O => \N__35289\,
            I => \N__35285\
        );

    \I__6997\ : InMux
    port map (
            O => \N__35288\,
            I => \N__35282\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__35285\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__35282\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\
        );

    \I__6994\ : InMux
    port map (
            O => \N__35277\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\
        );

    \I__6993\ : InMux
    port map (
            O => \N__35274\,
            I => \N__35270\
        );

    \I__6992\ : InMux
    port map (
            O => \N__35273\,
            I => \N__35267\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__35270\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6990\ : LocalMux
    port map (
            O => \N__35267\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\
        );

    \I__6989\ : InMux
    port map (
            O => \N__35262\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\
        );

    \I__6988\ : InMux
    port map (
            O => \N__35259\,
            I => \N__35255\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35258\,
            I => \N__35252\
        );

    \I__6986\ : LocalMux
    port map (
            O => \N__35255\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__35252\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\
        );

    \I__6984\ : InMux
    port map (
            O => \N__35247\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35244\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\
        );

    \I__6982\ : InMux
    port map (
            O => \N__35241\,
            I => \bfn_14_9_0_\
        );

    \I__6981\ : InMux
    port map (
            O => \N__35238\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\
        );

    \I__6980\ : InMux
    port map (
            O => \N__35235\,
            I => \N__35231\
        );

    \I__6979\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35228\
        );

    \I__6978\ : LocalMux
    port map (
            O => \N__35231\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6977\ : LocalMux
    port map (
            O => \N__35228\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\
        );

    \I__6976\ : InMux
    port map (
            O => \N__35223\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\
        );

    \I__6975\ : CascadeMux
    port map (
            O => \N__35220\,
            I => \N__35217\
        );

    \I__6974\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35214\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__35214\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\
        );

    \I__6972\ : InMux
    port map (
            O => \N__35211\,
            I => \N__35207\
        );

    \I__6971\ : InMux
    port map (
            O => \N__35210\,
            I => \N__35204\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35207\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6969\ : LocalMux
    port map (
            O => \N__35204\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\
        );

    \I__6968\ : InMux
    port map (
            O => \N__35199\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\
        );

    \I__6967\ : InMux
    port map (
            O => \N__35196\,
            I => \N__35192\
        );

    \I__6966\ : InMux
    port map (
            O => \N__35195\,
            I => \N__35189\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__35192\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6964\ : LocalMux
    port map (
            O => \N__35189\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\
        );

    \I__6963\ : InMux
    port map (
            O => \N__35184\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\
        );

    \I__6962\ : InMux
    port map (
            O => \N__35181\,
            I => \N__35177\
        );

    \I__6961\ : InMux
    port map (
            O => \N__35180\,
            I => \N__35174\
        );

    \I__6960\ : LocalMux
    port map (
            O => \N__35177\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__35174\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\
        );

    \I__6958\ : InMux
    port map (
            O => \N__35169\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\
        );

    \I__6957\ : InMux
    port map (
            O => \N__35166\,
            I => \N__35162\
        );

    \I__6956\ : InMux
    port map (
            O => \N__35165\,
            I => \N__35159\
        );

    \I__6955\ : LocalMux
    port map (
            O => \N__35162\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6954\ : LocalMux
    port map (
            O => \N__35159\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\
        );

    \I__6953\ : InMux
    port map (
            O => \N__35154\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\
        );

    \I__6952\ : InMux
    port map (
            O => \N__35151\,
            I => \N__35147\
        );

    \I__6951\ : InMux
    port map (
            O => \N__35150\,
            I => \N__35144\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35147\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6949\ : LocalMux
    port map (
            O => \N__35144\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\
        );

    \I__6948\ : InMux
    port map (
            O => \N__35139\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\
        );

    \I__6947\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35132\
        );

    \I__6946\ : InMux
    port map (
            O => \N__35135\,
            I => \N__35129\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__35132\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__35129\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\
        );

    \I__6943\ : InMux
    port map (
            O => \N__35124\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\
        );

    \I__6942\ : InMux
    port map (
            O => \N__35121\,
            I => \N__35117\
        );

    \I__6941\ : InMux
    port map (
            O => \N__35120\,
            I => \N__35114\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__35117\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6939\ : LocalMux
    port map (
            O => \N__35114\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\
        );

    \I__6938\ : InMux
    port map (
            O => \N__35109\,
            I => \bfn_14_8_0_\
        );

    \I__6937\ : InMux
    port map (
            O => \N__35106\,
            I => \N__35102\
        );

    \I__6936\ : InMux
    port map (
            O => \N__35105\,
            I => \N__35099\
        );

    \I__6935\ : LocalMux
    port map (
            O => \N__35102\,
            I => \N__35094\
        );

    \I__6934\ : LocalMux
    port map (
            O => \N__35099\,
            I => \N__35094\
        );

    \I__6933\ : Span4Mux_s3_v
    port map (
            O => \N__35094\,
            I => \N__35091\
        );

    \I__6932\ : Span4Mux_h
    port map (
            O => \N__35091\,
            I => \N__35088\
        );

    \I__6931\ : Sp12to4
    port map (
            O => \N__35088\,
            I => \N__35079\
        );

    \I__6930\ : InMux
    port map (
            O => \N__35087\,
            I => \N__35076\
        );

    \I__6929\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35071\
        );

    \I__6928\ : InMux
    port map (
            O => \N__35085\,
            I => \N__35071\
        );

    \I__6927\ : InMux
    port map (
            O => \N__35084\,
            I => \N__35064\
        );

    \I__6926\ : InMux
    port map (
            O => \N__35083\,
            I => \N__35064\
        );

    \I__6925\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35064\
        );

    \I__6924\ : Span12Mux_v
    port map (
            O => \N__35079\,
            I => \N__35061\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35054\
        );

    \I__6922\ : LocalMux
    port map (
            O => \N__35071\,
            I => \N__35054\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__35054\
        );

    \I__6920\ : Span12Mux_v
    port map (
            O => \N__35061\,
            I => \N__35051\
        );

    \I__6919\ : Span4Mux_v
    port map (
            O => \N__35054\,
            I => \N__35048\
        );

    \I__6918\ : Span12Mux_h
    port map (
            O => \N__35051\,
            I => \N__35045\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__35048\,
            I => \N__35042\
        );

    \I__6916\ : Odrv12
    port map (
            O => \N__35045\,
            I => start_stop_c
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__35042\,
            I => start_stop_c
        );

    \I__6914\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35032\
        );

    \I__6913\ : InMux
    port map (
            O => \N__35036\,
            I => \N__35027\
        );

    \I__6912\ : InMux
    port map (
            O => \N__35035\,
            I => \N__35027\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__35032\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__35027\,
            I => \phase_controller_inst2.stateZ0Z_4\
        );

    \I__6909\ : CascadeMux
    port map (
            O => \N__35022\,
            I => \N__35018\
        );

    \I__6908\ : InMux
    port map (
            O => \N__35021\,
            I => \N__35014\
        );

    \I__6907\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35009\
        );

    \I__6906\ : InMux
    port map (
            O => \N__35017\,
            I => \N__35009\
        );

    \I__6905\ : LocalMux
    port map (
            O => \N__35014\,
            I => \phase_controller_inst2.start_flagZ0\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__35009\,
            I => \phase_controller_inst2.start_flagZ0\
        );

    \I__6903\ : CascadeMux
    port map (
            O => \N__35004\,
            I => \N__35001\
        );

    \I__6902\ : InMux
    port map (
            O => \N__35001\,
            I => \N__34998\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__34998\,
            I => \N__34995\
        );

    \I__6900\ : Span4Mux_v
    port map (
            O => \N__34995\,
            I => \N__34992\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__34992\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt24\
        );

    \I__6898\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34986\
        );

    \I__6897\ : LocalMux
    port map (
            O => \N__34986\,
            I => \N__34983\
        );

    \I__6896\ : Span4Mux_v
    port map (
            O => \N__34983\,
            I => \N__34980\
        );

    \I__6895\ : Odrv4
    port map (
            O => \N__34980\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\
        );

    \I__6894\ : CascadeMux
    port map (
            O => \N__34977\,
            I => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\
        );

    \I__6893\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34971\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__34971\,
            I => \N__34968\
        );

    \I__6891\ : Odrv4
    port map (
            O => \N__34968\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\
        );

    \I__6890\ : CascadeMux
    port map (
            O => \N__34965\,
            I => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\
        );

    \I__6889\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34956\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34961\,
            I => \N__34956\
        );

    \I__6887\ : LocalMux
    port map (
            O => \N__34956\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\
        );

    \I__6886\ : InMux
    port map (
            O => \N__34953\,
            I => \N__34950\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__34950\,
            I => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\
        );

    \I__6884\ : CascadeMux
    port map (
            O => \N__34947\,
            I => \N__34943\
        );

    \I__6883\ : InMux
    port map (
            O => \N__34946\,
            I => \N__34939\
        );

    \I__6882\ : InMux
    port map (
            O => \N__34943\,
            I => \N__34936\
        );

    \I__6881\ : InMux
    port map (
            O => \N__34942\,
            I => \N__34933\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__34939\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6879\ : LocalMux
    port map (
            O => \N__34936\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6878\ : LocalMux
    port map (
            O => \N__34933\,
            I => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\
        );

    \I__6877\ : IoInMux
    port map (
            O => \N__34926\,
            I => \N__34923\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__6875\ : Odrv12
    port map (
            O => \N__34920\,
            I => s2_phy_c
        );

    \I__6874\ : CascadeMux
    port map (
            O => \N__34917\,
            I => \N__34911\
        );

    \I__6873\ : CascadeMux
    port map (
            O => \N__34916\,
            I => \N__34907\
        );

    \I__6872\ : InMux
    port map (
            O => \N__34915\,
            I => \N__34902\
        );

    \I__6871\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34902\
        );

    \I__6870\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34899\
        );

    \I__6869\ : CascadeMux
    port map (
            O => \N__34910\,
            I => \N__34896\
        );

    \I__6868\ : InMux
    port map (
            O => \N__34907\,
            I => \N__34893\
        );

    \I__6867\ : LocalMux
    port map (
            O => \N__34902\,
            I => \N__34888\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__34899\,
            I => \N__34888\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34896\,
            I => \N__34884\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__34893\,
            I => \N__34879\
        );

    \I__6863\ : Span12Mux_v
    port map (
            O => \N__34888\,
            I => \N__34879\
        );

    \I__6862\ : InMux
    port map (
            O => \N__34887\,
            I => \N__34876\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34884\,
            I => state_3
        );

    \I__6860\ : Odrv12
    port map (
            O => \N__34879\,
            I => state_3
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__34876\,
            I => state_3
        );

    \I__6858\ : IoInMux
    port map (
            O => \N__34869\,
            I => \N__34866\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__34866\,
            I => \N__34863\
        );

    \I__6856\ : Span4Mux_s0_v
    port map (
            O => \N__34863\,
            I => \N__34860\
        );

    \I__6855\ : Span4Mux_v
    port map (
            O => \N__34860\,
            I => \N__34857\
        );

    \I__6854\ : Span4Mux_v
    port map (
            O => \N__34857\,
            I => \N__34852\
        );

    \I__6853\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34849\
        );

    \I__6852\ : InMux
    port map (
            O => \N__34855\,
            I => \N__34846\
        );

    \I__6851\ : Odrv4
    port map (
            O => \N__34852\,
            I => s1_phy_c
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__34849\,
            I => s1_phy_c
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__34846\,
            I => s1_phy_c
        );

    \I__6848\ : InMux
    port map (
            O => \N__34839\,
            I => \N__34833\
        );

    \I__6847\ : InMux
    port map (
            O => \N__34838\,
            I => \N__34828\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34837\,
            I => \N__34828\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34836\,
            I => \N__34825\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__34833\,
            I => \N__34822\
        );

    \I__6843\ : LocalMux
    port map (
            O => \N__34828\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__34825\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6841\ : Odrv4
    port map (
            O => \N__34822\,
            I => \current_shift_inst.start_timer_sZ0Z1\
        );

    \I__6840\ : InMux
    port map (
            O => \N__34815\,
            I => \N__34807\
        );

    \I__6839\ : InMux
    port map (
            O => \N__34814\,
            I => \N__34807\
        );

    \I__6838\ : InMux
    port map (
            O => \N__34813\,
            I => \N__34804\
        );

    \I__6837\ : InMux
    port map (
            O => \N__34812\,
            I => \N__34801\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34807\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34804\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__34801\,
            I => \current_shift_inst.stop_timer_sZ0Z1\
        );

    \I__6833\ : IoInMux
    port map (
            O => \N__34794\,
            I => \N__34791\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__34791\,
            I => \N__34788\
        );

    \I__6831\ : Span4Mux_s3_v
    port map (
            O => \N__34788\,
            I => \N__34785\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__34785\,
            I => \current_shift_inst.timer_s1.N_161_i\
        );

    \I__6829\ : InMux
    port map (
            O => \N__34782\,
            I => \N__34779\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__34779\,
            I => \N__34774\
        );

    \I__6827\ : InMux
    port map (
            O => \N__34778\,
            I => \N__34771\
        );

    \I__6826\ : InMux
    port map (
            O => \N__34777\,
            I => \N__34768\
        );

    \I__6825\ : IoSpan4Mux
    port map (
            O => \N__34774\,
            I => \N__34765\
        );

    \I__6824\ : LocalMux
    port map (
            O => \N__34771\,
            I => \N__34762\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__34768\,
            I => \N__34759\
        );

    \I__6822\ : IoSpan4Mux
    port map (
            O => \N__34765\,
            I => \N__34756\
        );

    \I__6821\ : IoSpan4Mux
    port map (
            O => \N__34762\,
            I => \N__34751\
        );

    \I__6820\ : IoSpan4Mux
    port map (
            O => \N__34759\,
            I => \N__34751\
        );

    \I__6819\ : Odrv4
    port map (
            O => \N__34756\,
            I => il_min_comp1_c
        );

    \I__6818\ : Odrv4
    port map (
            O => \N__34751\,
            I => il_min_comp1_c
        );

    \I__6817\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34742\
        );

    \I__6816\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34739\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__34742\,
            I => \phase_controller_inst1.N_61\
        );

    \I__6814\ : LocalMux
    port map (
            O => \N__34739\,
            I => \phase_controller_inst1.N_61\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__34731\,
            I => \N__34728\
        );

    \I__6811\ : Sp12to4
    port map (
            O => \N__34728\,
            I => \N__34723\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34727\,
            I => \N__34719\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34726\,
            I => \N__34716\
        );

    \I__6808\ : Span12Mux_v
    port map (
            O => \N__34723\,
            I => \N__34713\
        );

    \I__6807\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34710\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34719\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__34716\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6804\ : Odrv12
    port map (
            O => \N__34713\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6803\ : LocalMux
    port map (
            O => \N__34710\,
            I => \phase_controller_inst1.stateZ0Z_1\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34701\,
            I => \bfn_13_19_0_\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34698\,
            I => \current_shift_inst.un38_control_input_cry_24_s1\
        );

    \I__6800\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34692\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__34692\,
            I => \N__34689\
        );

    \I__6798\ : Odrv4
    port map (
            O => \N__34689\,
            I => \current_shift_inst.un38_control_input_0_s1_26\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34686\,
            I => \current_shift_inst.un38_control_input_cry_25_s1\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34683\,
            I => \N__34680\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__6794\ : Odrv4
    port map (
            O => \N__34677\,
            I => \current_shift_inst.un38_control_input_0_s1_27\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34674\,
            I => \current_shift_inst.un38_control_input_cry_26_s1\
        );

    \I__6792\ : InMux
    port map (
            O => \N__34671\,
            I => \N__34668\
        );

    \I__6791\ : LocalMux
    port map (
            O => \N__34668\,
            I => \N__34665\
        );

    \I__6790\ : Odrv4
    port map (
            O => \N__34665\,
            I => \current_shift_inst.un38_control_input_0_s1_28\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34662\,
            I => \current_shift_inst.un38_control_input_cry_27_s1\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34659\,
            I => \N__34656\
        );

    \I__6787\ : LocalMux
    port map (
            O => \N__34656\,
            I => \N__34653\
        );

    \I__6786\ : Span4Mux_h
    port map (
            O => \N__34653\,
            I => \N__34650\
        );

    \I__6785\ : Odrv4
    port map (
            O => \N__34650\,
            I => \current_shift_inst.un38_control_input_0_s1_29\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34647\,
            I => \current_shift_inst.un38_control_input_cry_28_s1\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34644\,
            I => \N__34641\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__34641\,
            I => \N__34638\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__34638\,
            I => \N__34635\
        );

    \I__6780\ : Odrv4
    port map (
            O => \N__34635\,
            I => \current_shift_inst.un38_control_input_0_s1_30\
        );

    \I__6779\ : InMux
    port map (
            O => \N__34632\,
            I => \current_shift_inst.un38_control_input_cry_29_s1\
        );

    \I__6778\ : InMux
    port map (
            O => \N__34629\,
            I => \current_shift_inst.un38_control_input_cry_30_s1\
        );

    \I__6777\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34623\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__34623\,
            I => \N__34620\
        );

    \I__6775\ : Odrv4
    port map (
            O => \N__34620\,
            I => \current_shift_inst.un38_control_input_0_s1_15\
        );

    \I__6774\ : InMux
    port map (
            O => \N__34617\,
            I => \current_shift_inst.un38_control_input_cry_14_s1\
        );

    \I__6773\ : InMux
    port map (
            O => \N__34614\,
            I => \N__34611\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__34611\,
            I => \N__34608\
        );

    \I__6771\ : Odrv4
    port map (
            O => \N__34608\,
            I => \current_shift_inst.un38_control_input_0_s1_16\
        );

    \I__6770\ : InMux
    port map (
            O => \N__34605\,
            I => \bfn_13_18_0_\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34602\,
            I => \N__34599\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__34599\,
            I => \N__34596\
        );

    \I__6767\ : Odrv4
    port map (
            O => \N__34596\,
            I => \current_shift_inst.un38_control_input_0_s1_17\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34593\,
            I => \current_shift_inst.un38_control_input_cry_16_s1\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34587\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__34587\,
            I => \N__34584\
        );

    \I__6763\ : Odrv4
    port map (
            O => \N__34584\,
            I => \current_shift_inst.un38_control_input_0_s1_18\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34581\,
            I => \current_shift_inst.un38_control_input_cry_17_s1\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34578\,
            I => \N__34575\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34572\
        );

    \I__6759\ : Odrv4
    port map (
            O => \N__34572\,
            I => \current_shift_inst.un38_control_input_0_s1_19\
        );

    \I__6758\ : InMux
    port map (
            O => \N__34569\,
            I => \current_shift_inst.un38_control_input_cry_18_s1\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34563\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__34563\,
            I => \N__34560\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__34560\,
            I => \current_shift_inst.un38_control_input_0_s1_20\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34557\,
            I => \current_shift_inst.un38_control_input_cry_19_s1\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34554\,
            I => \N__34551\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__34551\,
            I => \N__34548\
        );

    \I__6751\ : Odrv4
    port map (
            O => \N__34548\,
            I => \current_shift_inst.un38_control_input_0_s1_21\
        );

    \I__6750\ : InMux
    port map (
            O => \N__34545\,
            I => \current_shift_inst.un38_control_input_cry_20_s1\
        );

    \I__6749\ : InMux
    port map (
            O => \N__34542\,
            I => \N__34539\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34539\,
            I => \N__34536\
        );

    \I__6747\ : Odrv4
    port map (
            O => \N__34536\,
            I => \current_shift_inst.un38_control_input_0_s1_22\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34533\,
            I => \current_shift_inst.un38_control_input_cry_21_s1\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34530\,
            I => \N__34527\
        );

    \I__6744\ : LocalMux
    port map (
            O => \N__34527\,
            I => \N__34524\
        );

    \I__6743\ : Odrv4
    port map (
            O => \N__34524\,
            I => \current_shift_inst.un38_control_input_0_s1_23\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34521\,
            I => \current_shift_inst.un38_control_input_cry_22_s1\
        );

    \I__6741\ : InMux
    port map (
            O => \N__34518\,
            I => \current_shift_inst.un38_control_input_cry_6_s1\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34515\,
            I => \bfn_13_17_0_\
        );

    \I__6739\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34509\
        );

    \I__6738\ : LocalMux
    port map (
            O => \N__34509\,
            I => \N__34506\
        );

    \I__6737\ : Span4Mux_v
    port map (
            O => \N__34506\,
            I => \N__34503\
        );

    \I__6736\ : Odrv4
    port map (
            O => \N__34503\,
            I => \current_shift_inst.un38_control_input_0_s1_9\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34500\,
            I => \current_shift_inst.un38_control_input_cry_8_s1\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34497\,
            I => \current_shift_inst.un38_control_input_cry_9_s1\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34494\,
            I => \current_shift_inst.un38_control_input_cry_10_s1\
        );

    \I__6732\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34488\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__34488\,
            I => \N__34485\
        );

    \I__6730\ : Odrv4
    port map (
            O => \N__34485\,
            I => \current_shift_inst.un38_control_input_0_s1_12\
        );

    \I__6729\ : InMux
    port map (
            O => \N__34482\,
            I => \current_shift_inst.un38_control_input_cry_11_s1\
        );

    \I__6728\ : InMux
    port map (
            O => \N__34479\,
            I => \N__34476\
        );

    \I__6727\ : LocalMux
    port map (
            O => \N__34476\,
            I => \current_shift_inst.un38_control_input_0_s1_13\
        );

    \I__6726\ : InMux
    port map (
            O => \N__34473\,
            I => \current_shift_inst.un38_control_input_cry_12_s1\
        );

    \I__6725\ : InMux
    port map (
            O => \N__34470\,
            I => \N__34467\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__34467\,
            I => \N__34464\
        );

    \I__6723\ : Odrv4
    port map (
            O => \N__34464\,
            I => \current_shift_inst.un38_control_input_0_s1_14\
        );

    \I__6722\ : InMux
    port map (
            O => \N__34461\,
            I => \current_shift_inst.un38_control_input_cry_13_s1\
        );

    \I__6721\ : CascadeMux
    port map (
            O => \N__34458\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\
        );

    \I__6720\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34450\
        );

    \I__6719\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34447\
        );

    \I__6718\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34444\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__34450\,
            I => \N__34439\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__34447\,
            I => \N__34439\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__34444\,
            I => \N__34436\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__34439\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__6713\ : Odrv4
    port map (
            O => \N__34436\,
            I => \elapsed_time_ns_1_RNI04EN9_0_31\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34431\,
            I => \N__34427\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34430\,
            I => \N__34424\
        );

    \I__6710\ : LocalMux
    port map (
            O => \N__34427\,
            I => \N__34421\
        );

    \I__6709\ : LocalMux
    port map (
            O => \N__34424\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__6708\ : Odrv4
    port map (
            O => \N__34421\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34416\,
            I => \N__34412\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34415\,
            I => \N__34409\
        );

    \I__6705\ : LocalMux
    port map (
            O => \N__34412\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__6704\ : LocalMux
    port map (
            O => \N__34409\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__34404\,
            I => \N__34401\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34401\,
            I => \N__34398\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__34398\,
            I => \N__34395\
        );

    \I__6700\ : Span4Mux_v
    port map (
            O => \N__34395\,
            I => \N__34392\
        );

    \I__6699\ : Odrv4
    port map (
            O => \N__34392\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34389\,
            I => \current_shift_inst.un38_control_input_cry_2_s1\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34386\,
            I => \current_shift_inst.un38_control_input_cry_3_s1\
        );

    \I__6696\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34380\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__34380\,
            I => \N__34377\
        );

    \I__6694\ : Span4Mux_h
    port map (
            O => \N__34377\,
            I => \N__34374\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__34374\,
            I => \current_shift_inst.un38_control_input_0_s1_5\
        );

    \I__6692\ : InMux
    port map (
            O => \N__34371\,
            I => \current_shift_inst.un38_control_input_cry_4_s1\
        );

    \I__6691\ : InMux
    port map (
            O => \N__34368\,
            I => \current_shift_inst.un38_control_input_cry_5_s1\
        );

    \I__6690\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34362\
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__34362\,
            I => \N__34359\
        );

    \I__6688\ : Odrv12
    port map (
            O => \N__34359\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\
        );

    \I__6687\ : InMux
    port map (
            O => \N__34356\,
            I => \N__34353\
        );

    \I__6686\ : LocalMux
    port map (
            O => \N__34353\,
            I => \N__34350\
        );

    \I__6685\ : Odrv12
    port map (
            O => \N__34350\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34347\,
            I => \N__34342\
        );

    \I__6683\ : InMux
    port map (
            O => \N__34346\,
            I => \N__34339\
        );

    \I__6682\ : InMux
    port map (
            O => \N__34345\,
            I => \N__34336\
        );

    \I__6681\ : LocalMux
    port map (
            O => \N__34342\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__34339\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__6679\ : LocalMux
    port map (
            O => \N__34336\,
            I => \elapsed_time_ns_1_RNIV2EN9_0_30\
        );

    \I__6678\ : InMux
    port map (
            O => \N__34329\,
            I => \N__34326\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__34326\,
            I => \N__34323\
        );

    \I__6676\ : Odrv12
    port map (
            O => \N__34323\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\
        );

    \I__6675\ : CascadeMux
    port map (
            O => \N__34320\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34317\,
            I => \N__34314\
        );

    \I__6673\ : LocalMux
    port map (
            O => \N__34314\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\
        );

    \I__6672\ : CascadeMux
    port map (
            O => \N__34311\,
            I => \N__34308\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34308\,
            I => \N__34305\
        );

    \I__6670\ : LocalMux
    port map (
            O => \N__34305\,
            I => \N__34302\
        );

    \I__6669\ : Odrv12
    port map (
            O => \N__34302\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34296\
        );

    \I__6667\ : LocalMux
    port map (
            O => \N__34296\,
            I => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\
        );

    \I__6666\ : CascadeMux
    port map (
            O => \N__34293\,
            I => \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34284\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34284\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__34284\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__34281\,
            I => \N__34278\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34278\,
            I => \N__34275\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__34275\,
            I => \N__34272\
        );

    \I__6659\ : Odrv4
    port map (
            O => \N__34272\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt28\
        );

    \I__6658\ : InMux
    port map (
            O => \N__34269\,
            I => \N__34266\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__34266\,
            I => \N__34262\
        );

    \I__6656\ : InMux
    port map (
            O => \N__34265\,
            I => \N__34259\
        );

    \I__6655\ : Odrv4
    port map (
            O => \N__34262\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__34259\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28\
        );

    \I__6653\ : CascadeMux
    port map (
            O => \N__34254\,
            I => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\
        );

    \I__6652\ : InMux
    port map (
            O => \N__34251\,
            I => \N__34247\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34250\,
            I => \N__34243\
        );

    \I__6650\ : LocalMux
    port map (
            O => \N__34247\,
            I => \N__34240\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34246\,
            I => \N__34237\
        );

    \I__6648\ : LocalMux
    port map (
            O => \N__34243\,
            I => \N__34234\
        );

    \I__6647\ : Span4Mux_h
    port map (
            O => \N__34240\,
            I => \N__34231\
        );

    \I__6646\ : LocalMux
    port map (
            O => \N__34237\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6645\ : Odrv12
    port map (
            O => \N__34234\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6644\ : Odrv4
    port map (
            O => \N__34231\,
            I => \elapsed_time_ns_1_RNI7ADN9_0_29\
        );

    \I__6643\ : CascadeMux
    port map (
            O => \N__34224\,
            I => \N__34220\
        );

    \I__6642\ : CascadeMux
    port map (
            O => \N__34223\,
            I => \N__34217\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34220\,
            I => \N__34212\
        );

    \I__6640\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34212\
        );

    \I__6639\ : LocalMux
    port map (
            O => \N__34212\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34209\,
            I => \N__34203\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34208\,
            I => \N__34203\
        );

    \I__6636\ : LocalMux
    port map (
            O => \N__34203\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34200\,
            I => \N__34197\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__6633\ : Odrv4
    port map (
            O => \N__34194\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\
        );

    \I__6632\ : InMux
    port map (
            O => \N__34191\,
            I => \N__34188\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__34188\,
            I => \N__34185\
        );

    \I__6630\ : Odrv12
    port map (
            O => \N__34185\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\
        );

    \I__6629\ : InMux
    port map (
            O => \N__34182\,
            I => \N__34179\
        );

    \I__6628\ : LocalMux
    port map (
            O => \N__34179\,
            I => \N__34176\
        );

    \I__6627\ : Span4Mux_h
    port map (
            O => \N__34176\,
            I => \N__34173\
        );

    \I__6626\ : Odrv4
    port map (
            O => \N__34173\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34167\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__34167\,
            I => \N__34164\
        );

    \I__6623\ : Span4Mux_h
    port map (
            O => \N__34164\,
            I => \N__34161\
        );

    \I__6622\ : Odrv4
    port map (
            O => \N__34161\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\
        );

    \I__6621\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34155\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__34155\,
            I => \N__34152\
        );

    \I__6619\ : Span4Mux_h
    port map (
            O => \N__34152\,
            I => \N__34149\
        );

    \I__6618\ : Odrv4
    port map (
            O => \N__34149\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt30\
        );

    \I__6617\ : InMux
    port map (
            O => \N__34146\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30\
        );

    \I__6616\ : CascadeMux
    port map (
            O => \N__34143\,
            I => \N__34139\
        );

    \I__6615\ : InMux
    port map (
            O => \N__34142\,
            I => \N__34135\
        );

    \I__6614\ : InMux
    port map (
            O => \N__34139\,
            I => \N__34130\
        );

    \I__6613\ : InMux
    port map (
            O => \N__34138\,
            I => \N__34130\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__34135\,
            I => \N__34127\
        );

    \I__6611\ : LocalMux
    port map (
            O => \N__34130\,
            I => \N__34124\
        );

    \I__6610\ : Span4Mux_v
    port map (
            O => \N__34127\,
            I => \N__34119\
        );

    \I__6609\ : Span4Mux_h
    port map (
            O => \N__34124\,
            I => \N__34119\
        );

    \I__6608\ : Odrv4
    port map (
            O => \N__34119\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__34116\,
            I => \N__34113\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34110\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__34110\,
            I => \phase_controller_inst1.stoper_hc.un4_running_lt26\
        );

    \I__6604\ : InMux
    port map (
            O => \N__34107\,
            I => \N__34104\
        );

    \I__6603\ : LocalMux
    port map (
            O => \N__34104\,
            I => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\
        );

    \I__6602\ : CascadeMux
    port map (
            O => \N__34101\,
            I => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\
        );

    \I__6601\ : CascadeMux
    port map (
            O => \N__34098\,
            I => \N__34095\
        );

    \I__6600\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34092\
        );

    \I__6599\ : LocalMux
    port map (
            O => \N__34092\,
            I => \N__34089\
        );

    \I__6598\ : Odrv4
    port map (
            O => \N__34089\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__34086\,
            I => \N__34082\
        );

    \I__6596\ : InMux
    port map (
            O => \N__34085\,
            I => \N__34077\
        );

    \I__6595\ : InMux
    port map (
            O => \N__34082\,
            I => \N__34077\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34077\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\
        );

    \I__6593\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34071\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__34071\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\
        );

    \I__6591\ : CascadeMux
    port map (
            O => \N__34068\,
            I => \N__34065\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34065\,
            I => \N__34062\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__34062\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\
        );

    \I__6588\ : CascadeMux
    port map (
            O => \N__34059\,
            I => \N__34056\
        );

    \I__6587\ : InMux
    port map (
            O => \N__34056\,
            I => \N__34053\
        );

    \I__6586\ : LocalMux
    port map (
            O => \N__34053\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\
        );

    \I__6585\ : CascadeMux
    port map (
            O => \N__34050\,
            I => \N__34047\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34047\,
            I => \N__34044\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__34044\,
            I => \N__34041\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__34041\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\
        );

    \I__6581\ : InMux
    port map (
            O => \N__34038\,
            I => \N__34035\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__34035\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\
        );

    \I__6579\ : CascadeMux
    port map (
            O => \N__34032\,
            I => \N__34029\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34029\,
            I => \N__34026\
        );

    \I__6577\ : LocalMux
    port map (
            O => \N__34026\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\
        );

    \I__6576\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34020\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__34020\,
            I => \N__34017\
        );

    \I__6574\ : Span4Mux_v
    port map (
            O => \N__34017\,
            I => \N__34014\
        );

    \I__6573\ : Odrv4
    port map (
            O => \N__34014\,
            I => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\
        );

    \I__6572\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \N__34008\
        );

    \I__6571\ : InMux
    port map (
            O => \N__34008\,
            I => \N__34005\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__6569\ : Odrv4
    port map (
            O => \N__34002\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__33999\,
            I => \N__33996\
        );

    \I__6567\ : InMux
    port map (
            O => \N__33996\,
            I => \N__33993\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__33993\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\
        );

    \I__6565\ : InMux
    port map (
            O => \N__33990\,
            I => \N__33987\
        );

    \I__6564\ : LocalMux
    port map (
            O => \N__33987\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\
        );

    \I__6563\ : CascadeMux
    port map (
            O => \N__33984\,
            I => \N__33981\
        );

    \I__6562\ : InMux
    port map (
            O => \N__33981\,
            I => \N__33978\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__33978\,
            I => \N__33975\
        );

    \I__6560\ : Odrv4
    port map (
            O => \N__33975\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\
        );

    \I__6559\ : CascadeMux
    port map (
            O => \N__33972\,
            I => \N__33969\
        );

    \I__6558\ : InMux
    port map (
            O => \N__33969\,
            I => \N__33966\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__33966\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\
        );

    \I__6556\ : CascadeMux
    port map (
            O => \N__33963\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\
        );

    \I__6555\ : InMux
    port map (
            O => \N__33960\,
            I => \N__33954\
        );

    \I__6554\ : InMux
    port map (
            O => \N__33959\,
            I => \N__33954\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__33954\,
            I => \phase_controller_inst1.stoper_hc.runningZ0\
        );

    \I__6552\ : CascadeMux
    port map (
            O => \N__33951\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\
        );

    \I__6551\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33945\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__33945\,
            I => \N__33939\
        );

    \I__6549\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33932\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33943\,
            I => \N__33932\
        );

    \I__6547\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33932\
        );

    \I__6546\ : Odrv4
    port map (
            O => \N__33939\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6545\ : LocalMux
    port map (
            O => \N__33932\,
            I => \phase_controller_inst1.stoper_hc.un2_start_0\
        );

    \I__6544\ : CascadeMux
    port map (
            O => \N__33927\,
            I => \N__33924\
        );

    \I__6543\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33918\
        );

    \I__6542\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33918\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__33918\,
            I => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\
        );

    \I__6540\ : CascadeMux
    port map (
            O => \N__33915\,
            I => \N__33912\
        );

    \I__6539\ : InMux
    port map (
            O => \N__33912\,
            I => \N__33909\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__33909\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\
        );

    \I__6537\ : CascadeMux
    port map (
            O => \N__33906\,
            I => \N__33903\
        );

    \I__6536\ : InMux
    port map (
            O => \N__33903\,
            I => \N__33900\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__33900\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\
        );

    \I__6534\ : CascadeMux
    port map (
            O => \N__33897\,
            I => \N__33894\
        );

    \I__6533\ : InMux
    port map (
            O => \N__33894\,
            I => \N__33891\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33891\,
            I => \N__33888\
        );

    \I__6531\ : Odrv4
    port map (
            O => \N__33888\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\
        );

    \I__6530\ : CascadeMux
    port map (
            O => \N__33885\,
            I => \N__33882\
        );

    \I__6529\ : InMux
    port map (
            O => \N__33882\,
            I => \N__33879\
        );

    \I__6528\ : LocalMux
    port map (
            O => \N__33879\,
            I => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\
        );

    \I__6527\ : CascadeMux
    port map (
            O => \N__33876\,
            I => \N__33872\
        );

    \I__6526\ : CascadeMux
    port map (
            O => \N__33875\,
            I => \N__33869\
        );

    \I__6525\ : InMux
    port map (
            O => \N__33872\,
            I => \N__33861\
        );

    \I__6524\ : InMux
    port map (
            O => \N__33869\,
            I => \N__33861\
        );

    \I__6523\ : InMux
    port map (
            O => \N__33868\,
            I => \N__33861\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__33861\,
            I => \phase_controller_inst1.start_flagZ0\
        );

    \I__6521\ : CascadeMux
    port map (
            O => \N__33858\,
            I => \N__33853\
        );

    \I__6520\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33850\
        );

    \I__6519\ : InMux
    port map (
            O => \N__33856\,
            I => \N__33845\
        );

    \I__6518\ : InMux
    port map (
            O => \N__33853\,
            I => \N__33845\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__33850\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6516\ : LocalMux
    port map (
            O => \N__33845\,
            I => \phase_controller_inst1.stateZ0Z_2\
        );

    \I__6515\ : InMux
    port map (
            O => \N__33840\,
            I => \N__33837\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__33837\,
            I => \phase_controller_inst1.N_54_0\
        );

    \I__6513\ : InMux
    port map (
            O => \N__33834\,
            I => \N__33830\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33833\,
            I => \N__33825\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__33830\,
            I => \N__33822\
        );

    \I__6510\ : InMux
    port map (
            O => \N__33829\,
            I => \N__33817\
        );

    \I__6509\ : InMux
    port map (
            O => \N__33828\,
            I => \N__33817\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__33825\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6507\ : Odrv4
    port map (
            O => \N__33822\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6506\ : LocalMux
    port map (
            O => \N__33817\,
            I => \phase_controller_inst1.hc_time_passed\
        );

    \I__6505\ : InMux
    port map (
            O => \N__33810\,
            I => \N__33806\
        );

    \I__6504\ : InMux
    port map (
            O => \N__33809\,
            I => \N__33803\
        );

    \I__6503\ : LocalMux
    port map (
            O => \N__33806\,
            I => \N__33799\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__33803\,
            I => \N__33796\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33793\
        );

    \I__6500\ : Span4Mux_h
    port map (
            O => \N__33799\,
            I => \N__33790\
        );

    \I__6499\ : Span4Mux_h
    port map (
            O => \N__33796\,
            I => \N__33787\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33784\
        );

    \I__6497\ : Span4Mux_h
    port map (
            O => \N__33790\,
            I => \N__33781\
        );

    \I__6496\ : Span4Mux_h
    port map (
            O => \N__33787\,
            I => \N__33778\
        );

    \I__6495\ : IoSpan4Mux
    port map (
            O => \N__33784\,
            I => \N__33775\
        );

    \I__6494\ : Odrv4
    port map (
            O => \N__33781\,
            I => il_max_comp1_c
        );

    \I__6493\ : Odrv4
    port map (
            O => \N__33778\,
            I => il_max_comp1_c
        );

    \I__6492\ : Odrv4
    port map (
            O => \N__33775\,
            I => il_max_comp1_c
        );

    \I__6491\ : CascadeMux
    port map (
            O => \N__33768\,
            I => \N__33765\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33765\,
            I => \N__33762\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__33762\,
            I => \phase_controller_inst2.state_ns_0_0_1\
        );

    \I__6488\ : InMux
    port map (
            O => \N__33759\,
            I => \N__33756\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__33756\,
            I => \N__33753\
        );

    \I__6486\ : Sp12to4
    port map (
            O => \N__33753\,
            I => \N__33750\
        );

    \I__6485\ : Span12Mux_v
    port map (
            O => \N__33750\,
            I => \N__33744\
        );

    \I__6484\ : InMux
    port map (
            O => \N__33749\,
            I => \N__33739\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33748\,
            I => \N__33739\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33736\
        );

    \I__6481\ : Odrv12
    port map (
            O => \N__33744\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__33739\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6479\ : LocalMux
    port map (
            O => \N__33736\,
            I => \phase_controller_inst2.stateZ0Z_3\
        );

    \I__6478\ : CascadeMux
    port map (
            O => \N__33729\,
            I => \N__33726\
        );

    \I__6477\ : InMux
    port map (
            O => \N__33726\,
            I => \N__33721\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33725\,
            I => \N__33718\
        );

    \I__6475\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33715\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__33721\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__33718\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__33715\,
            I => \phase_controller_inst2.stateZ0Z_2\
        );

    \I__6471\ : InMux
    port map (
            O => \N__33708\,
            I => \N__33702\
        );

    \I__6470\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33702\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__33702\,
            I => \phase_controller_inst2.N_61\
        );

    \I__6468\ : InMux
    port map (
            O => \N__33699\,
            I => \N__33659\
        );

    \I__6467\ : InMux
    port map (
            O => \N__33698\,
            I => \N__33659\
        );

    \I__6466\ : InMux
    port map (
            O => \N__33697\,
            I => \N__33659\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33659\
        );

    \I__6464\ : InMux
    port map (
            O => \N__33695\,
            I => \N__33650\
        );

    \I__6463\ : InMux
    port map (
            O => \N__33694\,
            I => \N__33650\
        );

    \I__6462\ : InMux
    port map (
            O => \N__33693\,
            I => \N__33650\
        );

    \I__6461\ : InMux
    port map (
            O => \N__33692\,
            I => \N__33650\
        );

    \I__6460\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33643\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33690\,
            I => \N__33643\
        );

    \I__6458\ : InMux
    port map (
            O => \N__33689\,
            I => \N__33643\
        );

    \I__6457\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33634\
        );

    \I__6456\ : InMux
    port map (
            O => \N__33687\,
            I => \N__33634\
        );

    \I__6455\ : InMux
    port map (
            O => \N__33686\,
            I => \N__33634\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33634\
        );

    \I__6453\ : IoInMux
    port map (
            O => \N__33684\,
            I => \N__33631\
        );

    \I__6452\ : InMux
    port map (
            O => \N__33683\,
            I => \N__33628\
        );

    \I__6451\ : InMux
    port map (
            O => \N__33682\,
            I => \N__33619\
        );

    \I__6450\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33619\
        );

    \I__6449\ : InMux
    port map (
            O => \N__33680\,
            I => \N__33619\
        );

    \I__6448\ : InMux
    port map (
            O => \N__33679\,
            I => \N__33619\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33612\
        );

    \I__6446\ : InMux
    port map (
            O => \N__33677\,
            I => \N__33612\
        );

    \I__6445\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33612\
        );

    \I__6444\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33603\
        );

    \I__6443\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33603\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33603\
        );

    \I__6441\ : InMux
    port map (
            O => \N__33672\,
            I => \N__33603\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33671\,
            I => \N__33594\
        );

    \I__6439\ : InMux
    port map (
            O => \N__33670\,
            I => \N__33594\
        );

    \I__6438\ : InMux
    port map (
            O => \N__33669\,
            I => \N__33594\
        );

    \I__6437\ : InMux
    port map (
            O => \N__33668\,
            I => \N__33594\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__33659\,
            I => \N__33589\
        );

    \I__6435\ : LocalMux
    port map (
            O => \N__33650\,
            I => \N__33589\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__33643\,
            I => \N__33586\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__33634\,
            I => \N__33583\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__33631\,
            I => \N__33580\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33628\,
            I => \N__33573\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33619\,
            I => \N__33573\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__33612\,
            I => \N__33573\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__33603\,
            I => \N__33562\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__33594\,
            I => \N__33562\
        );

    \I__6426\ : Span4Mux_h
    port map (
            O => \N__33589\,
            I => \N__33562\
        );

    \I__6425\ : Span4Mux_v
    port map (
            O => \N__33586\,
            I => \N__33562\
        );

    \I__6424\ : Span4Mux_v
    port map (
            O => \N__33583\,
            I => \N__33562\
        );

    \I__6423\ : Span4Mux_s1_v
    port map (
            O => \N__33580\,
            I => \N__33559\
        );

    \I__6422\ : Span4Mux_v
    port map (
            O => \N__33573\,
            I => \N__33552\
        );

    \I__6421\ : Span4Mux_v
    port map (
            O => \N__33562\,
            I => \N__33552\
        );

    \I__6420\ : Span4Mux_v
    port map (
            O => \N__33559\,
            I => \N__33552\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__33552\,
            I => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\
        );

    \I__6418\ : InMux
    port map (
            O => \N__33549\,
            I => \N__33546\
        );

    \I__6417\ : LocalMux
    port map (
            O => \N__33546\,
            I => \current_shift_inst.control_input_axb_27\
        );

    \I__6416\ : ClkMux
    port map (
            O => \N__33543\,
            I => \N__33540\
        );

    \I__6415\ : GlobalMux
    port map (
            O => \N__33540\,
            I => \N__33537\
        );

    \I__6414\ : gio2CtrlBuf
    port map (
            O => \N__33537\,
            I => delay_hc_input_c_g
        );

    \I__6413\ : IoInMux
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__6412\ : LocalMux
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__6411\ : IoSpan4Mux
    port map (
            O => \N__33528\,
            I => \N__33525\
        );

    \I__6410\ : Span4Mux_s3_v
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__6409\ : Sp12to4
    port map (
            O => \N__33522\,
            I => \N__33519\
        );

    \I__6408\ : Odrv12
    port map (
            O => \N__33519\,
            I => s3_phy_c
        );

    \I__6407\ : IoInMux
    port map (
            O => \N__33516\,
            I => \N__33513\
        );

    \I__6406\ : LocalMux
    port map (
            O => \N__33513\,
            I => \N__33510\
        );

    \I__6405\ : Span4Mux_s0_v
    port map (
            O => \N__33510\,
            I => \N__33507\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__33507\,
            I => \GB_BUFFER_red_c_g_THRU_CO\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33504\,
            I => \N__33501\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__33501\,
            I => \phase_controller_inst1.state_ns_0_0_1\
        );

    \I__6401\ : CascadeMux
    port map (
            O => \N__33498\,
            I => \N__33492\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33489\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33496\,
            I => \N__33484\
        );

    \I__6398\ : InMux
    port map (
            O => \N__33495\,
            I => \N__33484\
        );

    \I__6397\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33481\
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33489\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__33484\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6394\ : LocalMux
    port map (
            O => \N__33481\,
            I => \phase_controller_inst1.tr_time_passed\
        );

    \I__6393\ : CascadeMux
    port map (
            O => \N__33474\,
            I => \N__33470\
        );

    \I__6392\ : InMux
    port map (
            O => \N__33473\,
            I => \N__33466\
        );

    \I__6391\ : InMux
    port map (
            O => \N__33470\,
            I => \N__33463\
        );

    \I__6390\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33460\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33466\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6388\ : LocalMux
    port map (
            O => \N__33463\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__33460\,
            I => \phase_controller_inst1.stateZ0Z_0\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33453\,
            I => \N__33444\
        );

    \I__6385\ : InMux
    port map (
            O => \N__33452\,
            I => \N__33444\
        );

    \I__6384\ : InMux
    port map (
            O => \N__33451\,
            I => \N__33444\
        );

    \I__6383\ : LocalMux
    port map (
            O => \N__33444\,
            I => \phase_controller_inst1.stateZ0Z_4\
        );

    \I__6382\ : InMux
    port map (
            O => \N__33441\,
            I => \N__33438\
        );

    \I__6381\ : LocalMux
    port map (
            O => \N__33438\,
            I => \current_shift_inst.control_input_axb_14\
        );

    \I__6380\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33432\
        );

    \I__6379\ : LocalMux
    port map (
            O => \N__33432\,
            I => \current_shift_inst.control_input_axb_16\
        );

    \I__6378\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33426\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__33426\,
            I => \current_shift_inst.control_input_axb_18\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33423\,
            I => \N__33420\
        );

    \I__6375\ : LocalMux
    port map (
            O => \N__33420\,
            I => \current_shift_inst.control_input_axb_19\
        );

    \I__6374\ : InMux
    port map (
            O => \N__33417\,
            I => \N__33414\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__33414\,
            I => \current_shift_inst.control_input_axb_20\
        );

    \I__6372\ : InMux
    port map (
            O => \N__33411\,
            I => \N__33408\
        );

    \I__6371\ : LocalMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__6370\ : Odrv4
    port map (
            O => \N__33405\,
            I => \current_shift_inst.control_input_axb_10\
        );

    \I__6369\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__33399\,
            I => \current_shift_inst.control_input_axb_23\
        );

    \I__6367\ : InMux
    port map (
            O => \N__33396\,
            I => \N__33393\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__33393\,
            I => \current_shift_inst.control_input_axb_24\
        );

    \I__6365\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__6364\ : LocalMux
    port map (
            O => \N__33387\,
            I => \current_shift_inst.control_input_axb_25\
        );

    \I__6363\ : InMux
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__33381\,
            I => \current_shift_inst.control_input_axb_9\
        );

    \I__6361\ : InMux
    port map (
            O => \N__33378\,
            I => \N__33375\
        );

    \I__6360\ : LocalMux
    port map (
            O => \N__33375\,
            I => \current_shift_inst.control_input_axb_12\
        );

    \I__6359\ : InMux
    port map (
            O => \N__33372\,
            I => \N__33369\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__33369\,
            I => \current_shift_inst.control_input_axb_13\
        );

    \I__6357\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33363\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33363\,
            I => \current_shift_inst.control_input_axb_11\
        );

    \I__6355\ : InMux
    port map (
            O => \N__33360\,
            I => \N__33357\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__33357\,
            I => \current_shift_inst.control_input_axb_15\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33350\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33347\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__33350\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__33347\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\
        );

    \I__6349\ : CEMux
    port map (
            O => \N__33342\,
            I => \N__33306\
        );

    \I__6348\ : CEMux
    port map (
            O => \N__33341\,
            I => \N__33306\
        );

    \I__6347\ : CEMux
    port map (
            O => \N__33340\,
            I => \N__33306\
        );

    \I__6346\ : CEMux
    port map (
            O => \N__33339\,
            I => \N__33306\
        );

    \I__6345\ : CEMux
    port map (
            O => \N__33338\,
            I => \N__33306\
        );

    \I__6344\ : CEMux
    port map (
            O => \N__33337\,
            I => \N__33306\
        );

    \I__6343\ : CEMux
    port map (
            O => \N__33336\,
            I => \N__33306\
        );

    \I__6342\ : CEMux
    port map (
            O => \N__33335\,
            I => \N__33306\
        );

    \I__6341\ : CEMux
    port map (
            O => \N__33334\,
            I => \N__33306\
        );

    \I__6340\ : CEMux
    port map (
            O => \N__33333\,
            I => \N__33306\
        );

    \I__6339\ : CEMux
    port map (
            O => \N__33332\,
            I => \N__33306\
        );

    \I__6338\ : CEMux
    port map (
            O => \N__33331\,
            I => \N__33306\
        );

    \I__6337\ : GlobalMux
    port map (
            O => \N__33306\,
            I => \N__33303\
        );

    \I__6336\ : gio2CtrlBuf
    port map (
            O => \N__33303\,
            I => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33297\
        );

    \I__6334\ : LocalMux
    port map (
            O => \N__33297\,
            I => \current_shift_inst.control_input_axb_2\
        );

    \I__6333\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33290\
        );

    \I__6332\ : InMux
    port map (
            O => \N__33293\,
            I => \N__33287\
        );

    \I__6331\ : LocalMux
    port map (
            O => \N__33290\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__6330\ : LocalMux
    port map (
            O => \N__33287\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\
        );

    \I__6329\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33277\
        );

    \I__6328\ : InMux
    port map (
            O => \N__33281\,
            I => \N__33274\
        );

    \I__6327\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33271\
        );

    \I__6326\ : LocalMux
    port map (
            O => \N__33277\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6325\ : LocalMux
    port map (
            O => \N__33274\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6324\ : LocalMux
    port map (
            O => \N__33271\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__6323\ : CascadeMux
    port map (
            O => \N__33264\,
            I => \N__33260\
        );

    \I__6322\ : CascadeMux
    port map (
            O => \N__33263\,
            I => \N__33257\
        );

    \I__6321\ : InMux
    port map (
            O => \N__33260\,
            I => \N__33254\
        );

    \I__6320\ : InMux
    port map (
            O => \N__33257\,
            I => \N__33251\
        );

    \I__6319\ : LocalMux
    port map (
            O => \N__33254\,
            I => \N__33246\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__33251\,
            I => \N__33246\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__33246\,
            I => \N__33243\
        );

    \I__6316\ : Odrv4
    port map (
            O => \N__33243\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\
        );

    \I__6315\ : InMux
    port map (
            O => \N__33240\,
            I => \N__33235\
        );

    \I__6314\ : InMux
    port map (
            O => \N__33239\,
            I => \N__33232\
        );

    \I__6313\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33229\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__33235\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__6311\ : LocalMux
    port map (
            O => \N__33232\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__33229\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__6309\ : InMux
    port map (
            O => \N__33222\,
            I => \N__33219\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__33219\,
            I => \N__33216\
        );

    \I__6307\ : Span4Mux_h
    port map (
            O => \N__33216\,
            I => \N__33213\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__33213\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt28\
        );

    \I__6305\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__33207\,
            I => \current_shift_inst.control_input_axb_6\
        );

    \I__6303\ : CascadeMux
    port map (
            O => \N__33204\,
            I => \N__33198\
        );

    \I__6302\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33195\
        );

    \I__6301\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33192\
        );

    \I__6300\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33189\
        );

    \I__6299\ : InMux
    port map (
            O => \N__33198\,
            I => \N__33186\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__33195\,
            I => \N__33183\
        );

    \I__6297\ : LocalMux
    port map (
            O => \N__33192\,
            I => \N__33180\
        );

    \I__6296\ : LocalMux
    port map (
            O => \N__33189\,
            I => \N__33175\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__33186\,
            I => \N__33175\
        );

    \I__6294\ : Span4Mux_v
    port map (
            O => \N__33183\,
            I => \N__33172\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__33180\,
            I => \N__33169\
        );

    \I__6292\ : Span4Mux_v
    port map (
            O => \N__33175\,
            I => \N__33166\
        );

    \I__6291\ : Odrv4
    port map (
            O => \N__33172\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__6290\ : Odrv4
    port map (
            O => \N__33169\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__6289\ : Odrv4
    port map (
            O => \N__33166\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\
        );

    \I__6288\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33156\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33152\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33155\,
            I => \N__33149\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__33152\,
            I => \N__33143\
        );

    \I__6284\ : LocalMux
    port map (
            O => \N__33149\,
            I => \N__33143\
        );

    \I__6283\ : InMux
    port map (
            O => \N__33148\,
            I => \N__33140\
        );

    \I__6282\ : Span4Mux_h
    port map (
            O => \N__33143\,
            I => \N__33137\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__33140\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__6280\ : Odrv4
    port map (
            O => \N__33137\,
            I => \elapsed_time_ns_1_RNIU8PBB_0_20\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__33132\,
            I => \N__33129\
        );

    \I__6278\ : InMux
    port map (
            O => \N__33129\,
            I => \N__33126\
        );

    \I__6277\ : LocalMux
    port map (
            O => \N__33126\,
            I => \N__33123\
        );

    \I__6276\ : Odrv4
    port map (
            O => \N__33123\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\
        );

    \I__6275\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33114\
        );

    \I__6274\ : InMux
    port map (
            O => \N__33119\,
            I => \N__33114\
        );

    \I__6273\ : LocalMux
    port map (
            O => \N__33114\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__6271\ : InMux
    port map (
            O => \N__33108\,
            I => \N__33102\
        );

    \I__6270\ : InMux
    port map (
            O => \N__33107\,
            I => \N__33102\
        );

    \I__6269\ : LocalMux
    port map (
            O => \N__33102\,
            I => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\
        );

    \I__6268\ : InMux
    port map (
            O => \N__33099\,
            I => \N__33096\
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__33096\,
            I => \N__33093\
        );

    \I__6266\ : Span4Mux_h
    port map (
            O => \N__33093\,
            I => \N__33090\
        );

    \I__6265\ : Odrv4
    port map (
            O => \N__33090\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt16\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__6263\ : InMux
    port map (
            O => \N__33084\,
            I => \N__33081\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33081\,
            I => \N__33078\
        );

    \I__6261\ : Span4Mux_v
    port map (
            O => \N__33078\,
            I => \N__33075\
        );

    \I__6260\ : Odrv4
    port map (
            O => \N__33075\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\
        );

    \I__6259\ : InMux
    port map (
            O => \N__33072\,
            I => \N__33069\
        );

    \I__6258\ : LocalMux
    port map (
            O => \N__33069\,
            I => \N__33064\
        );

    \I__6257\ : InMux
    port map (
            O => \N__33068\,
            I => \N__33061\
        );

    \I__6256\ : InMux
    port map (
            O => \N__33067\,
            I => \N__33058\
        );

    \I__6255\ : Span4Mux_h
    port map (
            O => \N__33064\,
            I => \N__33054\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__33061\,
            I => \N__33051\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__33058\,
            I => \N__33048\
        );

    \I__6252\ : InMux
    port map (
            O => \N__33057\,
            I => \N__33045\
        );

    \I__6251\ : Span4Mux_v
    port map (
            O => \N__33054\,
            I => \N__33042\
        );

    \I__6250\ : Span4Mux_h
    port map (
            O => \N__33051\,
            I => \N__33037\
        );

    \I__6249\ : Span4Mux_v
    port map (
            O => \N__33048\,
            I => \N__33037\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__33045\,
            I => \N__33034\
        );

    \I__6247\ : Odrv4
    port map (
            O => \N__33042\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__6246\ : Odrv4
    port map (
            O => \N__33037\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__6245\ : Odrv12
    port map (
            O => \N__33034\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\
        );

    \I__6244\ : InMux
    port map (
            O => \N__33027\,
            I => \N__33023\
        );

    \I__6243\ : InMux
    port map (
            O => \N__33026\,
            I => \N__33019\
        );

    \I__6242\ : LocalMux
    port map (
            O => \N__33023\,
            I => \N__33016\
        );

    \I__6241\ : InMux
    port map (
            O => \N__33022\,
            I => \N__33013\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__33019\,
            I => \N__33008\
        );

    \I__6239\ : Span4Mux_v
    port map (
            O => \N__33016\,
            I => \N__33008\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__33013\,
            I => \N__33005\
        );

    \I__6237\ : Odrv4
    port map (
            O => \N__33008\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__6236\ : Odrv4
    port map (
            O => \N__33005\,
            I => \elapsed_time_ns_1_RNI6HPBB_0_28\
        );

    \I__6235\ : InMux
    port map (
            O => \N__33000\,
            I => \N__32995\
        );

    \I__6234\ : InMux
    port map (
            O => \N__32999\,
            I => \N__32992\
        );

    \I__6233\ : InMux
    port map (
            O => \N__32998\,
            I => \N__32989\
        );

    \I__6232\ : LocalMux
    port map (
            O => \N__32995\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6231\ : LocalMux
    port map (
            O => \N__32992\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__32989\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__6229\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32978\
        );

    \I__6228\ : InMux
    port map (
            O => \N__32981\,
            I => \N__32975\
        );

    \I__6227\ : LocalMux
    port map (
            O => \N__32978\,
            I => \N__32970\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32970\
        );

    \I__6225\ : Odrv12
    port map (
            O => \N__32970\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\
        );

    \I__6224\ : CascadeMux
    port map (
            O => \N__32967\,
            I => \N__32963\
        );

    \I__6223\ : CascadeMux
    port map (
            O => \N__32966\,
            I => \N__32959\
        );

    \I__6222\ : InMux
    port map (
            O => \N__32963\,
            I => \N__32956\
        );

    \I__6221\ : InMux
    port map (
            O => \N__32962\,
            I => \N__32953\
        );

    \I__6220\ : InMux
    port map (
            O => \N__32959\,
            I => \N__32950\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__32956\,
            I => \N__32947\
        );

    \I__6218\ : LocalMux
    port map (
            O => \N__32953\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6217\ : LocalMux
    port map (
            O => \N__32950\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6216\ : Odrv4
    port map (
            O => \N__32947\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__6215\ : CascadeMux
    port map (
            O => \N__32940\,
            I => \N__32937\
        );

    \I__6214\ : InMux
    port map (
            O => \N__32937\,
            I => \N__32934\
        );

    \I__6213\ : LocalMux
    port map (
            O => \N__32934\,
            I => \N__32931\
        );

    \I__6212\ : Span4Mux_h
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__6211\ : Span4Mux_h
    port map (
            O => \N__32928\,
            I => \N__32925\
        );

    \I__6210\ : Odrv4
    port map (
            O => \N__32925\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\
        );

    \I__6209\ : InMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__6207\ : Span4Mux_v
    port map (
            O => \N__32916\,
            I => \N__32911\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32915\,
            I => \N__32906\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32914\,
            I => \N__32906\
        );

    \I__6204\ : Sp12to4
    port map (
            O => \N__32911\,
            I => \N__32901\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32906\,
            I => \N__32901\
        );

    \I__6202\ : Span12Mux_h
    port map (
            O => \N__32901\,
            I => \N__32898\
        );

    \I__6201\ : Odrv12
    port map (
            O => \N__32898\,
            I => il_max_comp2_c
        );

    \I__6200\ : InMux
    port map (
            O => \N__32895\,
            I => \N__32892\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__32892\,
            I => \N__32889\
        );

    \I__6198\ : Span4Mux_v
    port map (
            O => \N__32889\,
            I => \N__32884\
        );

    \I__6197\ : InMux
    port map (
            O => \N__32888\,
            I => \N__32881\
        );

    \I__6196\ : InMux
    port map (
            O => \N__32887\,
            I => \N__32878\
        );

    \I__6195\ : Sp12to4
    port map (
            O => \N__32884\,
            I => \N__32871\
        );

    \I__6194\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32871\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__32878\,
            I => \N__32871\
        );

    \I__6192\ : Span12Mux_h
    port map (
            O => \N__32871\,
            I => \N__32868\
        );

    \I__6191\ : Odrv12
    port map (
            O => \N__32868\,
            I => il_min_comp2_c
        );

    \I__6190\ : InMux
    port map (
            O => \N__32865\,
            I => \N__32862\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__6188\ : Span4Mux_v
    port map (
            O => \N__32859\,
            I => \N__32855\
        );

    \I__6187\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32851\
        );

    \I__6186\ : Sp12to4
    port map (
            O => \N__32855\,
            I => \N__32848\
        );

    \I__6185\ : InMux
    port map (
            O => \N__32854\,
            I => \N__32844\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__32851\,
            I => \N__32839\
        );

    \I__6183\ : Span12Mux_v
    port map (
            O => \N__32848\,
            I => \N__32839\
        );

    \I__6182\ : InMux
    port map (
            O => \N__32847\,
            I => \N__32836\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__32844\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6180\ : Odrv12
    port map (
            O => \N__32839\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__32836\,
            I => \phase_controller_inst2.stateZ0Z_1\
        );

    \I__6178\ : InMux
    port map (
            O => \N__32829\,
            I => \N__32824\
        );

    \I__6177\ : InMux
    port map (
            O => \N__32828\,
            I => \N__32821\
        );

    \I__6176\ : InMux
    port map (
            O => \N__32827\,
            I => \N__32818\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32824\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__32821\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__32818\,
            I => \phase_controller_inst2.stateZ0Z_0\
        );

    \I__6172\ : InMux
    port map (
            O => \N__32811\,
            I => \N__32808\
        );

    \I__6171\ : LocalMux
    port map (
            O => \N__32808\,
            I => \N__32805\
        );

    \I__6170\ : Odrv4
    port map (
            O => \N__32805\,
            I => \phase_controller_inst2.N_54_0\
        );

    \I__6169\ : CascadeMux
    port map (
            O => \N__32802\,
            I => \N__32798\
        );

    \I__6168\ : CascadeMux
    port map (
            O => \N__32801\,
            I => \N__32793\
        );

    \I__6167\ : InMux
    port map (
            O => \N__32798\,
            I => \N__32790\
        );

    \I__6166\ : InMux
    port map (
            O => \N__32797\,
            I => \N__32785\
        );

    \I__6165\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32785\
        );

    \I__6164\ : InMux
    port map (
            O => \N__32793\,
            I => \N__32782\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32790\,
            I => \N__32779\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__32785\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__32782\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__32779\,
            I => \phase_controller_inst2.tr_time_passed\
        );

    \I__6159\ : CascadeMux
    port map (
            O => \N__32772\,
            I => \N__32767\
        );

    \I__6158\ : CascadeMux
    port map (
            O => \N__32771\,
            I => \N__32764\
        );

    \I__6157\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32761\
        );

    \I__6156\ : InMux
    port map (
            O => \N__32767\,
            I => \N__32758\
        );

    \I__6155\ : InMux
    port map (
            O => \N__32764\,
            I => \N__32755\
        );

    \I__6154\ : LocalMux
    port map (
            O => \N__32761\,
            I => \N__32752\
        );

    \I__6153\ : LocalMux
    port map (
            O => \N__32758\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32755\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__32752\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__6150\ : CascadeMux
    port map (
            O => \N__32745\,
            I => \N__32741\
        );

    \I__6149\ : CascadeMux
    port map (
            O => \N__32744\,
            I => \N__32738\
        );

    \I__6148\ : InMux
    port map (
            O => \N__32741\,
            I => \N__32734\
        );

    \I__6147\ : InMux
    port map (
            O => \N__32738\,
            I => \N__32729\
        );

    \I__6146\ : InMux
    port map (
            O => \N__32737\,
            I => \N__32729\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__32734\,
            I => \N__32726\
        );

    \I__6144\ : LocalMux
    port map (
            O => \N__32729\,
            I => \N__32723\
        );

    \I__6143\ : Span4Mux_h
    port map (
            O => \N__32726\,
            I => \N__32720\
        );

    \I__6142\ : Span4Mux_h
    port map (
            O => \N__32723\,
            I => \N__32717\
        );

    \I__6141\ : Odrv4
    port map (
            O => \N__32720\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6140\ : Odrv4
    port map (
            O => \N__32717\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6139\ : CascadeMux
    port map (
            O => \N__32712\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__6138\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32706\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__32706\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\
        );

    \I__6136\ : InMux
    port map (
            O => \N__32703\,
            I => \N__32699\
        );

    \I__6135\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32696\
        );

    \I__6134\ : LocalMux
    port map (
            O => \N__32699\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__32696\,
            I => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\
        );

    \I__6132\ : InMux
    port map (
            O => \N__32691\,
            I => \N__32688\
        );

    \I__6131\ : LocalMux
    port map (
            O => \N__32688\,
            I => \N__32685\
        );

    \I__6130\ : Span4Mux_v
    port map (
            O => \N__32685\,
            I => \N__32680\
        );

    \I__6129\ : InMux
    port map (
            O => \N__32684\,
            I => \N__32677\
        );

    \I__6128\ : InMux
    port map (
            O => \N__32683\,
            I => \N__32674\
        );

    \I__6127\ : Span4Mux_h
    port map (
            O => \N__32680\,
            I => \N__32669\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__32677\,
            I => \N__32669\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__32674\,
            I => \N__32666\
        );

    \I__6124\ : Sp12to4
    port map (
            O => \N__32669\,
            I => \N__32663\
        );

    \I__6123\ : Span4Mux_h
    port map (
            O => \N__32666\,
            I => \N__32659\
        );

    \I__6122\ : Span12Mux_s10_v
    port map (
            O => \N__32663\,
            I => \N__32656\
        );

    \I__6121\ : InMux
    port map (
            O => \N__32662\,
            I => \N__32653\
        );

    \I__6120\ : Odrv4
    port map (
            O => \N__32659\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__6119\ : Odrv12
    port map (
            O => \N__32656\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32653\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\
        );

    \I__6117\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32643\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__32643\,
            I => \N__32640\
        );

    \I__6115\ : Span4Mux_h
    port map (
            O => \N__32640\,
            I => \N__32635\
        );

    \I__6114\ : InMux
    port map (
            O => \N__32639\,
            I => \N__32632\
        );

    \I__6113\ : InMux
    port map (
            O => \N__32638\,
            I => \N__32629\
        );

    \I__6112\ : Span4Mux_v
    port map (
            O => \N__32635\,
            I => \N__32626\
        );

    \I__6111\ : LocalMux
    port map (
            O => \N__32632\,
            I => \N__32623\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__32629\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__6109\ : Odrv4
    port map (
            O => \N__32626\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__6108\ : Odrv12
    port map (
            O => \N__32623\,
            I => \elapsed_time_ns_1_RNIDC91B_0_1\
        );

    \I__6107\ : InMux
    port map (
            O => \N__32616\,
            I => \N__32612\
        );

    \I__6106\ : CascadeMux
    port map (
            O => \N__32615\,
            I => \N__32609\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__32612\,
            I => \N__32606\
        );

    \I__6104\ : InMux
    port map (
            O => \N__32609\,
            I => \N__32600\
        );

    \I__6103\ : Span4Mux_s2_v
    port map (
            O => \N__32606\,
            I => \N__32597\
        );

    \I__6102\ : InMux
    port map (
            O => \N__32605\,
            I => \N__32590\
        );

    \I__6101\ : InMux
    port map (
            O => \N__32604\,
            I => \N__32590\
        );

    \I__6100\ : InMux
    port map (
            O => \N__32603\,
            I => \N__32590\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__32600\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6098\ : Odrv4
    port map (
            O => \N__32597\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__32590\,
            I => \phase_controller_inst1.stoper_tr.un2_start_0\
        );

    \I__6096\ : CascadeMux
    port map (
            O => \N__32583\,
            I => \N__32579\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32582\,
            I => \N__32576\
        );

    \I__6094\ : InMux
    port map (
            O => \N__32579\,
            I => \N__32572\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__32576\,
            I => \N__32569\
        );

    \I__6092\ : InMux
    port map (
            O => \N__32575\,
            I => \N__32566\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__32572\,
            I => \N__32559\
        );

    \I__6090\ : Span4Mux_h
    port map (
            O => \N__32569\,
            I => \N__32559\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__32566\,
            I => \N__32559\
        );

    \I__6088\ : Odrv4
    port map (
            O => \N__32559\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\
        );

    \I__6087\ : CascadeMux
    port map (
            O => \N__32556\,
            I => \N__32552\
        );

    \I__6086\ : InMux
    port map (
            O => \N__32555\,
            I => \N__32545\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32552\,
            I => \N__32545\
        );

    \I__6084\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32540\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32550\,
            I => \N__32540\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__32545\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6081\ : LocalMux
    port map (
            O => \N__32540\,
            I => \phase_controller_inst1.start_timer_trZ0\
        );

    \I__6080\ : InMux
    port map (
            O => \N__32535\,
            I => \N__32528\
        );

    \I__6079\ : InMux
    port map (
            O => \N__32534\,
            I => \N__32528\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32533\,
            I => \N__32523\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__32528\,
            I => \N__32520\
        );

    \I__6076\ : InMux
    port map (
            O => \N__32527\,
            I => \N__32515\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32526\,
            I => \N__32515\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32523\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6073\ : Odrv4
    port map (
            O => \N__32520\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32515\,
            I => \phase_controller_inst1.stoper_tr.start_latchedZ0\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32508\,
            I => \N__32503\
        );

    \I__6070\ : InMux
    port map (
            O => \N__32507\,
            I => \N__32500\
        );

    \I__6069\ : InMux
    port map (
            O => \N__32506\,
            I => \N__32497\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__32503\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6067\ : LocalMux
    port map (
            O => \N__32500\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32497\,
            I => \elapsed_time_ns_1_RNI3DOBB_0_16\
        );

    \I__6065\ : InMux
    port map (
            O => \N__32490\,
            I => \N__32487\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__32487\,
            I => \N__32482\
        );

    \I__6063\ : InMux
    port map (
            O => \N__32486\,
            I => \N__32479\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32485\,
            I => \N__32476\
        );

    \I__6061\ : Span4Mux_h
    port map (
            O => \N__32482\,
            I => \N__32471\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32479\,
            I => \N__32471\
        );

    \I__6059\ : LocalMux
    port map (
            O => \N__32476\,
            I => \N__32467\
        );

    \I__6058\ : Span4Mux_h
    port map (
            O => \N__32471\,
            I => \N__32464\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32461\
        );

    \I__6056\ : Span12Mux_s11_v
    port map (
            O => \N__32467\,
            I => \N__32458\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__32464\,
            I => \N__32453\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__32461\,
            I => \N__32453\
        );

    \I__6053\ : Odrv12
    port map (
            O => \N__32458\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6052\ : Odrv4
    port map (
            O => \N__32453\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\
        );

    \I__6051\ : InMux
    port map (
            O => \N__32448\,
            I => \N__32445\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32445\,
            I => \N__32442\
        );

    \I__6049\ : Odrv4
    port map (
            O => \N__32442\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\
        );

    \I__6048\ : InMux
    port map (
            O => \N__32439\,
            I => \current_shift_inst.control_input_cry_25\
        );

    \I__6047\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32433\
        );

    \I__6046\ : LocalMux
    port map (
            O => \N__32433\,
            I => \N__32430\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__32430\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\
        );

    \I__6044\ : InMux
    port map (
            O => \N__32427\,
            I => \current_shift_inst.control_input_cry_26\
        );

    \I__6043\ : CascadeMux
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__32418\,
            I => \N__32415\
        );

    \I__6040\ : Odrv4
    port map (
            O => \N__32415\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\
        );

    \I__6039\ : InMux
    port map (
            O => \N__32412\,
            I => \current_shift_inst.control_input_cry_27\
        );

    \I__6038\ : CascadeMux
    port map (
            O => \N__32409\,
            I => \N__32406\
        );

    \I__6037\ : InMux
    port map (
            O => \N__32406\,
            I => \N__32403\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__32403\,
            I => \N__32400\
        );

    \I__6035\ : Odrv4
    port map (
            O => \N__32400\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32397\,
            I => \current_shift_inst.control_input_cry_28\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32394\,
            I => \current_shift_inst.control_input_cry_29\
        );

    \I__6032\ : InMux
    port map (
            O => \N__32391\,
            I => \N__32388\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__32388\,
            I => \N__32384\
        );

    \I__6030\ : InMux
    port map (
            O => \N__32387\,
            I => \N__32381\
        );

    \I__6029\ : Odrv4
    port map (
            O => \N__32384\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6028\ : LocalMux
    port map (
            O => \N__32381\,
            I => \current_shift_inst.control_input_31\
        );

    \I__6027\ : InMux
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__6026\ : LocalMux
    port map (
            O => \N__32373\,
            I => \current_shift_inst.control_input_axb_26\
        );

    \I__6025\ : InMux
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32367\,
            I => \current_shift_inst.control_input_axb_29\
        );

    \I__6023\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32361\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__32361\,
            I => \N__32358\
        );

    \I__6021\ : Odrv4
    port map (
            O => \N__32358\,
            I => \current_shift_inst.control_input_axb_17\
        );

    \I__6020\ : IoInMux
    port map (
            O => \N__32355\,
            I => \N__32352\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__32352\,
            I => \N__32349\
        );

    \I__6018\ : IoSpan4Mux
    port map (
            O => \N__32349\,
            I => \N__32346\
        );

    \I__6017\ : Span4Mux_s2_v
    port map (
            O => \N__32346\,
            I => \N__32343\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__32343\,
            I => s4_phy_c
        );

    \I__6015\ : InMux
    port map (
            O => \N__32340\,
            I => \N__32337\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__32337\,
            I => \N__32334\
        );

    \I__6013\ : Odrv4
    port map (
            O => \N__32334\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\
        );

    \I__6012\ : InMux
    port map (
            O => \N__32331\,
            I => \current_shift_inst.control_input_cry_17\
        );

    \I__6011\ : InMux
    port map (
            O => \N__32328\,
            I => \N__32325\
        );

    \I__6010\ : LocalMux
    port map (
            O => \N__32325\,
            I => \N__32322\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__32322\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\
        );

    \I__6008\ : InMux
    port map (
            O => \N__32319\,
            I => \current_shift_inst.control_input_cry_18\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__32316\,
            I => \N__32313\
        );

    \I__6006\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32310\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__32310\,
            I => \N__32307\
        );

    \I__6004\ : Odrv4
    port map (
            O => \N__32307\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\
        );

    \I__6003\ : InMux
    port map (
            O => \N__32304\,
            I => \current_shift_inst.control_input_cry_19\
        );

    \I__6002\ : InMux
    port map (
            O => \N__32301\,
            I => \N__32298\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__32298\,
            I => \N__32295\
        );

    \I__6000\ : Odrv4
    port map (
            O => \N__32295\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\
        );

    \I__5999\ : InMux
    port map (
            O => \N__32292\,
            I => \current_shift_inst.control_input_cry_20\
        );

    \I__5998\ : CascadeMux
    port map (
            O => \N__32289\,
            I => \N__32286\
        );

    \I__5997\ : InMux
    port map (
            O => \N__32286\,
            I => \N__32283\
        );

    \I__5996\ : LocalMux
    port map (
            O => \N__32283\,
            I => \N__32280\
        );

    \I__5995\ : Odrv4
    port map (
            O => \N__32280\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\
        );

    \I__5994\ : InMux
    port map (
            O => \N__32277\,
            I => \current_shift_inst.control_input_cry_21\
        );

    \I__5993\ : CascadeMux
    port map (
            O => \N__32274\,
            I => \N__32271\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32268\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__32268\,
            I => \N__32265\
        );

    \I__5990\ : Odrv4
    port map (
            O => \N__32265\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\
        );

    \I__5989\ : InMux
    port map (
            O => \N__32262\,
            I => \current_shift_inst.control_input_cry_22\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32259\,
            I => \N__32256\
        );

    \I__5987\ : LocalMux
    port map (
            O => \N__32256\,
            I => \N__32253\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__32253\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\
        );

    \I__5985\ : InMux
    port map (
            O => \N__32250\,
            I => \bfn_11_16_0_\
        );

    \I__5984\ : InMux
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__5983\ : LocalMux
    port map (
            O => \N__32244\,
            I => \N__32241\
        );

    \I__5982\ : Odrv4
    port map (
            O => \N__32241\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\
        );

    \I__5981\ : InMux
    port map (
            O => \N__32238\,
            I => \current_shift_inst.control_input_cry_24\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__32235\,
            I => \N__32232\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32232\,
            I => \N__32229\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__32229\,
            I => \N__32226\
        );

    \I__5977\ : Odrv4
    port map (
            O => \N__32226\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\
        );

    \I__5976\ : InMux
    port map (
            O => \N__32223\,
            I => \current_shift_inst.control_input_cry_9\
        );

    \I__5975\ : InMux
    port map (
            O => \N__32220\,
            I => \N__32217\
        );

    \I__5974\ : LocalMux
    port map (
            O => \N__32217\,
            I => \N__32214\
        );

    \I__5973\ : Odrv4
    port map (
            O => \N__32214\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\
        );

    \I__5972\ : InMux
    port map (
            O => \N__32211\,
            I => \current_shift_inst.control_input_cry_10\
        );

    \I__5971\ : InMux
    port map (
            O => \N__32208\,
            I => \N__32205\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__32205\,
            I => \N__32202\
        );

    \I__5969\ : Odrv4
    port map (
            O => \N__32202\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32199\,
            I => \current_shift_inst.control_input_cry_11\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__32196\,
            I => \N__32193\
        );

    \I__5966\ : InMux
    port map (
            O => \N__32193\,
            I => \N__32190\
        );

    \I__5965\ : LocalMux
    port map (
            O => \N__32190\,
            I => \N__32187\
        );

    \I__5964\ : Odrv4
    port map (
            O => \N__32187\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\
        );

    \I__5963\ : InMux
    port map (
            O => \N__32184\,
            I => \current_shift_inst.control_input_cry_12\
        );

    \I__5962\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32178\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__32178\,
            I => \N__32175\
        );

    \I__5960\ : Odrv4
    port map (
            O => \N__32175\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32172\,
            I => \current_shift_inst.control_input_cry_13\
        );

    \I__5958\ : CascadeMux
    port map (
            O => \N__32169\,
            I => \N__32166\
        );

    \I__5957\ : InMux
    port map (
            O => \N__32166\,
            I => \N__32163\
        );

    \I__5956\ : LocalMux
    port map (
            O => \N__32163\,
            I => \N__32160\
        );

    \I__5955\ : Odrv4
    port map (
            O => \N__32160\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\
        );

    \I__5954\ : InMux
    port map (
            O => \N__32157\,
            I => \current_shift_inst.control_input_cry_14\
        );

    \I__5953\ : InMux
    port map (
            O => \N__32154\,
            I => \N__32151\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__32151\,
            I => \N__32148\
        );

    \I__5951\ : Odrv4
    port map (
            O => \N__32148\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32145\,
            I => \bfn_11_15_0_\
        );

    \I__5949\ : CascadeMux
    port map (
            O => \N__32142\,
            I => \N__32139\
        );

    \I__5948\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__32136\,
            I => \N__32133\
        );

    \I__5946\ : Odrv4
    port map (
            O => \N__32133\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\
        );

    \I__5945\ : InMux
    port map (
            O => \N__32130\,
            I => \current_shift_inst.control_input_cry_16\
        );

    \I__5944\ : InMux
    port map (
            O => \N__32127\,
            I => \N__32124\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32124\,
            I => \N__32121\
        );

    \I__5942\ : Odrv4
    port map (
            O => \N__32121\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32118\,
            I => \current_shift_inst.control_input_cry_0\
        );

    \I__5940\ : CascadeMux
    port map (
            O => \N__32115\,
            I => \N__32112\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32112\,
            I => \N__32109\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__32109\,
            I => \N__32106\
        );

    \I__5937\ : Odrv4
    port map (
            O => \N__32106\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32103\,
            I => \current_shift_inst.control_input_cry_1\
        );

    \I__5935\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32097\
        );

    \I__5934\ : LocalMux
    port map (
            O => \N__32097\,
            I => \N__32094\
        );

    \I__5933\ : Odrv4
    port map (
            O => \N__32094\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\
        );

    \I__5932\ : InMux
    port map (
            O => \N__32091\,
            I => \current_shift_inst.control_input_cry_2\
        );

    \I__5931\ : InMux
    port map (
            O => \N__32088\,
            I => \N__32085\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__5929\ : Odrv4
    port map (
            O => \N__32082\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\
        );

    \I__5928\ : InMux
    port map (
            O => \N__32079\,
            I => \current_shift_inst.control_input_cry_3\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__32076\,
            I => \N__32073\
        );

    \I__5926\ : InMux
    port map (
            O => \N__32073\,
            I => \N__32070\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__32070\,
            I => \N__32067\
        );

    \I__5924\ : Odrv4
    port map (
            O => \N__32067\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\
        );

    \I__5923\ : InMux
    port map (
            O => \N__32064\,
            I => \current_shift_inst.control_input_cry_4\
        );

    \I__5922\ : InMux
    port map (
            O => \N__32061\,
            I => \N__32058\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__32058\,
            I => \N__32055\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__32055\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\
        );

    \I__5919\ : InMux
    port map (
            O => \N__32052\,
            I => \current_shift_inst.control_input_cry_5\
        );

    \I__5918\ : CascadeMux
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__5917\ : InMux
    port map (
            O => \N__32046\,
            I => \N__32043\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__32043\,
            I => \N__32040\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__32040\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\
        );

    \I__5914\ : InMux
    port map (
            O => \N__32037\,
            I => \current_shift_inst.control_input_cry_6\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__32034\,
            I => \N__32031\
        );

    \I__5912\ : InMux
    port map (
            O => \N__32031\,
            I => \N__32028\
        );

    \I__5911\ : LocalMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__5910\ : Odrv4
    port map (
            O => \N__32025\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32022\,
            I => \bfn_11_14_0_\
        );

    \I__5908\ : InMux
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__5907\ : LocalMux
    port map (
            O => \N__32016\,
            I => \N__32013\
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__32013\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\
        );

    \I__5905\ : InMux
    port map (
            O => \N__32010\,
            I => \current_shift_inst.control_input_cry_8\
        );

    \I__5904\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32002\
        );

    \I__5903\ : InMux
    port map (
            O => \N__32006\,
            I => \N__31997\
        );

    \I__5902\ : InMux
    port map (
            O => \N__32005\,
            I => \N__31997\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__32002\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__31997\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__5899\ : InMux
    port map (
            O => \N__31992\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__5898\ : CascadeMux
    port map (
            O => \N__31989\,
            I => \N__31985\
        );

    \I__5897\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31979\
        );

    \I__5896\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31979\
        );

    \I__5895\ : InMux
    port map (
            O => \N__31984\,
            I => \N__31976\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31973\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__31976\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5892\ : Odrv4
    port map (
            O => \N__31973\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__5891\ : InMux
    port map (
            O => \N__31968\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__5890\ : InMux
    port map (
            O => \N__31965\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__5889\ : InMux
    port map (
            O => \N__31962\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__5888\ : CascadeMux
    port map (
            O => \N__31959\,
            I => \N__31954\
        );

    \I__5887\ : InMux
    port map (
            O => \N__31958\,
            I => \N__31951\
        );

    \I__5886\ : InMux
    port map (
            O => \N__31957\,
            I => \N__31946\
        );

    \I__5885\ : InMux
    port map (
            O => \N__31954\,
            I => \N__31946\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__31951\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__31946\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__5882\ : InMux
    port map (
            O => \N__31941\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31938\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__5880\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31930\
        );

    \I__5879\ : InMux
    port map (
            O => \N__31934\,
            I => \N__31925\
        );

    \I__5878\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31925\
        );

    \I__5877\ : LocalMux
    port map (
            O => \N__31930\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__31925\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__5875\ : CascadeMux
    port map (
            O => \N__31920\,
            I => \N__31915\
        );

    \I__5874\ : InMux
    port map (
            O => \N__31919\,
            I => \N__31912\
        );

    \I__5873\ : InMux
    port map (
            O => \N__31918\,
            I => \N__31909\
        );

    \I__5872\ : InMux
    port map (
            O => \N__31915\,
            I => \N__31906\
        );

    \I__5871\ : LocalMux
    port map (
            O => \N__31912\,
            I => \current_shift_inst.N_1263_i\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__31909\,
            I => \current_shift_inst.N_1263_i\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__31906\,
            I => \current_shift_inst.N_1263_i\
        );

    \I__5868\ : InMux
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__31896\,
            I => \N__31893\
        );

    \I__5866\ : Odrv4
    port map (
            O => \N__31893\,
            I => \current_shift_inst.control_input_1\
        );

    \I__5865\ : InMux
    port map (
            O => \N__31890\,
            I => \bfn_11_10_0_\
        );

    \I__5864\ : CascadeMux
    port map (
            O => \N__31887\,
            I => \N__31883\
        );

    \I__5863\ : InMux
    port map (
            O => \N__31886\,
            I => \N__31877\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31877\
        );

    \I__5861\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31874\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__31877\,
            I => \N__31871\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__31874\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__31871\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31866\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__5856\ : InMux
    port map (
            O => \N__31863\,
            I => \N__31856\
        );

    \I__5855\ : InMux
    port map (
            O => \N__31862\,
            I => \N__31856\
        );

    \I__5854\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31853\
        );

    \I__5853\ : LocalMux
    port map (
            O => \N__31856\,
            I => \N__31850\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__31853\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5851\ : Odrv4
    port map (
            O => \N__31850\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__5850\ : InMux
    port map (
            O => \N__31845\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__5849\ : InMux
    port map (
            O => \N__31842\,
            I => \N__31835\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31841\,
            I => \N__31835\
        );

    \I__5847\ : InMux
    port map (
            O => \N__31840\,
            I => \N__31832\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__31835\,
            I => \N__31829\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31832\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5844\ : Odrv4
    port map (
            O => \N__31829\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__5843\ : InMux
    port map (
            O => \N__31824\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__5842\ : CascadeMux
    port map (
            O => \N__31821\,
            I => \N__31817\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31820\,
            I => \N__31811\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31817\,
            I => \N__31811\
        );

    \I__5839\ : InMux
    port map (
            O => \N__31816\,
            I => \N__31808\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31811\,
            I => \N__31805\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__31808\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5836\ : Odrv4
    port map (
            O => \N__31805\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31800\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__5834\ : CascadeMux
    port map (
            O => \N__31797\,
            I => \N__31793\
        );

    \I__5833\ : InMux
    port map (
            O => \N__31796\,
            I => \N__31787\
        );

    \I__5832\ : InMux
    port map (
            O => \N__31793\,
            I => \N__31787\
        );

    \I__5831\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31784\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31787\,
            I => \N__31781\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31784\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__5828\ : Odrv12
    port map (
            O => \N__31781\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__5827\ : InMux
    port map (
            O => \N__31776\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__5826\ : InMux
    port map (
            O => \N__31773\,
            I => \N__31766\
        );

    \I__5825\ : InMux
    port map (
            O => \N__31772\,
            I => \N__31766\
        );

    \I__5824\ : InMux
    port map (
            O => \N__31771\,
            I => \N__31763\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31766\,
            I => \N__31760\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__31763\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5821\ : Odrv12
    port map (
            O => \N__31760\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__5820\ : InMux
    port map (
            O => \N__31755\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__5819\ : InMux
    port map (
            O => \N__31752\,
            I => \N__31746\
        );

    \I__5818\ : InMux
    port map (
            O => \N__31751\,
            I => \N__31746\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31746\,
            I => \N__31742\
        );

    \I__5816\ : InMux
    port map (
            O => \N__31745\,
            I => \N__31739\
        );

    \I__5815\ : Span4Mux_h
    port map (
            O => \N__31742\,
            I => \N__31736\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__31739\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5813\ : Odrv4
    port map (
            O => \N__31736\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__5812\ : InMux
    port map (
            O => \N__31731\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__5811\ : CascadeMux
    port map (
            O => \N__31728\,
            I => \N__31724\
        );

    \I__5810\ : InMux
    port map (
            O => \N__31727\,
            I => \N__31719\
        );

    \I__5809\ : InMux
    port map (
            O => \N__31724\,
            I => \N__31719\
        );

    \I__5808\ : LocalMux
    port map (
            O => \N__31719\,
            I => \N__31715\
        );

    \I__5807\ : InMux
    port map (
            O => \N__31718\,
            I => \N__31712\
        );

    \I__5806\ : Span4Mux_h
    port map (
            O => \N__31715\,
            I => \N__31709\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__31712\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5804\ : Odrv4
    port map (
            O => \N__31709\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__5803\ : InMux
    port map (
            O => \N__31704\,
            I => \bfn_11_11_0_\
        );

    \I__5802\ : InMux
    port map (
            O => \N__31701\,
            I => \N__31697\
        );

    \I__5801\ : InMux
    port map (
            O => \N__31700\,
            I => \N__31694\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__31697\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__31694\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__5798\ : InMux
    port map (
            O => \N__31689\,
            I => \bfn_11_9_0_\
        );

    \I__5797\ : InMux
    port map (
            O => \N__31686\,
            I => \N__31682\
        );

    \I__5796\ : InMux
    port map (
            O => \N__31685\,
            I => \N__31679\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__31682\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31679\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__5793\ : InMux
    port map (
            O => \N__31674\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__5792\ : InMux
    port map (
            O => \N__31671\,
            I => \N__31667\
        );

    \I__5791\ : InMux
    port map (
            O => \N__31670\,
            I => \N__31664\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__31667\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__5789\ : LocalMux
    port map (
            O => \N__31664\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__5788\ : InMux
    port map (
            O => \N__31659\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__5787\ : InMux
    port map (
            O => \N__31656\,
            I => \N__31652\
        );

    \I__5786\ : InMux
    port map (
            O => \N__31655\,
            I => \N__31649\
        );

    \I__5785\ : LocalMux
    port map (
            O => \N__31652\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__31649\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__5783\ : InMux
    port map (
            O => \N__31644\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__5782\ : InMux
    port map (
            O => \N__31641\,
            I => \N__31637\
        );

    \I__5781\ : InMux
    port map (
            O => \N__31640\,
            I => \N__31634\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31637\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__31634\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__5778\ : InMux
    port map (
            O => \N__31629\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__5777\ : InMux
    port map (
            O => \N__31626\,
            I => \N__31622\
        );

    \I__5776\ : InMux
    port map (
            O => \N__31625\,
            I => \N__31619\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__31622\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__31619\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__5773\ : InMux
    port map (
            O => \N__31614\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__5772\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31607\
        );

    \I__5771\ : InMux
    port map (
            O => \N__31610\,
            I => \N__31604\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__31607\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__31604\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__5768\ : InMux
    port map (
            O => \N__31599\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__5767\ : InMux
    port map (
            O => \N__31596\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__5766\ : InMux
    port map (
            O => \N__31593\,
            I => \N__31588\
        );

    \I__5765\ : InMux
    port map (
            O => \N__31592\,
            I => \N__31583\
        );

    \I__5764\ : InMux
    port map (
            O => \N__31591\,
            I => \N__31583\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__31588\,
            I => \N__31580\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__31583\,
            I => \N__31577\
        );

    \I__5761\ : Span4Mux_v
    port map (
            O => \N__31580\,
            I => \N__31571\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__31577\,
            I => \N__31571\
        );

    \I__5759\ : InMux
    port map (
            O => \N__31576\,
            I => \N__31568\
        );

    \I__5758\ : Span4Mux_h
    port map (
            O => \N__31571\,
            I => \N__31563\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__31568\,
            I => \N__31563\
        );

    \I__5756\ : Odrv4
    port map (
            O => \N__31563\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\
        );

    \I__5755\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31556\
        );

    \I__5754\ : InMux
    port map (
            O => \N__31559\,
            I => \N__31553\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__31556\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__31553\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__5750\ : InMux
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__31542\,
            I => \N__31539\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__31539\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\
        );

    \I__5747\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31532\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31535\,
            I => \N__31529\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__31532\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__31529\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__5743\ : InMux
    port map (
            O => \N__31524\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__5742\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31517\
        );

    \I__5741\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31514\
        );

    \I__5740\ : LocalMux
    port map (
            O => \N__31517\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__31514\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__5738\ : InMux
    port map (
            O => \N__31509\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__5737\ : InMux
    port map (
            O => \N__31506\,
            I => \N__31502\
        );

    \I__5736\ : InMux
    port map (
            O => \N__31505\,
            I => \N__31499\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__31502\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__31499\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31494\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__5732\ : InMux
    port map (
            O => \N__31491\,
            I => \N__31487\
        );

    \I__5731\ : InMux
    port map (
            O => \N__31490\,
            I => \N__31484\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31487\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__31484\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__5728\ : InMux
    port map (
            O => \N__31479\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__5727\ : InMux
    port map (
            O => \N__31476\,
            I => \N__31472\
        );

    \I__5726\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31469\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31472\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__31469\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__5723\ : InMux
    port map (
            O => \N__31464\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__5722\ : InMux
    port map (
            O => \N__31461\,
            I => \N__31457\
        );

    \I__5721\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31454\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__31457\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__31454\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__5718\ : InMux
    port map (
            O => \N__31449\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__5717\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31442\
        );

    \I__5716\ : InMux
    port map (
            O => \N__31445\,
            I => \N__31439\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__31442\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__31439\,
            I => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__5713\ : InMux
    port map (
            O => \N__31434\,
            I => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__5712\ : InMux
    port map (
            O => \N__31431\,
            I => \N__31427\
        );

    \I__5711\ : InMux
    port map (
            O => \N__31430\,
            I => \N__31424\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__31427\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__31424\,
            I => \phase_controller_inst1.stoper_tr.runningZ0\
        );

    \I__5708\ : InMux
    port map (
            O => \N__31419\,
            I => \N__31415\
        );

    \I__5707\ : InMux
    port map (
            O => \N__31418\,
            I => \N__31411\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__31415\,
            I => \N__31408\
        );

    \I__5705\ : InMux
    port map (
            O => \N__31414\,
            I => \N__31405\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__31411\,
            I => \N__31402\
        );

    \I__5703\ : Span4Mux_s2_v
    port map (
            O => \N__31408\,
            I => \N__31397\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__31405\,
            I => \N__31397\
        );

    \I__5701\ : Span4Mux_h
    port map (
            O => \N__31402\,
            I => \N__31392\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__31397\,
            I => \N__31392\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__31392\,
            I => \N__31388\
        );

    \I__5698\ : InMux
    port map (
            O => \N__31391\,
            I => \N__31385\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__31388\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__31385\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\
        );

    \I__5695\ : InMux
    port map (
            O => \N__31380\,
            I => \N__31377\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__31377\,
            I => \N__31372\
        );

    \I__5693\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31369\
        );

    \I__5692\ : InMux
    port map (
            O => \N__31375\,
            I => \N__31366\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__31372\,
            I => \N__31361\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__31369\,
            I => \N__31361\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__31366\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__5688\ : Odrv4
    port map (
            O => \N__31361\,
            I => \elapsed_time_ns_1_RNIFE91B_0_3\
        );

    \I__5687\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31352\
        );

    \I__5686\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31349\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__31352\,
            I => \N__31345\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__31349\,
            I => \N__31342\
        );

    \I__5683\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31339\
        );

    \I__5682\ : Span4Mux_h
    port map (
            O => \N__31345\,
            I => \N__31333\
        );

    \I__5681\ : Span4Mux_h
    port map (
            O => \N__31342\,
            I => \N__31333\
        );

    \I__5680\ : LocalMux
    port map (
            O => \N__31339\,
            I => \N__31330\
        );

    \I__5679\ : InMux
    port map (
            O => \N__31338\,
            I => \N__31327\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__31333\,
            I => \N__31324\
        );

    \I__5677\ : Span4Mux_v
    port map (
            O => \N__31330\,
            I => \N__31321\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__31327\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5675\ : Odrv4
    port map (
            O => \N__31324\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5674\ : Odrv4
    port map (
            O => \N__31321\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\
        );

    \I__5673\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31308\
        );

    \I__5671\ : Span4Mux_h
    port map (
            O => \N__31308\,
            I => \N__31303\
        );

    \I__5670\ : InMux
    port map (
            O => \N__31307\,
            I => \N__31300\
        );

    \I__5669\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31297\
        );

    \I__5668\ : Span4Mux_v
    port map (
            O => \N__31303\,
            I => \N__31294\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31300\,
            I => \N__31291\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__31297\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__31294\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__5664\ : Odrv12
    port map (
            O => \N__31291\,
            I => \elapsed_time_ns_1_RNI5FOBB_0_18\
        );

    \I__5663\ : CascadeMux
    port map (
            O => \N__31284\,
            I => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\
        );

    \I__5662\ : InMux
    port map (
            O => \N__31281\,
            I => \N__31278\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__31278\,
            I => \N__31275\
        );

    \I__5660\ : Span4Mux_s1_v
    port map (
            O => \N__31275\,
            I => \N__31272\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__31272\,
            I => \N__31269\
        );

    \I__5658\ : Odrv4
    port map (
            O => \N__31269\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\
        );

    \I__5657\ : CEMux
    port map (
            O => \N__31266\,
            I => \N__31260\
        );

    \I__5656\ : CEMux
    port map (
            O => \N__31265\,
            I => \N__31257\
        );

    \I__5655\ : CEMux
    port map (
            O => \N__31264\,
            I => \N__31251\
        );

    \I__5654\ : CEMux
    port map (
            O => \N__31263\,
            I => \N__31245\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__31260\,
            I => \N__31240\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__31257\,
            I => \N__31240\
        );

    \I__5651\ : CEMux
    port map (
            O => \N__31256\,
            I => \N__31220\
        );

    \I__5650\ : CEMux
    port map (
            O => \N__31255\,
            I => \N__31208\
        );

    \I__5649\ : CEMux
    port map (
            O => \N__31254\,
            I => \N__31205\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31202\
        );

    \I__5647\ : CEMux
    port map (
            O => \N__31250\,
            I => \N__31196\
        );

    \I__5646\ : CEMux
    port map (
            O => \N__31249\,
            I => \N__31193\
        );

    \I__5645\ : CEMux
    port map (
            O => \N__31248\,
            I => \N__31190\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__31245\,
            I => \N__31185\
        );

    \I__5643\ : Span4Mux_h
    port map (
            O => \N__31240\,
            I => \N__31185\
        );

    \I__5642\ : InMux
    port map (
            O => \N__31239\,
            I => \N__31178\
        );

    \I__5641\ : InMux
    port map (
            O => \N__31238\,
            I => \N__31178\
        );

    \I__5640\ : InMux
    port map (
            O => \N__31237\,
            I => \N__31178\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31236\,
            I => \N__31169\
        );

    \I__5638\ : InMux
    port map (
            O => \N__31235\,
            I => \N__31169\
        );

    \I__5637\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31169\
        );

    \I__5636\ : InMux
    port map (
            O => \N__31233\,
            I => \N__31169\
        );

    \I__5635\ : InMux
    port map (
            O => \N__31232\,
            I => \N__31166\
        );

    \I__5634\ : InMux
    port map (
            O => \N__31231\,
            I => \N__31157\
        );

    \I__5633\ : InMux
    port map (
            O => \N__31230\,
            I => \N__31157\
        );

    \I__5632\ : InMux
    port map (
            O => \N__31229\,
            I => \N__31157\
        );

    \I__5631\ : InMux
    port map (
            O => \N__31228\,
            I => \N__31157\
        );

    \I__5630\ : InMux
    port map (
            O => \N__31227\,
            I => \N__31148\
        );

    \I__5629\ : InMux
    port map (
            O => \N__31226\,
            I => \N__31148\
        );

    \I__5628\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31148\
        );

    \I__5627\ : InMux
    port map (
            O => \N__31224\,
            I => \N__31148\
        );

    \I__5626\ : CEMux
    port map (
            O => \N__31223\,
            I => \N__31145\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__31220\,
            I => \N__31142\
        );

    \I__5624\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31133\
        );

    \I__5623\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31133\
        );

    \I__5622\ : InMux
    port map (
            O => \N__31217\,
            I => \N__31133\
        );

    \I__5621\ : InMux
    port map (
            O => \N__31216\,
            I => \N__31133\
        );

    \I__5620\ : InMux
    port map (
            O => \N__31215\,
            I => \N__31124\
        );

    \I__5619\ : InMux
    port map (
            O => \N__31214\,
            I => \N__31124\
        );

    \I__5618\ : InMux
    port map (
            O => \N__31213\,
            I => \N__31124\
        );

    \I__5617\ : InMux
    port map (
            O => \N__31212\,
            I => \N__31124\
        );

    \I__5616\ : CEMux
    port map (
            O => \N__31211\,
            I => \N__31114\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__31208\,
            I => \N__31109\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__31205\,
            I => \N__31109\
        );

    \I__5613\ : Span4Mux_h
    port map (
            O => \N__31202\,
            I => \N__31106\
        );

    \I__5612\ : CEMux
    port map (
            O => \N__31201\,
            I => \N__31103\
        );

    \I__5611\ : CEMux
    port map (
            O => \N__31200\,
            I => \N__31100\
        );

    \I__5610\ : CEMux
    port map (
            O => \N__31199\,
            I => \N__31097\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__31196\,
            I => \N__31092\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__31193\,
            I => \N__31092\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__31190\,
            I => \N__31083\
        );

    \I__5606\ : Span4Mux_v
    port map (
            O => \N__31185\,
            I => \N__31083\
        );

    \I__5605\ : LocalMux
    port map (
            O => \N__31178\,
            I => \N__31083\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__31169\,
            I => \N__31083\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31166\,
            I => \N__31080\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__31157\,
            I => \N__31075\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__31148\,
            I => \N__31075\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__31145\,
            I => \N__31068\
        );

    \I__5599\ : Span4Mux_s3_v
    port map (
            O => \N__31142\,
            I => \N__31068\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__31133\,
            I => \N__31068\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__31124\,
            I => \N__31065\
        );

    \I__5596\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31058\
        );

    \I__5595\ : InMux
    port map (
            O => \N__31122\,
            I => \N__31058\
        );

    \I__5594\ : InMux
    port map (
            O => \N__31121\,
            I => \N__31058\
        );

    \I__5593\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31049\
        );

    \I__5592\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31049\
        );

    \I__5591\ : InMux
    port map (
            O => \N__31118\,
            I => \N__31049\
        );

    \I__5590\ : InMux
    port map (
            O => \N__31117\,
            I => \N__31049\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__31114\,
            I => \N__31038\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__31109\,
            I => \N__31038\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__31106\,
            I => \N__31038\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__31103\,
            I => \N__31038\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__31100\,
            I => \N__31038\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31097\,
            I => \N__31031\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__31092\,
            I => \N__31031\
        );

    \I__5582\ : Span4Mux_h
    port map (
            O => \N__31083\,
            I => \N__31031\
        );

    \I__5581\ : Span4Mux_h
    port map (
            O => \N__31080\,
            I => \N__31026\
        );

    \I__5580\ : Span4Mux_h
    port map (
            O => \N__31075\,
            I => \N__31026\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__31068\,
            I => \N__31021\
        );

    \I__5578\ : Span4Mux_h
    port map (
            O => \N__31065\,
            I => \N__31021\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__31058\,
            I => \N__31014\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__31049\,
            I => \N__31014\
        );

    \I__5575\ : Span4Mux_v
    port map (
            O => \N__31038\,
            I => \N__31014\
        );

    \I__5574\ : Odrv4
    port map (
            O => \N__31031\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__31026\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__5572\ : Odrv4
    port map (
            O => \N__31021\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__31014\,
            I => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\
        );

    \I__5570\ : InMux
    port map (
            O => \N__31005\,
            I => \N__31001\
        );

    \I__5569\ : InMux
    port map (
            O => \N__31004\,
            I => \N__30997\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__31001\,
            I => \N__30994\
        );

    \I__5567\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30991\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__30997\,
            I => \N__30988\
        );

    \I__5565\ : Span4Mux_h
    port map (
            O => \N__30994\,
            I => \N__30985\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__30991\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__5563\ : Odrv4
    port map (
            O => \N__30988\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__5562\ : Odrv4
    port map (
            O => \N__30985\,
            I => \elapsed_time_ns_1_RNIKJ91B_0_8\
        );

    \I__5561\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30974\
        );

    \I__5560\ : InMux
    port map (
            O => \N__30977\,
            I => \N__30971\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__30974\,
            I => \N__30967\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__30971\,
            I => \N__30964\
        );

    \I__5557\ : InMux
    port map (
            O => \N__30970\,
            I => \N__30961\
        );

    \I__5556\ : Span4Mux_h
    port map (
            O => \N__30967\,
            I => \N__30953\
        );

    \I__5555\ : Span4Mux_v
    port map (
            O => \N__30964\,
            I => \N__30953\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__30961\,
            I => \N__30953\
        );

    \I__5553\ : InMux
    port map (
            O => \N__30960\,
            I => \N__30950\
        );

    \I__5552\ : Odrv4
    port map (
            O => \N__30953\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__30950\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30945\,
            I => \N__30942\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__30942\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\
        );

    \I__5548\ : CascadeMux
    port map (
            O => \N__30939\,
            I => \N__30935\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30938\,
            I => \N__30930\
        );

    \I__5546\ : InMux
    port map (
            O => \N__30935\,
            I => \N__30930\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__30930\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\
        );

    \I__5544\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30924\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__30924\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt30\
        );

    \I__5542\ : InMux
    port map (
            O => \N__30921\,
            I => \N__30917\
        );

    \I__5541\ : InMux
    port map (
            O => \N__30920\,
            I => \N__30913\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__30917\,
            I => \N__30910\
        );

    \I__5539\ : InMux
    port map (
            O => \N__30916\,
            I => \N__30907\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__30913\,
            I => \N__30904\
        );

    \I__5537\ : Span4Mux_h
    port map (
            O => \N__30910\,
            I => \N__30901\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__30907\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__5535\ : Odrv12
    port map (
            O => \N__30904\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__5534\ : Odrv4
    port map (
            O => \N__30901\,
            I => \elapsed_time_ns_1_RNIVAQBB_0_30\
        );

    \I__5533\ : InMux
    port map (
            O => \N__30894\,
            I => \N__30890\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30893\,
            I => \N__30886\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__30890\,
            I => \N__30882\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30889\,
            I => \N__30879\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__30886\,
            I => \N__30876\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30873\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__30882\,
            I => \N__30868\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__30879\,
            I => \N__30868\
        );

    \I__5525\ : Sp12to4
    port map (
            O => \N__30876\,
            I => \N__30863\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30873\,
            I => \N__30863\
        );

    \I__5523\ : Odrv4
    port map (
            O => \N__30868\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__5522\ : Odrv12
    port map (
            O => \N__30863\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\
        );

    \I__5521\ : InMux
    port map (
            O => \N__30858\,
            I => \N__30852\
        );

    \I__5520\ : InMux
    port map (
            O => \N__30857\,
            I => \N__30852\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__30852\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\
        );

    \I__5518\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \N__30846\
        );

    \I__5517\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30843\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__30843\,
            I => \N__30840\
        );

    \I__5515\ : Odrv12
    port map (
            O => \N__30840\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt18\
        );

    \I__5514\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30831\
        );

    \I__5513\ : InMux
    port map (
            O => \N__30836\,
            I => \N__30831\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30831\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\
        );

    \I__5511\ : CascadeMux
    port map (
            O => \N__30828\,
            I => \N__30825\
        );

    \I__5510\ : InMux
    port map (
            O => \N__30825\,
            I => \N__30819\
        );

    \I__5509\ : InMux
    port map (
            O => \N__30824\,
            I => \N__30819\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__30819\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\
        );

    \I__5507\ : InMux
    port map (
            O => \N__30816\,
            I => \N__30813\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__5505\ : Odrv4
    port map (
            O => \N__30810\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\
        );

    \I__5504\ : InMux
    port map (
            O => \N__30807\,
            I => \N__30804\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30800\
        );

    \I__5502\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30797\
        );

    \I__5501\ : Span4Mux_v
    port map (
            O => \N__30800\,
            I => \N__30794\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__30797\,
            I => \N__30791\
        );

    \I__5499\ : Sp12to4
    port map (
            O => \N__30794\,
            I => \N__30788\
        );

    \I__5498\ : Span12Mux_v
    port map (
            O => \N__30791\,
            I => \N__30785\
        );

    \I__5497\ : Span12Mux_s10_h
    port map (
            O => \N__30788\,
            I => \N__30782\
        );

    \I__5496\ : Odrv12
    port map (
            O => \N__30785\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5495\ : Odrv12
    port map (
            O => \N__30782\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_0\
        );

    \I__5494\ : InMux
    port map (
            O => \N__30777\,
            I => \N__30774\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30774\,
            I => \N__30770\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30773\,
            I => \N__30766\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__30770\,
            I => \N__30763\
        );

    \I__5490\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30760\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__30766\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__5488\ : Odrv4
    port map (
            O => \N__30763\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__30760\,
            I => \elapsed_time_ns_1_RNI7IPBB_0_29\
        );

    \I__5486\ : InMux
    port map (
            O => \N__30753\,
            I => \N__30748\
        );

    \I__5485\ : InMux
    port map (
            O => \N__30752\,
            I => \N__30745\
        );

    \I__5484\ : InMux
    port map (
            O => \N__30751\,
            I => \N__30741\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__30748\,
            I => \N__30736\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__30745\,
            I => \N__30736\
        );

    \I__5481\ : InMux
    port map (
            O => \N__30744\,
            I => \N__30733\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__30741\,
            I => \N__30730\
        );

    \I__5479\ : Span4Mux_v
    port map (
            O => \N__30736\,
            I => \N__30727\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__30733\,
            I => \N__30724\
        );

    \I__5477\ : Odrv4
    port map (
            O => \N__30730\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__5476\ : Odrv4
    port map (
            O => \N__30727\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__5475\ : Odrv12
    port map (
            O => \N__30724\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__30714\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\
        );

    \I__5472\ : InMux
    port map (
            O => \N__30711\,
            I => \N__30708\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__30708\,
            I => \N__30705\
        );

    \I__5470\ : Span4Mux_v
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__5469\ : Sp12to4
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__5468\ : Span12Mux_h
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__5467\ : Odrv12
    port map (
            O => \N__30696\,
            I => \pwm_generator_inst.un2_threshold_2_1_16\
        );

    \I__5466\ : InMux
    port map (
            O => \N__30693\,
            I => \N__30690\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__30690\,
            I => \N__30687\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__30687\,
            I => \N__30684\
        );

    \I__5463\ : Span4Mux_h
    port map (
            O => \N__30684\,
            I => \N__30681\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__30681\,
            I => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30675\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\
        );

    \I__5459\ : CascadeMux
    port map (
            O => \N__30672\,
            I => \N__30669\
        );

    \I__5458\ : InMux
    port map (
            O => \N__30669\,
            I => \N__30666\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__30666\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt24\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30663\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_30\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__30660\,
            I => \N__30657\
        );

    \I__5454\ : InMux
    port map (
            O => \N__30657\,
            I => \N__30654\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30654\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt26\
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__30651\,
            I => \N__30647\
        );

    \I__5451\ : InMux
    port map (
            O => \N__30650\,
            I => \N__30642\
        );

    \I__5450\ : InMux
    port map (
            O => \N__30647\,
            I => \N__30642\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__30642\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\
        );

    \I__5448\ : InMux
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__30636\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\
        );

    \I__5446\ : InMux
    port map (
            O => \N__30633\,
            I => \N__30628\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30632\,
            I => \N__30625\
        );

    \I__5444\ : InMux
    port map (
            O => \N__30631\,
            I => \N__30622\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__30628\,
            I => \N__30619\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__30625\,
            I => \N__30616\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30622\,
            I => \N__30611\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__30619\,
            I => \N__30611\
        );

    \I__5439\ : Odrv12
    port map (
            O => \N__30616\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__30611\,
            I => \elapsed_time_ns_1_RNI4FPBB_0_26\
        );

    \I__5437\ : InMux
    port map (
            O => \N__30606\,
            I => \N__30601\
        );

    \I__5436\ : CascadeMux
    port map (
            O => \N__30605\,
            I => \N__30598\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30604\,
            I => \N__30594\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__30601\,
            I => \N__30591\
        );

    \I__5433\ : InMux
    port map (
            O => \N__30598\,
            I => \N__30588\
        );

    \I__5432\ : InMux
    port map (
            O => \N__30597\,
            I => \N__30585\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__30594\,
            I => \N__30582\
        );

    \I__5430\ : Span4Mux_v
    port map (
            O => \N__30591\,
            I => \N__30579\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__30588\,
            I => \N__30576\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30585\,
            I => \N__30573\
        );

    \I__5427\ : Span4Mux_h
    port map (
            O => \N__30582\,
            I => \N__30566\
        );

    \I__5426\ : Span4Mux_v
    port map (
            O => \N__30579\,
            I => \N__30566\
        );

    \I__5425\ : Span4Mux_v
    port map (
            O => \N__30576\,
            I => \N__30566\
        );

    \I__5424\ : Odrv12
    port map (
            O => \N__30573\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5423\ : Odrv4
    port map (
            O => \N__30566\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\
        );

    \I__5422\ : InMux
    port map (
            O => \N__30561\,
            I => \N__30555\
        );

    \I__5421\ : InMux
    port map (
            O => \N__30560\,
            I => \N__30555\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__30555\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\
        );

    \I__5419\ : CascadeMux
    port map (
            O => \N__30552\,
            I => \N__30549\
        );

    \I__5418\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30546\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__30546\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\
        );

    \I__5416\ : CascadeMux
    port map (
            O => \N__30543\,
            I => \N__30540\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30540\,
            I => \N__30537\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__30537\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\
        );

    \I__5413\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30531\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__30531\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__30525\,
            I => \N__30522\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__30522\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\
        );

    \I__5408\ : CascadeMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__5407\ : InMux
    port map (
            O => \N__30516\,
            I => \N__30513\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__30513\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30510\,
            I => \N__30507\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30507\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\
        );

    \I__5403\ : InMux
    port map (
            O => \N__30504\,
            I => \N__30501\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__30501\,
            I => \N__30498\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__30498\,
            I => \N__30495\
        );

    \I__5400\ : Span4Mux_h
    port map (
            O => \N__30495\,
            I => \N__30492\
        );

    \I__5399\ : Odrv4
    port map (
            O => \N__30492\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\
        );

    \I__5398\ : CascadeMux
    port map (
            O => \N__30489\,
            I => \N__30486\
        );

    \I__5397\ : InMux
    port map (
            O => \N__30486\,
            I => \N__30483\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__30483\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\
        );

    \I__5395\ : InMux
    port map (
            O => \N__30480\,
            I => \N__30477\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__30477\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__30474\,
            I => \N__30471\
        );

    \I__5392\ : InMux
    port map (
            O => \N__30471\,
            I => \N__30468\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__30468\,
            I => \N__30465\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__30465\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt20\
        );

    \I__5389\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30459\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__30459\,
            I => \N__30456\
        );

    \I__5387\ : Odrv4
    port map (
            O => \N__30456\,
            I => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__30453\,
            I => \N__30450\
        );

    \I__5385\ : InMux
    port map (
            O => \N__30450\,
            I => \N__30447\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__30447\,
            I => \N__30444\
        );

    \I__5383\ : Odrv4
    port map (
            O => \N__30444\,
            I => \phase_controller_inst2.stoper_tr.un4_running_lt22\
        );

    \I__5382\ : InMux
    port map (
            O => \N__30441\,
            I => \N__30438\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__30438\,
            I => \N__30435\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__30435\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__30432\,
            I => \N__30429\
        );

    \I__5378\ : InMux
    port map (
            O => \N__30429\,
            I => \N__30426\
        );

    \I__5377\ : LocalMux
    port map (
            O => \N__30426\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\
        );

    \I__5376\ : InMux
    port map (
            O => \N__30423\,
            I => \N__30420\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__30420\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__30417\,
            I => \N__30414\
        );

    \I__5373\ : InMux
    port map (
            O => \N__30414\,
            I => \N__30411\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__30411\,
            I => \N__30408\
        );

    \I__5371\ : Odrv4
    port map (
            O => \N__30408\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\
        );

    \I__5370\ : InMux
    port map (
            O => \N__30405\,
            I => \N__30402\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30402\,
            I => \N__30399\
        );

    \I__5368\ : Odrv4
    port map (
            O => \N__30399\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\
        );

    \I__5367\ : CascadeMux
    port map (
            O => \N__30396\,
            I => \N__30393\
        );

    \I__5366\ : InMux
    port map (
            O => \N__30393\,
            I => \N__30390\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__30390\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\
        );

    \I__5364\ : InMux
    port map (
            O => \N__30387\,
            I => \N__30384\
        );

    \I__5363\ : LocalMux
    port map (
            O => \N__30384\,
            I => \N__30381\
        );

    \I__5362\ : Span4Mux_v
    port map (
            O => \N__30381\,
            I => \N__30378\
        );

    \I__5361\ : Odrv4
    port map (
            O => \N__30378\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__30375\,
            I => \N__30372\
        );

    \I__5359\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30369\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__30369\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__30366\,
            I => \N__30363\
        );

    \I__5356\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__30360\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\
        );

    \I__5354\ : InMux
    port map (
            O => \N__30357\,
            I => \N__30354\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__5352\ : Odrv4
    port map (
            O => \N__30351\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\
        );

    \I__5351\ : CascadeMux
    port map (
            O => \N__30348\,
            I => \N__30345\
        );

    \I__5350\ : InMux
    port map (
            O => \N__30345\,
            I => \N__30342\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__30342\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30339\,
            I => \N__30336\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__30336\,
            I => \N__30333\
        );

    \I__5346\ : Odrv4
    port map (
            O => \N__30333\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__30330\,
            I => \N__30327\
        );

    \I__5344\ : InMux
    port map (
            O => \N__30327\,
            I => \N__30324\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__30324\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30321\,
            I => \N__30318\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30318\,
            I => \N__30315\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__30315\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\
        );

    \I__5339\ : CascadeMux
    port map (
            O => \N__30312\,
            I => \N__30309\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30309\,
            I => \N__30306\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__30306\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\
        );

    \I__5336\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30300\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__30300\,
            I => \N__30295\
        );

    \I__5334\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30292\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30298\,
            I => \N__30289\
        );

    \I__5332\ : Span4Mux_s3_v
    port map (
            O => \N__30295\,
            I => \N__30284\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__30292\,
            I => \N__30284\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__30289\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__5329\ : Odrv4
    port map (
            O => \N__30284\,
            I => \elapsed_time_ns_1_RNI0AOBB_0_13\
        );

    \I__5328\ : InMux
    port map (
            O => \N__30279\,
            I => \N__30275\
        );

    \I__5327\ : InMux
    port map (
            O => \N__30278\,
            I => \N__30272\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30275\,
            I => \N__30268\
        );

    \I__5325\ : LocalMux
    port map (
            O => \N__30272\,
            I => \N__30265\
        );

    \I__5324\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30261\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__30268\,
            I => \N__30256\
        );

    \I__5322\ : Span4Mux_v
    port map (
            O => \N__30265\,
            I => \N__30256\
        );

    \I__5321\ : CascadeMux
    port map (
            O => \N__30264\,
            I => \N__30253\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__30261\,
            I => \N__30250\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__30256\,
            I => \N__30247\
        );

    \I__5318\ : InMux
    port map (
            O => \N__30253\,
            I => \N__30244\
        );

    \I__5317\ : Span12Mux_h
    port map (
            O => \N__30250\,
            I => \N__30241\
        );

    \I__5316\ : Sp12to4
    port map (
            O => \N__30247\,
            I => \N__30238\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__30244\,
            I => \N__30235\
        );

    \I__5314\ : Odrv12
    port map (
            O => \N__30241\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5313\ : Odrv12
    port map (
            O => \N__30238\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__30235\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\
        );

    \I__5311\ : InMux
    port map (
            O => \N__30228\,
            I => \N__30224\
        );

    \I__5310\ : InMux
    port map (
            O => \N__30227\,
            I => \N__30220\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__30224\,
            I => \N__30217\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30223\,
            I => \N__30214\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__30220\,
            I => \N__30210\
        );

    \I__5306\ : Span4Mux_s2_v
    port map (
            O => \N__30217\,
            I => \N__30205\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__30214\,
            I => \N__30205\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30213\,
            I => \N__30202\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__30210\,
            I => \N__30197\
        );

    \I__5302\ : Span4Mux_v
    port map (
            O => \N__30205\,
            I => \N__30197\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__30202\,
            I => \N__30194\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__30197\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__30194\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\
        );

    \I__5298\ : InMux
    port map (
            O => \N__30189\,
            I => \N__30186\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__30186\,
            I => \N__30181\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30178\
        );

    \I__5295\ : InMux
    port map (
            O => \N__30184\,
            I => \N__30175\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__30181\,
            I => \N__30172\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__30178\,
            I => \N__30169\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__30175\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__5291\ : Odrv4
    port map (
            O => \N__30172\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__30169\,
            I => \elapsed_time_ns_1_RNIHG91B_0_5\
        );

    \I__5289\ : InMux
    port map (
            O => \N__30162\,
            I => \N__30158\
        );

    \I__5288\ : InMux
    port map (
            O => \N__30161\,
            I => \N__30155\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__30158\,
            I => \N__30149\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__30155\,
            I => \N__30149\
        );

    \I__5285\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30146\
        );

    \I__5284\ : Sp12to4
    port map (
            O => \N__30149\,
            I => \N__30140\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__30146\,
            I => \N__30140\
        );

    \I__5282\ : InMux
    port map (
            O => \N__30145\,
            I => \N__30137\
        );

    \I__5281\ : Span12Mux_s10_v
    port map (
            O => \N__30140\,
            I => \N__30134\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30131\
        );

    \I__5279\ : Odrv12
    port map (
            O => \N__30134\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__5278\ : Odrv12
    port map (
            O => \N__30131\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\
        );

    \I__5277\ : InMux
    port map (
            O => \N__30126\,
            I => \N__30122\
        );

    \I__5276\ : InMux
    port map (
            O => \N__30125\,
            I => \N__30118\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__30122\,
            I => \N__30115\
        );

    \I__5274\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30112\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__30118\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__30115\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__30112\,
            I => \elapsed_time_ns_1_RNILK91B_0_9\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30100\
        );

    \I__5269\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30097\
        );

    \I__5268\ : InMux
    port map (
            O => \N__30103\,
            I => \N__30094\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__30100\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__30097\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__30094\,
            I => \elapsed_time_ns_1_RNIT6OBB_0_10\
        );

    \I__5264\ : InMux
    port map (
            O => \N__30087\,
            I => \N__30084\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__30084\,
            I => \N__30080\
        );

    \I__5262\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30077\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__30080\,
            I => \N__30072\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__30077\,
            I => \N__30069\
        );

    \I__5259\ : InMux
    port map (
            O => \N__30076\,
            I => \N__30064\
        );

    \I__5258\ : InMux
    port map (
            O => \N__30075\,
            I => \N__30064\
        );

    \I__5257\ : Span4Mux_v
    port map (
            O => \N__30072\,
            I => \N__30061\
        );

    \I__5256\ : Span4Mux_h
    port map (
            O => \N__30069\,
            I => \N__30058\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__30064\,
            I => \N__30055\
        );

    \I__5254\ : Odrv4
    port map (
            O => \N__30061\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__5253\ : Odrv4
    port map (
            O => \N__30058\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__5252\ : Odrv12
    port map (
            O => \N__30055\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\
        );

    \I__5251\ : CascadeMux
    port map (
            O => \N__30048\,
            I => \N__30045\
        );

    \I__5250\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30042\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__30042\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\
        );

    \I__5248\ : InMux
    port map (
            O => \N__30039\,
            I => \N__30036\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__30036\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__30033\,
            I => \N__30030\
        );

    \I__5245\ : InMux
    port map (
            O => \N__30030\,
            I => \N__30027\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__30027\,
            I => \N__30024\
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__30024\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\
        );

    \I__5242\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30018\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__30018\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\
        );

    \I__5240\ : CascadeMux
    port map (
            O => \N__30015\,
            I => \N__30012\
        );

    \I__5239\ : InMux
    port map (
            O => \N__30012\,
            I => \N__30009\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__30009\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\
        );

    \I__5237\ : InMux
    port map (
            O => \N__30006\,
            I => \N__30003\
        );

    \I__5236\ : LocalMux
    port map (
            O => \N__30003\,
            I => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29997\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__29997\,
            I => \N__29993\
        );

    \I__5233\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29990\
        );

    \I__5232\ : Odrv4
    port map (
            O => \N__29993\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__29990\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\
        );

    \I__5230\ : CascadeMux
    port map (
            O => \N__29985\,
            I => \N__29982\
        );

    \I__5229\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29979\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29976\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__29976\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\
        );

    \I__5226\ : InMux
    port map (
            O => \N__29973\,
            I => \N__29970\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__29970\,
            I => \N__29967\
        );

    \I__5224\ : Span12Mux_s10_h
    port map (
            O => \N__29967\,
            I => \N__29964\
        );

    \I__5223\ : Odrv12
    port map (
            O => \N__29964\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\
        );

    \I__5222\ : InMux
    port map (
            O => \N__29961\,
            I => \N__29958\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29955\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__29955\,
            I => \N__29952\
        );

    \I__5219\ : Odrv4
    port map (
            O => \N__29952\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt16\
        );

    \I__5218\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29943\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29948\,
            I => \N__29943\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__29943\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\
        );

    \I__5215\ : CascadeMux
    port map (
            O => \N__29940\,
            I => \N__29935\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29939\,
            I => \N__29932\
        );

    \I__5213\ : InMux
    port map (
            O => \N__29938\,
            I => \N__29927\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29927\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__29932\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__29927\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\
        );

    \I__5209\ : CascadeMux
    port map (
            O => \N__29922\,
            I => \N__29918\
        );

    \I__5208\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29914\
        );

    \I__5207\ : InMux
    port map (
            O => \N__29918\,
            I => \N__29911\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29917\,
            I => \N__29908\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__29914\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29911\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__29908\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\
        );

    \I__5202\ : CascadeMux
    port map (
            O => \N__29901\,
            I => \N__29898\
        );

    \I__5201\ : InMux
    port map (
            O => \N__29898\,
            I => \N__29895\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__29895\,
            I => \N__29892\
        );

    \I__5199\ : Span4Mux_h
    port map (
            O => \N__29892\,
            I => \N__29889\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__29889\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\
        );

    \I__5197\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29882\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29885\,
            I => \N__29879\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__29882\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__29879\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\
        );

    \I__5193\ : InMux
    port map (
            O => \N__29874\,
            I => \N__29868\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29868\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__29868\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\
        );

    \I__5190\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29862\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__29862\,
            I => \N__29858\
        );

    \I__5188\ : InMux
    port map (
            O => \N__29861\,
            I => \N__29855\
        );

    \I__5187\ : Span4Mux_v
    port map (
            O => \N__29858\,
            I => \N__29852\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29855\,
            I => \N__29849\
        );

    \I__5185\ : Sp12to4
    port map (
            O => \N__29852\,
            I => \N__29844\
        );

    \I__5184\ : Span12Mux_v
    port map (
            O => \N__29849\,
            I => \N__29844\
        );

    \I__5183\ : Odrv12
    port map (
            O => \N__29844\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_29\
        );

    \I__5182\ : InMux
    port map (
            O => \N__29841\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_28\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29831\
        );

    \I__5179\ : InMux
    port map (
            O => \N__29834\,
            I => \N__29828\
        );

    \I__5178\ : Span4Mux_s2_h
    port map (
            O => \N__29831\,
            I => \N__29825\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__29828\,
            I => \N__29822\
        );

    \I__5176\ : Span4Mux_v
    port map (
            O => \N__29825\,
            I => \N__29819\
        );

    \I__5175\ : Span4Mux_v
    port map (
            O => \N__29822\,
            I => \N__29814\
        );

    \I__5174\ : Span4Mux_h
    port map (
            O => \N__29819\,
            I => \N__29814\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__29814\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_30\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29811\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_29\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29808\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_30\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29805\,
            I => \N__29802\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29802\,
            I => \N__29799\
        );

    \I__5168\ : Odrv12
    port map (
            O => \N__29799\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_31\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__5165\ : Odrv12
    port map (
            O => \N__29790\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29779\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29786\,
            I => \N__29768\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29785\,
            I => \N__29768\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29768\
        );

    \I__5160\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29768\
        );

    \I__5159\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29768\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__29779\,
            I => \N__29765\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29759\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__29765\,
            I => \N__29755\
        );

    \I__5155\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29748\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29763\,
            I => \N__29748\
        );

    \I__5153\ : InMux
    port map (
            O => \N__29762\,
            I => \N__29748\
        );

    \I__5152\ : Span4Mux_s3_h
    port map (
            O => \N__29759\,
            I => \N__29745\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29758\,
            I => \N__29742\
        );

    \I__5150\ : Span4Mux_h
    port map (
            O => \N__29755\,
            I => \N__29737\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__29748\,
            I => \N__29737\
        );

    \I__5148\ : Odrv4
    port map (
            O => \N__29745\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__29742\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__5146\ : Odrv4
    port map (
            O => \N__29737\,
            I => \current_shift_inst.PI_CTRL.un8_enablelto31\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29727\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29727\,
            I => \N__29724\
        );

    \I__5143\ : Odrv12
    port map (
            O => \N__29724\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__29721\,
            I => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29718\,
            I => \N__29715\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__29715\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29708\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29711\,
            I => \N__29705\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29708\,
            I => \N__29702\
        );

    \I__5136\ : LocalMux
    port map (
            O => \N__29705\,
            I => \N__29699\
        );

    \I__5135\ : Span12Mux_s9_h
    port map (
            O => \N__29702\,
            I => \N__29696\
        );

    \I__5134\ : Span12Mux_v
    port map (
            O => \N__29699\,
            I => \N__29693\
        );

    \I__5133\ : Odrv12
    port map (
            O => \N__29696\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__5132\ : Odrv12
    port map (
            O => \N__29693\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_21\
        );

    \I__5131\ : InMux
    port map (
            O => \N__29688\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_20\
        );

    \I__5130\ : InMux
    port map (
            O => \N__29685\,
            I => \N__29682\
        );

    \I__5129\ : LocalMux
    port map (
            O => \N__29682\,
            I => \N__29679\
        );

    \I__5128\ : Span4Mux_s2_h
    port map (
            O => \N__29679\,
            I => \N__29675\
        );

    \I__5127\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29672\
        );

    \I__5126\ : Span4Mux_h
    port map (
            O => \N__29675\,
            I => \N__29669\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29672\,
            I => \N__29666\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__29669\,
            I => \N__29663\
        );

    \I__5123\ : Odrv12
    port map (
            O => \N__29666\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__5122\ : Odrv4
    port map (
            O => \N__29663\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_22\
        );

    \I__5121\ : InMux
    port map (
            O => \N__29658\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_21\
        );

    \I__5120\ : InMux
    port map (
            O => \N__29655\,
            I => \N__29651\
        );

    \I__5119\ : InMux
    port map (
            O => \N__29654\,
            I => \N__29648\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__29651\,
            I => \N__29645\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__29648\,
            I => \N__29642\
        );

    \I__5116\ : Span4Mux_v
    port map (
            O => \N__29645\,
            I => \N__29637\
        );

    \I__5115\ : Span4Mux_v
    port map (
            O => \N__29642\,
            I => \N__29637\
        );

    \I__5114\ : Sp12to4
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__29634\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_23\
        );

    \I__5112\ : InMux
    port map (
            O => \N__29631\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_22\
        );

    \I__5111\ : InMux
    port map (
            O => \N__29628\,
            I => \N__29625\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__29625\,
            I => \N__29621\
        );

    \I__5109\ : InMux
    port map (
            O => \N__29624\,
            I => \N__29618\
        );

    \I__5108\ : Span4Mux_h
    port map (
            O => \N__29621\,
            I => \N__29615\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29618\,
            I => \N__29612\
        );

    \I__5106\ : Span4Mux_h
    port map (
            O => \N__29615\,
            I => \N__29609\
        );

    \I__5105\ : Span12Mux_s9_h
    port map (
            O => \N__29612\,
            I => \N__29606\
        );

    \I__5104\ : Odrv4
    port map (
            O => \N__29609\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__5103\ : Odrv12
    port map (
            O => \N__29606\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_24\
        );

    \I__5102\ : InMux
    port map (
            O => \N__29601\,
            I => \bfn_9_16_0_\
        );

    \I__5101\ : InMux
    port map (
            O => \N__29598\,
            I => \N__29595\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__29595\,
            I => \N__29591\
        );

    \I__5099\ : InMux
    port map (
            O => \N__29594\,
            I => \N__29588\
        );

    \I__5098\ : Span4Mux_s1_h
    port map (
            O => \N__29591\,
            I => \N__29585\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__29588\,
            I => \N__29582\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__29585\,
            I => \N__29579\
        );

    \I__5095\ : Span12Mux_v
    port map (
            O => \N__29582\,
            I => \N__29576\
        );

    \I__5094\ : Span4Mux_h
    port map (
            O => \N__29579\,
            I => \N__29573\
        );

    \I__5093\ : Odrv12
    port map (
            O => \N__29576\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__5092\ : Odrv4
    port map (
            O => \N__29573\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_25\
        );

    \I__5091\ : InMux
    port map (
            O => \N__29568\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_24\
        );

    \I__5090\ : InMux
    port map (
            O => \N__29565\,
            I => \N__29561\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29564\,
            I => \N__29558\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__29561\,
            I => \N__29555\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__29558\,
            I => \N__29552\
        );

    \I__5086\ : Span4Mux_s1_h
    port map (
            O => \N__29555\,
            I => \N__29549\
        );

    \I__5085\ : Span4Mux_v
    port map (
            O => \N__29552\,
            I => \N__29546\
        );

    \I__5084\ : Span4Mux_h
    port map (
            O => \N__29549\,
            I => \N__29543\
        );

    \I__5083\ : Span4Mux_h
    port map (
            O => \N__29546\,
            I => \N__29538\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__29543\,
            I => \N__29538\
        );

    \I__5081\ : Odrv4
    port map (
            O => \N__29538\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_26\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29535\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_25\
        );

    \I__5079\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29528\
        );

    \I__5078\ : InMux
    port map (
            O => \N__29531\,
            I => \N__29525\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29528\,
            I => \N__29522\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__29525\,
            I => \N__29519\
        );

    \I__5075\ : Span4Mux_s1_h
    port map (
            O => \N__29522\,
            I => \N__29516\
        );

    \I__5074\ : Span4Mux_v
    port map (
            O => \N__29519\,
            I => \N__29513\
        );

    \I__5073\ : Span4Mux_h
    port map (
            O => \N__29516\,
            I => \N__29510\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__29513\,
            I => \N__29505\
        );

    \I__5071\ : Span4Mux_h
    port map (
            O => \N__29510\,
            I => \N__29505\
        );

    \I__5070\ : Odrv4
    port map (
            O => \N__29505\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_27\
        );

    \I__5069\ : InMux
    port map (
            O => \N__29502\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_26\
        );

    \I__5068\ : InMux
    port map (
            O => \N__29499\,
            I => \N__29496\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29496\,
            I => \N__29493\
        );

    \I__5066\ : Span4Mux_s1_h
    port map (
            O => \N__29493\,
            I => \N__29489\
        );

    \I__5065\ : InMux
    port map (
            O => \N__29492\,
            I => \N__29486\
        );

    \I__5064\ : Span4Mux_h
    port map (
            O => \N__29489\,
            I => \N__29483\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__29486\,
            I => \N__29480\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__29483\,
            I => \N__29477\
        );

    \I__5061\ : Odrv12
    port map (
            O => \N__29480\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__29477\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_28\
        );

    \I__5059\ : InMux
    port map (
            O => \N__29472\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_27\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29469\,
            I => \N__29465\
        );

    \I__5057\ : InMux
    port map (
            O => \N__29468\,
            I => \N__29462\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29465\,
            I => \N__29459\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__29462\,
            I => \N__29456\
        );

    \I__5054\ : Span12Mux_s9_h
    port map (
            O => \N__29459\,
            I => \N__29453\
        );

    \I__5053\ : Odrv12
    port map (
            O => \N__29456\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__5052\ : Odrv12
    port map (
            O => \N__29453\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_13\
        );

    \I__5051\ : InMux
    port map (
            O => \N__29448\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_12\
        );

    \I__5050\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29441\
        );

    \I__5049\ : InMux
    port map (
            O => \N__29444\,
            I => \N__29438\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__29441\,
            I => \N__29435\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__29438\,
            I => \N__29432\
        );

    \I__5046\ : Span4Mux_v
    port map (
            O => \N__29435\,
            I => \N__29429\
        );

    \I__5045\ : Span4Mux_v
    port map (
            O => \N__29432\,
            I => \N__29424\
        );

    \I__5044\ : Span4Mux_v
    port map (
            O => \N__29429\,
            I => \N__29424\
        );

    \I__5043\ : Sp12to4
    port map (
            O => \N__29424\,
            I => \N__29421\
        );

    \I__5042\ : Odrv12
    port map (
            O => \N__29421\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_14\
        );

    \I__5041\ : InMux
    port map (
            O => \N__29418\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_13\
        );

    \I__5040\ : InMux
    port map (
            O => \N__29415\,
            I => \N__29412\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__29412\,
            I => \N__29408\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29411\,
            I => \N__29405\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__29408\,
            I => \N__29402\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__29405\,
            I => \N__29397\
        );

    \I__5035\ : Sp12to4
    port map (
            O => \N__29402\,
            I => \N__29397\
        );

    \I__5034\ : Odrv12
    port map (
            O => \N__29397\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_15\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29394\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_14\
        );

    \I__5032\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29387\
        );

    \I__5031\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29384\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__29387\,
            I => \N__29381\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__29384\,
            I => \N__29378\
        );

    \I__5028\ : Span4Mux_s1_h
    port map (
            O => \N__29381\,
            I => \N__29375\
        );

    \I__5027\ : Span4Mux_v
    port map (
            O => \N__29378\,
            I => \N__29372\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__29375\,
            I => \N__29369\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__29372\,
            I => \N__29364\
        );

    \I__5024\ : Span4Mux_h
    port map (
            O => \N__29369\,
            I => \N__29364\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__29364\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_16\
        );

    \I__5022\ : InMux
    port map (
            O => \N__29361\,
            I => \bfn_9_15_0_\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29358\,
            I => \N__29354\
        );

    \I__5020\ : InMux
    port map (
            O => \N__29357\,
            I => \N__29351\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__29354\,
            I => \N__29348\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29351\,
            I => \N__29345\
        );

    \I__5017\ : Span12Mux_s9_h
    port map (
            O => \N__29348\,
            I => \N__29342\
        );

    \I__5016\ : Odrv12
    port map (
            O => \N__29345\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__5015\ : Odrv12
    port map (
            O => \N__29342\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_17\
        );

    \I__5014\ : InMux
    port map (
            O => \N__29337\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_16\
        );

    \I__5013\ : InMux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__5011\ : Span4Mux_s1_h
    port map (
            O => \N__29328\,
            I => \N__29324\
        );

    \I__5010\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29321\
        );

    \I__5009\ : Span4Mux_h
    port map (
            O => \N__29324\,
            I => \N__29318\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__29321\,
            I => \N__29315\
        );

    \I__5007\ : Span4Mux_h
    port map (
            O => \N__29318\,
            I => \N__29312\
        );

    \I__5006\ : Odrv12
    port map (
            O => \N__29315\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__29312\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_18\
        );

    \I__5004\ : InMux
    port map (
            O => \N__29307\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_17\
        );

    \I__5003\ : InMux
    port map (
            O => \N__29304\,
            I => \N__29300\
        );

    \I__5002\ : InMux
    port map (
            O => \N__29303\,
            I => \N__29297\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__29300\,
            I => \N__29294\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__29297\,
            I => \N__29291\
        );

    \I__4999\ : Span4Mux_s1_h
    port map (
            O => \N__29294\,
            I => \N__29288\
        );

    \I__4998\ : Span4Mux_v
    port map (
            O => \N__29291\,
            I => \N__29285\
        );

    \I__4997\ : Span4Mux_h
    port map (
            O => \N__29288\,
            I => \N__29282\
        );

    \I__4996\ : Span4Mux_h
    port map (
            O => \N__29285\,
            I => \N__29277\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__29282\,
            I => \N__29277\
        );

    \I__4994\ : Odrv4
    port map (
            O => \N__29277\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_19\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29274\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_18\
        );

    \I__4992\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29267\
        );

    \I__4991\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29264\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__29267\,
            I => \N__29261\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29264\,
            I => \N__29258\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__29261\,
            I => \N__29253\
        );

    \I__4987\ : Span4Mux_v
    port map (
            O => \N__29258\,
            I => \N__29253\
        );

    \I__4986\ : Sp12to4
    port map (
            O => \N__29253\,
            I => \N__29250\
        );

    \I__4985\ : Odrv12
    port map (
            O => \N__29250\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_20\
        );

    \I__4984\ : InMux
    port map (
            O => \N__29247\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_19\
        );

    \I__4983\ : InMux
    port map (
            O => \N__29244\,
            I => \N__29240\
        );

    \I__4982\ : InMux
    port map (
            O => \N__29243\,
            I => \N__29237\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__29240\,
            I => \N__29234\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__29237\,
            I => \N__29231\
        );

    \I__4979\ : Span4Mux_v
    port map (
            O => \N__29234\,
            I => \N__29228\
        );

    \I__4978\ : Sp12to4
    port map (
            O => \N__29231\,
            I => \N__29225\
        );

    \I__4977\ : Sp12to4
    port map (
            O => \N__29228\,
            I => \N__29220\
        );

    \I__4976\ : Span12Mux_v
    port map (
            O => \N__29225\,
            I => \N__29220\
        );

    \I__4975\ : Odrv12
    port map (
            O => \N__29220\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_4\
        );

    \I__4974\ : InMux
    port map (
            O => \N__29217\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_3\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29214\,
            I => \N__29210\
        );

    \I__4972\ : InMux
    port map (
            O => \N__29213\,
            I => \N__29207\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__29210\,
            I => \N__29204\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__29207\,
            I => \N__29199\
        );

    \I__4969\ : Span12Mux_v
    port map (
            O => \N__29204\,
            I => \N__29199\
        );

    \I__4968\ : Odrv12
    port map (
            O => \N__29199\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_5\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29196\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_4\
        );

    \I__4966\ : InMux
    port map (
            O => \N__29193\,
            I => \N__29189\
        );

    \I__4965\ : InMux
    port map (
            O => \N__29192\,
            I => \N__29186\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__29186\,
            I => \N__29180\
        );

    \I__4962\ : Span12Mux_s9_h
    port map (
            O => \N__29183\,
            I => \N__29177\
        );

    \I__4961\ : Odrv12
    port map (
            O => \N__29180\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__4960\ : Odrv12
    port map (
            O => \N__29177\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_6\
        );

    \I__4959\ : InMux
    port map (
            O => \N__29172\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_5\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29166\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__29166\,
            I => \N__29163\
        );

    \I__4956\ : Span4Mux_v
    port map (
            O => \N__29163\,
            I => \N__29159\
        );

    \I__4955\ : InMux
    port map (
            O => \N__29162\,
            I => \N__29156\
        );

    \I__4954\ : Span4Mux_h
    port map (
            O => \N__29159\,
            I => \N__29153\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__29156\,
            I => \N__29150\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__29153\,
            I => \N__29147\
        );

    \I__4951\ : Odrv12
    port map (
            O => \N__29150\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__29147\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_7\
        );

    \I__4949\ : InMux
    port map (
            O => \N__29142\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_6\
        );

    \I__4948\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29136\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__29136\,
            I => \N__29132\
        );

    \I__4946\ : InMux
    port map (
            O => \N__29135\,
            I => \N__29129\
        );

    \I__4945\ : Span4Mux_v
    port map (
            O => \N__29132\,
            I => \N__29126\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29129\,
            I => \N__29123\
        );

    \I__4943\ : Sp12to4
    port map (
            O => \N__29126\,
            I => \N__29120\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__29123\,
            I => \N__29117\
        );

    \I__4941\ : Span12Mux_s9_h
    port map (
            O => \N__29120\,
            I => \N__29114\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__29117\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__4939\ : Odrv12
    port map (
            O => \N__29114\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_8\
        );

    \I__4938\ : InMux
    port map (
            O => \N__29109\,
            I => \bfn_9_14_0_\
        );

    \I__4937\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29103\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__29103\,
            I => \N__29099\
        );

    \I__4935\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29096\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__29099\,
            I => \N__29093\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29090\
        );

    \I__4932\ : Sp12to4
    port map (
            O => \N__29093\,
            I => \N__29087\
        );

    \I__4931\ : Span12Mux_s4_h
    port map (
            O => \N__29090\,
            I => \N__29082\
        );

    \I__4930\ : Span12Mux_v
    port map (
            O => \N__29087\,
            I => \N__29082\
        );

    \I__4929\ : Odrv12
    port map (
            O => \N__29082\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_9\
        );

    \I__4928\ : InMux
    port map (
            O => \N__29079\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_8\
        );

    \I__4927\ : InMux
    port map (
            O => \N__29076\,
            I => \N__29073\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__29073\,
            I => \N__29069\
        );

    \I__4925\ : InMux
    port map (
            O => \N__29072\,
            I => \N__29066\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__29069\,
            I => \N__29063\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__29066\,
            I => \N__29060\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__29063\,
            I => \N__29057\
        );

    \I__4921\ : Span12Mux_v
    port map (
            O => \N__29060\,
            I => \N__29054\
        );

    \I__4920\ : Span4Mux_h
    port map (
            O => \N__29057\,
            I => \N__29051\
        );

    \I__4919\ : Odrv12
    port map (
            O => \N__29054\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__29051\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_10\
        );

    \I__4917\ : InMux
    port map (
            O => \N__29046\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_9\
        );

    \I__4916\ : InMux
    port map (
            O => \N__29043\,
            I => \N__29040\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__29040\,
            I => \N__29036\
        );

    \I__4914\ : InMux
    port map (
            O => \N__29039\,
            I => \N__29033\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__29036\,
            I => \N__29030\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__29033\,
            I => \N__29027\
        );

    \I__4911\ : Span4Mux_h
    port map (
            O => \N__29030\,
            I => \N__29024\
        );

    \I__4910\ : Span12Mux_s9_h
    port map (
            O => \N__29027\,
            I => \N__29021\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__29024\,
            I => \N__29018\
        );

    \I__4908\ : Odrv12
    port map (
            O => \N__29021\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__4907\ : Odrv4
    port map (
            O => \N__29018\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_11\
        );

    \I__4906\ : InMux
    port map (
            O => \N__29013\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_10\
        );

    \I__4905\ : InMux
    port map (
            O => \N__29010\,
            I => \N__29006\
        );

    \I__4904\ : InMux
    port map (
            O => \N__29009\,
            I => \N__29003\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__29006\,
            I => \N__29000\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__29003\,
            I => \N__28997\
        );

    \I__4901\ : Span4Mux_v
    port map (
            O => \N__29000\,
            I => \N__28994\
        );

    \I__4900\ : Span4Mux_v
    port map (
            O => \N__28997\,
            I => \N__28991\
        );

    \I__4899\ : Span4Mux_h
    port map (
            O => \N__28994\,
            I => \N__28988\
        );

    \I__4898\ : Span4Mux_h
    port map (
            O => \N__28991\,
            I => \N__28985\
        );

    \I__4897\ : Span4Mux_h
    port map (
            O => \N__28988\,
            I => \N__28982\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__28985\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__28982\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_12\
        );

    \I__4894\ : InMux
    port map (
            O => \N__28977\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_11\
        );

    \I__4893\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28970\
        );

    \I__4892\ : InMux
    port map (
            O => \N__28973\,
            I => \N__28967\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__28970\,
            I => \N__28962\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__28967\,
            I => \N__28959\
        );

    \I__4889\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28954\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28954\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__28962\,
            I => \N__28951\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__28959\,
            I => \N__28948\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28945\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__28951\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4883\ : Odrv4
    port map (
            O => \N__28948\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4882\ : Odrv12
    port map (
            O => \N__28945\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\
        );

    \I__4881\ : InMux
    port map (
            O => \N__28938\,
            I => \N__28933\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28937\,
            I => \N__28930\
        );

    \I__4879\ : InMux
    port map (
            O => \N__28936\,
            I => \N__28927\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28924\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__28930\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__28927\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__28924\,
            I => \elapsed_time_ns_1_RNI0CQBB_0_31\
        );

    \I__4874\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28911\
        );

    \I__4873\ : InMux
    port map (
            O => \N__28916\,
            I => \N__28911\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__28911\,
            I => \N__28906\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28903\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28900\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__28906\,
            I => \N__28897\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__28903\,
            I => \N__28894\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__28900\,
            I => \N__28887\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__28897\,
            I => \N__28887\
        );

    \I__4865\ : Span4Mux_h
    port map (
            O => \N__28894\,
            I => \N__28887\
        );

    \I__4864\ : Odrv4
    port map (
            O => \N__28887\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28884\,
            I => \N__28881\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28878\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__28878\,
            I => \N__28874\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28871\
        );

    \I__4859\ : Odrv4
    port map (
            O => \N__28874\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__28871\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27\
        );

    \I__4857\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28861\
        );

    \I__4856\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28858\
        );

    \I__4855\ : InMux
    port map (
            O => \N__28864\,
            I => \N__28855\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__28861\,
            I => \N__28852\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28849\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__28855\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__4851\ : Odrv4
    port map (
            O => \N__28852\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__4850\ : Odrv4
    port map (
            O => \N__28849\,
            I => \elapsed_time_ns_1_RNIV9PBB_0_21\
        );

    \I__4849\ : InMux
    port map (
            O => \N__28842\,
            I => \N__28835\
        );

    \I__4848\ : InMux
    port map (
            O => \N__28841\,
            I => \N__28835\
        );

    \I__4847\ : InMux
    port map (
            O => \N__28840\,
            I => \N__28831\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__28835\,
            I => \N__28828\
        );

    \I__4845\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28825\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__28831\,
            I => \N__28820\
        );

    \I__4843\ : Span4Mux_v
    port map (
            O => \N__28828\,
            I => \N__28820\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__28825\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__28820\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__28815\,
            I => \N__28812\
        );

    \I__4839\ : InMux
    port map (
            O => \N__28812\,
            I => \N__28806\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28811\,
            I => \N__28806\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__28806\,
            I => \N__28803\
        );

    \I__4836\ : Odrv4
    port map (
            O => \N__28803\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\
        );

    \I__4835\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28795\
        );

    \I__4834\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28792\
        );

    \I__4833\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28789\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__28795\,
            I => \N__28786\
        );

    \I__4831\ : LocalMux
    port map (
            O => \N__28792\,
            I => \N__28783\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__28789\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4829\ : Odrv4
    port map (
            O => \N__28786\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__28783\,
            I => \elapsed_time_ns_1_RNI6GOBB_0_19\
        );

    \I__4827\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28772\
        );

    \I__4826\ : CascadeMux
    port map (
            O => \N__28775\,
            I => \N__28769\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28765\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28769\,
            I => \N__28762\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28768\,
            I => \N__28759\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__28765\,
            I => \N__28751\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__28762\,
            I => \N__28751\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__28759\,
            I => \N__28751\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28748\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__28751\,
            I => \N__28745\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__28748\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4816\ : Odrv4
    port map (
            O => \N__28745\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__28737\,
            I => \current_shift_inst.PI_CTRL.error_control_2_axb_0\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28734\,
            I => \N__28730\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28733\,
            I => \N__28727\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__28730\,
            I => \N__28724\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__28727\,
            I => \N__28721\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__28724\,
            I => \N__28718\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__28721\,
            I => \N__28715\
        );

    \I__4807\ : Span4Mux_h
    port map (
            O => \N__28718\,
            I => \N__28712\
        );

    \I__4806\ : Span4Mux_h
    port map (
            O => \N__28715\,
            I => \N__28709\
        );

    \I__4805\ : Span4Mux_v
    port map (
            O => \N__28712\,
            I => \N__28706\
        );

    \I__4804\ : Span4Mux_h
    port map (
            O => \N__28709\,
            I => \N__28703\
        );

    \I__4803\ : Odrv4
    port map (
            O => \N__28706\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__4802\ : Odrv4
    port map (
            O => \N__28703\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_1\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28698\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_0\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28695\,
            I => \N__28692\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__4798\ : Span4Mux_v
    port map (
            O => \N__28689\,
            I => \N__28685\
        );

    \I__4797\ : InMux
    port map (
            O => \N__28688\,
            I => \N__28682\
        );

    \I__4796\ : Span4Mux_h
    port map (
            O => \N__28685\,
            I => \N__28679\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__28682\,
            I => \N__28676\
        );

    \I__4794\ : Span4Mux_h
    port map (
            O => \N__28679\,
            I => \N__28673\
        );

    \I__4793\ : Odrv12
    port map (
            O => \N__28676\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__28673\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_2\
        );

    \I__4791\ : InMux
    port map (
            O => \N__28668\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_1\
        );

    \I__4790\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28661\
        );

    \I__4789\ : InMux
    port map (
            O => \N__28664\,
            I => \N__28658\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__28661\,
            I => \N__28655\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28658\,
            I => \N__28652\
        );

    \I__4786\ : Span4Mux_v
    port map (
            O => \N__28655\,
            I => \N__28649\
        );

    \I__4785\ : Span4Mux_h
    port map (
            O => \N__28652\,
            I => \N__28646\
        );

    \I__4784\ : Span4Mux_h
    port map (
            O => \N__28649\,
            I => \N__28643\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__28646\,
            I => \N__28638\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__28643\,
            I => \N__28638\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__28638\,
            I => \current_shift_inst.PI_CTRL.prop_term_1_3\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28635\,
            I => \current_shift_inst.PI_CTRL.error_control_2_cry_2\
        );

    \I__4779\ : InMux
    port map (
            O => \N__28632\,
            I => \N__28628\
        );

    \I__4778\ : InMux
    port map (
            O => \N__28631\,
            I => \N__28624\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28628\,
            I => \N__28621\
        );

    \I__4776\ : InMux
    port map (
            O => \N__28627\,
            I => \N__28618\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__28624\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4774\ : Odrv12
    port map (
            O => \N__28621\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__28618\,
            I => \elapsed_time_ns_1_RNI2DPBB_0_24\
        );

    \I__4772\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28606\
        );

    \I__4771\ : CascadeMux
    port map (
            O => \N__28610\,
            I => \N__28602\
        );

    \I__4770\ : InMux
    port map (
            O => \N__28609\,
            I => \N__28599\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__28606\,
            I => \N__28596\
        );

    \I__4768\ : InMux
    port map (
            O => \N__28605\,
            I => \N__28593\
        );

    \I__4767\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28590\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28599\,
            I => \N__28587\
        );

    \I__4765\ : Span4Mux_h
    port map (
            O => \N__28596\,
            I => \N__28580\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28580\
        );

    \I__4763\ : LocalMux
    port map (
            O => \N__28590\,
            I => \N__28580\
        );

    \I__4762\ : Span4Mux_h
    port map (
            O => \N__28587\,
            I => \N__28575\
        );

    \I__4761\ : Span4Mux_v
    port map (
            O => \N__28580\,
            I => \N__28575\
        );

    \I__4760\ : Odrv4
    port map (
            O => \N__28575\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28572\,
            I => \N__28566\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28571\,
            I => \N__28566\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__28566\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\
        );

    \I__4756\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28559\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28562\,
            I => \N__28555\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__28559\,
            I => \N__28552\
        );

    \I__4753\ : InMux
    port map (
            O => \N__28558\,
            I => \N__28549\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28555\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__28552\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__28549\,
            I => \elapsed_time_ns_1_RNIV8OBB_0_12\
        );

    \I__4749\ : CascadeMux
    port map (
            O => \N__28542\,
            I => \N__28537\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28541\,
            I => \N__28533\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28540\,
            I => \N__28528\
        );

    \I__4746\ : InMux
    port map (
            O => \N__28537\,
            I => \N__28528\
        );

    \I__4745\ : InMux
    port map (
            O => \N__28536\,
            I => \N__28525\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__28533\,
            I => \N__28520\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__28528\,
            I => \N__28520\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__28525\,
            I => \N__28517\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__28520\,
            I => \N__28514\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__28517\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__28514\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\
        );

    \I__4738\ : InMux
    port map (
            O => \N__28509\,
            I => \N__28505\
        );

    \I__4737\ : InMux
    port map (
            O => \N__28508\,
            I => \N__28501\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__28505\,
            I => \N__28498\
        );

    \I__4735\ : InMux
    port map (
            O => \N__28504\,
            I => \N__28495\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__28501\,
            I => \N__28492\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__28498\,
            I => \N__28489\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__28495\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__28492\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__28489\,
            I => \elapsed_time_ns_1_RNIED91B_0_2\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28478\
        );

    \I__4728\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28474\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__28478\,
            I => \N__28471\
        );

    \I__4726\ : CascadeMux
    port map (
            O => \N__28477\,
            I => \N__28467\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28474\,
            I => \N__28464\
        );

    \I__4724\ : Span4Mux_h
    port map (
            O => \N__28471\,
            I => \N__28461\
        );

    \I__4723\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28458\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28467\,
            I => \N__28455\
        );

    \I__4721\ : Odrv12
    port map (
            O => \N__28464\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__28461\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__28458\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__28455\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\
        );

    \I__4717\ : InMux
    port map (
            O => \N__28446\,
            I => \N__28440\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28445\,
            I => \N__28440\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__28440\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\
        );

    \I__4714\ : InMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__28434\,
            I => \N__28431\
        );

    \I__4712\ : Span4Mux_s1_v
    port map (
            O => \N__28431\,
            I => \N__28427\
        );

    \I__4711\ : InMux
    port map (
            O => \N__28430\,
            I => \N__28424\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__28427\,
            I => \N__28419\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__28424\,
            I => \N__28416\
        );

    \I__4708\ : InMux
    port map (
            O => \N__28423\,
            I => \N__28413\
        );

    \I__4707\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28410\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__28419\,
            I => \N__28407\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__28416\,
            I => \N__28402\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28413\,
            I => \N__28402\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__28410\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__28407\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4701\ : Odrv4
    port map (
            O => \N__28402\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28395\,
            I => \N__28390\
        );

    \I__4699\ : InMux
    port map (
            O => \N__28394\,
            I => \N__28387\
        );

    \I__4698\ : InMux
    port map (
            O => \N__28393\,
            I => \N__28384\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__28390\,
            I => \N__28381\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__28387\,
            I => \N__28378\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__28384\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4694\ : Odrv12
    port map (
            O => \N__28381\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__28378\,
            I => \elapsed_time_ns_1_RNIIH91B_0_6\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__4690\ : Span4Mux_v
    port map (
            O => \N__28365\,
            I => \N__28359\
        );

    \I__4689\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28356\
        );

    \I__4688\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28351\
        );

    \I__4687\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28351\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__28359\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__28356\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__28351\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28344\,
            I => \N__28340\
        );

    \I__4682\ : InMux
    port map (
            O => \N__28343\,
            I => \N__28336\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28333\
        );

    \I__4680\ : InMux
    port map (
            O => \N__28339\,
            I => \N__28330\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__28336\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4678\ : Odrv12
    port map (
            O => \N__28333\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__28330\,
            I => \elapsed_time_ns_1_RNIGF91B_0_4\
        );

    \I__4676\ : CascadeMux
    port map (
            O => \N__28323\,
            I => \N__28320\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28320\,
            I => \N__28314\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28319\,
            I => \N__28314\
        );

    \I__4673\ : LocalMux
    port map (
            O => \N__28314\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\
        );

    \I__4672\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__28308\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\
        );

    \I__4670\ : InMux
    port map (
            O => \N__28305\,
            I => \N__28302\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__28302\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__28299\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_\
        );

    \I__4667\ : InMux
    port map (
            O => \N__28296\,
            I => \N__28293\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__28293\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\
        );

    \I__4665\ : InMux
    port map (
            O => \N__28290\,
            I => \N__28287\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__28287\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\
        );

    \I__4663\ : CascadeMux
    port map (
            O => \N__28284\,
            I => \N__28281\
        );

    \I__4662\ : InMux
    port map (
            O => \N__28281\,
            I => \N__28275\
        );

    \I__4661\ : InMux
    port map (
            O => \N__28280\,
            I => \N__28275\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__28275\,
            I => \N__28272\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__28272\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__4657\ : InMux
    port map (
            O => \N__28266\,
            I => \N__28259\
        );

    \I__4656\ : InMux
    port map (
            O => \N__28265\,
            I => \N__28259\
        );

    \I__4655\ : InMux
    port map (
            O => \N__28264\,
            I => \N__28256\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28259\,
            I => \N__28253\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__28256\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__28253\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28248\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\
        );

    \I__4650\ : InMux
    port map (
            O => \N__28245\,
            I => \N__28240\
        );

    \I__4649\ : InMux
    port map (
            O => \N__28244\,
            I => \N__28235\
        );

    \I__4648\ : InMux
    port map (
            O => \N__28243\,
            I => \N__28235\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__28240\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__28235\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\
        );

    \I__4645\ : InMux
    port map (
            O => \N__28230\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\
        );

    \I__4644\ : InMux
    port map (
            O => \N__28227\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28224\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\
        );

    \I__4642\ : InMux
    port map (
            O => \N__28221\,
            I => \N__28217\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28220\,
            I => \N__28213\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__28217\,
            I => \N__28210\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28207\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__28213\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4637\ : Odrv12
    port map (
            O => \N__28210\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__28207\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28200\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\
        );

    \I__4634\ : InMux
    port map (
            O => \N__28197\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\
        );

    \I__4633\ : InMux
    port map (
            O => \N__28194\,
            I => \N__28190\
        );

    \I__4632\ : InMux
    port map (
            O => \N__28193\,
            I => \N__28186\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__28190\,
            I => \N__28183\
        );

    \I__4630\ : InMux
    port map (
            O => \N__28189\,
            I => \N__28180\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__28186\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4628\ : Odrv12
    port map (
            O => \N__28183\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__28180\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\
        );

    \I__4626\ : InMux
    port map (
            O => \N__28173\,
            I => \N__28170\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__28170\,
            I => \N__28167\
        );

    \I__4624\ : Span4Mux_s2_v
    port map (
            O => \N__28167\,
            I => \N__28164\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__28164\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt28\
        );

    \I__4622\ : InMux
    port map (
            O => \N__28161\,
            I => \N__28156\
        );

    \I__4621\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28151\
        );

    \I__4620\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28151\
        );

    \I__4619\ : LocalMux
    port map (
            O => \N__28156\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__28151\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \N__28142\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28145\,
            I => \N__28138\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28133\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28133\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__28138\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__28133\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\
        );

    \I__4611\ : CascadeMux
    port map (
            O => \N__28128\,
            I => \N__28125\
        );

    \I__4610\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__28122\,
            I => \N__28119\
        );

    \I__4608\ : Span4Mux_h
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__4607\ : Odrv4
    port map (
            O => \N__28116\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\
        );

    \I__4606\ : InMux
    port map (
            O => \N__28113\,
            I => \bfn_9_5_0_\
        );

    \I__4605\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28106\
        );

    \I__4604\ : InMux
    port map (
            O => \N__28109\,
            I => \N__28103\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__28106\,
            I => \N__28099\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__28103\,
            I => \N__28096\
        );

    \I__4601\ : InMux
    port map (
            O => \N__28102\,
            I => \N__28093\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__28099\,
            I => \N__28090\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__28096\,
            I => \N__28087\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__28093\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__28090\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4596\ : Odrv4
    port map (
            O => \N__28087\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\
        );

    \I__4595\ : InMux
    port map (
            O => \N__28080\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\
        );

    \I__4594\ : InMux
    port map (
            O => \N__28077\,
            I => \N__28072\
        );

    \I__4593\ : InMux
    port map (
            O => \N__28076\,
            I => \N__28069\
        );

    \I__4592\ : InMux
    port map (
            O => \N__28075\,
            I => \N__28066\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__28072\,
            I => \N__28061\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28061\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__28066\,
            I => \N__28056\
        );

    \I__4588\ : Span4Mux_v
    port map (
            O => \N__28061\,
            I => \N__28056\
        );

    \I__4587\ : Odrv4
    port map (
            O => \N__28056\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\
        );

    \I__4586\ : InMux
    port map (
            O => \N__28053\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\
        );

    \I__4585\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28043\
        );

    \I__4584\ : InMux
    port map (
            O => \N__28049\,
            I => \N__28043\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28048\,
            I => \N__28040\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28037\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__28040\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4580\ : Odrv4
    port map (
            O => \N__28037\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\
        );

    \I__4579\ : InMux
    port map (
            O => \N__28032\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\
        );

    \I__4578\ : CascadeMux
    port map (
            O => \N__28029\,
            I => \N__28025\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__28028\,
            I => \N__28021\
        );

    \I__4576\ : InMux
    port map (
            O => \N__28025\,
            I => \N__28016\
        );

    \I__4575\ : InMux
    port map (
            O => \N__28024\,
            I => \N__28016\
        );

    \I__4574\ : InMux
    port map (
            O => \N__28021\,
            I => \N__28013\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__28016\,
            I => \N__28010\
        );

    \I__4572\ : LocalMux
    port map (
            O => \N__28013\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4571\ : Odrv4
    port map (
            O => \N__28010\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28005\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\
        );

    \I__4569\ : InMux
    port map (
            O => \N__28002\,
            I => \N__27997\
        );

    \I__4568\ : InMux
    port map (
            O => \N__28001\,
            I => \N__27992\
        );

    \I__4567\ : InMux
    port map (
            O => \N__28000\,
            I => \N__27992\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__27997\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__27992\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\
        );

    \I__4564\ : InMux
    port map (
            O => \N__27987\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\
        );

    \I__4563\ : InMux
    port map (
            O => \N__27984\,
            I => \N__27979\
        );

    \I__4562\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27974\
        );

    \I__4561\ : InMux
    port map (
            O => \N__27982\,
            I => \N__27974\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__27979\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__27974\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\
        );

    \I__4558\ : InMux
    port map (
            O => \N__27969\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\
        );

    \I__4557\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27961\
        );

    \I__4556\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27956\
        );

    \I__4555\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27956\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__27961\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4553\ : LocalMux
    port map (
            O => \N__27956\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\
        );

    \I__4552\ : InMux
    port map (
            O => \N__27951\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\
        );

    \I__4551\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27943\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27947\,
            I => \N__27938\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27946\,
            I => \N__27938\
        );

    \I__4548\ : LocalMux
    port map (
            O => \N__27943\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__27938\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\
        );

    \I__4546\ : InMux
    port map (
            O => \N__27933\,
            I => \bfn_9_6_0_\
        );

    \I__4545\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27926\
        );

    \I__4544\ : InMux
    port map (
            O => \N__27929\,
            I => \N__27923\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__27926\,
            I => \N__27920\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__27923\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__27920\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\
        );

    \I__4540\ : InMux
    port map (
            O => \N__27915\,
            I => \bfn_9_4_0_\
        );

    \I__4539\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27908\
        );

    \I__4538\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27905\
        );

    \I__4537\ : LocalMux
    port map (
            O => \N__27908\,
            I => \N__27902\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__27905\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4535\ : Odrv4
    port map (
            O => \N__27902\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\
        );

    \I__4534\ : InMux
    port map (
            O => \N__27897\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\
        );

    \I__4533\ : InMux
    port map (
            O => \N__27894\,
            I => \N__27890\
        );

    \I__4532\ : InMux
    port map (
            O => \N__27893\,
            I => \N__27887\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__27890\,
            I => \N__27884\
        );

    \I__4530\ : LocalMux
    port map (
            O => \N__27887\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4529\ : Odrv4
    port map (
            O => \N__27884\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27879\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\
        );

    \I__4527\ : InMux
    port map (
            O => \N__27876\,
            I => \N__27872\
        );

    \I__4526\ : InMux
    port map (
            O => \N__27875\,
            I => \N__27869\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27872\,
            I => \N__27866\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__27869\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4523\ : Odrv4
    port map (
            O => \N__27866\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\
        );

    \I__4522\ : InMux
    port map (
            O => \N__27861\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\
        );

    \I__4521\ : InMux
    port map (
            O => \N__27858\,
            I => \N__27855\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__27855\,
            I => \N__27851\
        );

    \I__4519\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27848\
        );

    \I__4518\ : Span4Mux_s1_v
    port map (
            O => \N__27851\,
            I => \N__27845\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__27848\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__27845\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\
        );

    \I__4515\ : InMux
    port map (
            O => \N__27840\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\
        );

    \I__4514\ : InMux
    port map (
            O => \N__27837\,
            I => \N__27834\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__27834\,
            I => \N__27830\
        );

    \I__4512\ : InMux
    port map (
            O => \N__27833\,
            I => \N__27827\
        );

    \I__4511\ : Span4Mux_s1_v
    port map (
            O => \N__27830\,
            I => \N__27824\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__27827\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4509\ : Odrv4
    port map (
            O => \N__27824\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\
        );

    \I__4508\ : InMux
    port map (
            O => \N__27819\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27816\,
            I => \N__27812\
        );

    \I__4506\ : InMux
    port map (
            O => \N__27815\,
            I => \N__27809\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__27812\,
            I => \N__27806\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__27809\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__27806\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27801\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\
        );

    \I__4501\ : InMux
    port map (
            O => \N__27798\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\
        );

    \I__4500\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27792\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__27792\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\
        );

    \I__4498\ : CascadeMux
    port map (
            O => \N__27789\,
            I => \N__27785\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__27788\,
            I => \N__27782\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27779\
        );

    \I__4495\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27775\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27779\,
            I => \N__27772\
        );

    \I__4493\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27769\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27775\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__27772\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__27769\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\
        );

    \I__4489\ : InMux
    port map (
            O => \N__27762\,
            I => \N__27758\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27761\,
            I => \N__27755\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__27758\,
            I => \N__27752\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__27755\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4485\ : Odrv4
    port map (
            O => \N__27752\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\
        );

    \I__4484\ : InMux
    port map (
            O => \N__27747\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\
        );

    \I__4483\ : InMux
    port map (
            O => \N__27744\,
            I => \N__27740\
        );

    \I__4482\ : InMux
    port map (
            O => \N__27743\,
            I => \N__27737\
        );

    \I__4481\ : LocalMux
    port map (
            O => \N__27740\,
            I => \N__27734\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__27737\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4479\ : Odrv4
    port map (
            O => \N__27734\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\
        );

    \I__4478\ : InMux
    port map (
            O => \N__27729\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\
        );

    \I__4477\ : InMux
    port map (
            O => \N__27726\,
            I => \N__27722\
        );

    \I__4476\ : InMux
    port map (
            O => \N__27725\,
            I => \N__27719\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__27722\,
            I => \N__27716\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__27719\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__27716\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27711\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\
        );

    \I__4471\ : InMux
    port map (
            O => \N__27708\,
            I => \N__27704\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27707\,
            I => \N__27701\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27698\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__27701\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4467\ : Odrv4
    port map (
            O => \N__27698\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\
        );

    \I__4466\ : InMux
    port map (
            O => \N__27693\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\
        );

    \I__4465\ : InMux
    port map (
            O => \N__27690\,
            I => \N__27686\
        );

    \I__4464\ : InMux
    port map (
            O => \N__27689\,
            I => \N__27683\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27686\,
            I => \N__27680\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27683\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4461\ : Odrv4
    port map (
            O => \N__27680\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\
        );

    \I__4460\ : InMux
    port map (
            O => \N__27675\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\
        );

    \I__4459\ : InMux
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__27669\,
            I => \N__27665\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27668\,
            I => \N__27662\
        );

    \I__4456\ : Span4Mux_s1_v
    port map (
            O => \N__27665\,
            I => \N__27659\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__27662\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4454\ : Odrv4
    port map (
            O => \N__27659\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\
        );

    \I__4453\ : InMux
    port map (
            O => \N__27654\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\
        );

    \I__4452\ : InMux
    port map (
            O => \N__27651\,
            I => \N__27647\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27650\,
            I => \N__27644\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__27647\,
            I => \N__27641\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__27644\,
            I => \N__27636\
        );

    \I__4448\ : Span4Mux_s2_v
    port map (
            O => \N__27641\,
            I => \N__27636\
        );

    \I__4447\ : Odrv4
    port map (
            O => \N__27636\,
            I => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\
        );

    \I__4446\ : InMux
    port map (
            O => \N__27633\,
            I => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\
        );

    \I__4445\ : InMux
    port map (
            O => \N__27630\,
            I => \N__27626\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27629\,
            I => \N__27622\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__27626\,
            I => \N__27619\
        );

    \I__4442\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27616\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__27622\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__27619\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4439\ : LocalMux
    port map (
            O => \N__27616\,
            I => \pwm_generator_inst.counterZ0Z_8\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27605\
        );

    \I__4437\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27601\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__27605\,
            I => \N__27598\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27604\,
            I => \N__27595\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27601\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4433\ : Odrv4
    port map (
            O => \N__27598\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__27595\,
            I => \pwm_generator_inst.counterZ0Z_9\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27583\
        );

    \I__4430\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27580\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27586\,
            I => \N__27577\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27583\,
            I => \N__27574\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__27580\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27577\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__27574\,
            I => \pwm_generator_inst.counterZ0Z_7\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27564\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__27564\,
            I => \N__27559\
        );

    \I__4422\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27556\
        );

    \I__4421\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27553\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__27559\,
            I => \N__27550\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__27556\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__27553\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__27550\,
            I => \pwm_generator_inst.counterZ0Z_0\
        );

    \I__4416\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27539\
        );

    \I__4415\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27535\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__27539\,
            I => \N__27532\
        );

    \I__4413\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27529\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__27535\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4411\ : Odrv4
    port map (
            O => \N__27532\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__27529\,
            I => \pwm_generator_inst.counterZ0Z_2\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27517\
        );

    \I__4408\ : InMux
    port map (
            O => \N__27521\,
            I => \N__27514\
        );

    \I__4407\ : InMux
    port map (
            O => \N__27520\,
            I => \N__27511\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27517\,
            I => \N__27508\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__27514\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__27511\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4403\ : Odrv4
    port map (
            O => \N__27508\,
            I => \pwm_generator_inst.counterZ0Z_4\
        );

    \I__4402\ : InMux
    port map (
            O => \N__27501\,
            I => \N__27496\
        );

    \I__4401\ : InMux
    port map (
            O => \N__27500\,
            I => \N__27493\
        );

    \I__4400\ : InMux
    port map (
            O => \N__27499\,
            I => \N__27490\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__27496\,
            I => \N__27487\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27493\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__27490\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4396\ : Odrv4
    port map (
            O => \N__27487\,
            I => \pwm_generator_inst.counterZ0Z_1\
        );

    \I__4395\ : CascadeMux
    port map (
            O => \N__27480\,
            I => \pwm_generator_inst.un1_counterlto2_0_cascade_\
        );

    \I__4394\ : InMux
    port map (
            O => \N__27477\,
            I => \N__27472\
        );

    \I__4393\ : InMux
    port map (
            O => \N__27476\,
            I => \N__27469\
        );

    \I__4392\ : InMux
    port map (
            O => \N__27475\,
            I => \N__27466\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__27472\,
            I => \N__27463\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__27469\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__27466\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__27463\,
            I => \pwm_generator_inst.counterZ0Z_3\
        );

    \I__4387\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__27453\,
            I => \pwm_generator_inst.un1_counterlto9_2\
        );

    \I__4385\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27445\
        );

    \I__4384\ : InMux
    port map (
            O => \N__27449\,
            I => \N__27442\
        );

    \I__4383\ : InMux
    port map (
            O => \N__27448\,
            I => \N__27439\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27436\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__27442\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__27439\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__27436\,
            I => \pwm_generator_inst.counterZ0Z_6\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__27429\,
            I => \pwm_generator_inst.un1_counterlt9_cascade_\
        );

    \I__4377\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27421\
        );

    \I__4376\ : InMux
    port map (
            O => \N__27425\,
            I => \N__27418\
        );

    \I__4375\ : InMux
    port map (
            O => \N__27424\,
            I => \N__27415\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27421\,
            I => \N__27412\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__27418\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__27415\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4371\ : Odrv4
    port map (
            O => \N__27412\,
            I => \pwm_generator_inst.counterZ0Z_5\
        );

    \I__4370\ : InMux
    port map (
            O => \N__27405\,
            I => \N__27393\
        );

    \I__4369\ : InMux
    port map (
            O => \N__27404\,
            I => \N__27393\
        );

    \I__4368\ : InMux
    port map (
            O => \N__27403\,
            I => \N__27393\
        );

    \I__4367\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27393\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__27393\,
            I => \N__27384\
        );

    \I__4365\ : InMux
    port map (
            O => \N__27392\,
            I => \N__27379\
        );

    \I__4364\ : InMux
    port map (
            O => \N__27391\,
            I => \N__27379\
        );

    \I__4363\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27370\
        );

    \I__4362\ : InMux
    port map (
            O => \N__27389\,
            I => \N__27370\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27370\
        );

    \I__4360\ : InMux
    port map (
            O => \N__27387\,
            I => \N__27370\
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__27384\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__27379\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27370\,
            I => \pwm_generator_inst.un1_counter_0\
        );

    \I__4356\ : InMux
    port map (
            O => \N__27363\,
            I => \N__27360\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__27360\,
            I => \N__27357\
        );

    \I__4354\ : Glb2LocalMux
    port map (
            O => \N__27357\,
            I => \N__27354\
        );

    \I__4353\ : GlobalMux
    port map (
            O => \N__27354\,
            I => clk_12mhz
        );

    \I__4352\ : IoInMux
    port map (
            O => \N__27351\,
            I => \N__27348\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__4350\ : IoSpan4Mux
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__4349\ : Odrv4
    port map (
            O => \N__27342\,
            I => \GB_BUFFER_clk_12mhz_THRU_CO\
        );

    \I__4348\ : InMux
    port map (
            O => \N__27339\,
            I => \N__27336\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__27336\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\
        );

    \I__4346\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__27330\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\
        );

    \I__4344\ : CascadeMux
    port map (
            O => \N__27327\,
            I => \N__27324\
        );

    \I__4343\ : InMux
    port map (
            O => \N__27324\,
            I => \N__27321\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__27321\,
            I => \pwm_generator_inst.threshold_3\
        );

    \I__4341\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27315\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27315\,
            I => \pwm_generator_inst.counter_i_3\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__27312\,
            I => \N__27309\
        );

    \I__4338\ : InMux
    port map (
            O => \N__27309\,
            I => \N__27306\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__27306\,
            I => \N__27303\
        );

    \I__4336\ : Sp12to4
    port map (
            O => \N__27303\,
            I => \N__27300\
        );

    \I__4335\ : Odrv12
    port map (
            O => \N__27300\,
            I => \pwm_generator_inst.threshold_4\
        );

    \I__4334\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27294\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__27294\,
            I => \pwm_generator_inst.counter_i_4\
        );

    \I__4332\ : CascadeMux
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__4331\ : InMux
    port map (
            O => \N__27288\,
            I => \N__27285\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__27282\,
            I => \N__27279\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__27279\,
            I => \pwm_generator_inst.threshold_5\
        );

    \I__4327\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27273\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__27273\,
            I => \pwm_generator_inst.counter_i_5\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__27270\,
            I => \N__27267\
        );

    \I__4324\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27264\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__27264\,
            I => \pwm_generator_inst.threshold_6\
        );

    \I__4322\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__27258\,
            I => \pwm_generator_inst.counter_i_6\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__4319\ : InMux
    port map (
            O => \N__27252\,
            I => \N__27249\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__27249\,
            I => \pwm_generator_inst.threshold_7\
        );

    \I__4317\ : InMux
    port map (
            O => \N__27246\,
            I => \N__27243\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__4315\ : Odrv4
    port map (
            O => \N__27240\,
            I => \pwm_generator_inst.counter_i_7\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__27237\,
            I => \N__27234\
        );

    \I__4313\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27231\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__27231\,
            I => \pwm_generator_inst.threshold_8\
        );

    \I__4311\ : InMux
    port map (
            O => \N__27228\,
            I => \N__27225\
        );

    \I__4310\ : LocalMux
    port map (
            O => \N__27225\,
            I => \pwm_generator_inst.counter_i_8\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__27222\,
            I => \N__27219\
        );

    \I__4308\ : InMux
    port map (
            O => \N__27219\,
            I => \N__27216\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__27216\,
            I => \N__27213\
        );

    \I__4306\ : Odrv12
    port map (
            O => \N__27213\,
            I => \pwm_generator_inst.threshold_9\
        );

    \I__4305\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27207\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__27207\,
            I => \pwm_generator_inst.counter_i_9\
        );

    \I__4303\ : InMux
    port map (
            O => \N__27204\,
            I => \pwm_generator_inst.un14_counter_cry_9\
        );

    \I__4302\ : IoInMux
    port map (
            O => \N__27201\,
            I => \N__27198\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__27198\,
            I => \N__27195\
        );

    \I__4300\ : IoSpan4Mux
    port map (
            O => \N__27195\,
            I => \N__27192\
        );

    \I__4299\ : Span4Mux_s0_v
    port map (
            O => \N__27192\,
            I => \N__27189\
        );

    \I__4298\ : Sp12to4
    port map (
            O => \N__27189\,
            I => \N__27186\
        );

    \I__4297\ : Span12Mux_v
    port map (
            O => \N__27186\,
            I => \N__27183\
        );

    \I__4296\ : Span12Mux_h
    port map (
            O => \N__27183\,
            I => \N__27180\
        );

    \I__4295\ : Odrv12
    port map (
            O => \N__27180\,
            I => pwm_output_c
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__27177\,
            I => \N__27174\
        );

    \I__4293\ : InMux
    port map (
            O => \N__27174\,
            I => \N__27169\
        );

    \I__4292\ : InMux
    port map (
            O => \N__27173\,
            I => \N__27166\
        );

    \I__4291\ : InMux
    port map (
            O => \N__27172\,
            I => \N__27163\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__27169\,
            I => \N__27158\
        );

    \I__4289\ : LocalMux
    port map (
            O => \N__27166\,
            I => \N__27158\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__27163\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__27158\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\
        );

    \I__4286\ : InMux
    port map (
            O => \N__27153\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27150\,
            I => \N__27146\
        );

    \I__4284\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27143\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__27146\,
            I => \N__27140\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__27143\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__27140\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\
        );

    \I__4280\ : CascadeMux
    port map (
            O => \N__27135\,
            I => \N__27132\
        );

    \I__4279\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27127\
        );

    \I__4278\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27124\
        );

    \I__4277\ : InMux
    port map (
            O => \N__27130\,
            I => \N__27121\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__27127\,
            I => \N__27116\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__27124\,
            I => \N__27116\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__27121\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4273\ : Odrv4
    port map (
            O => \N__27116\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\
        );

    \I__4272\ : InMux
    port map (
            O => \N__27111\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\
        );

    \I__4271\ : InMux
    port map (
            O => \N__27108\,
            I => \N__27104\
        );

    \I__4270\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27101\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__27104\,
            I => \N__27098\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__27101\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__4267\ : Odrv4
    port map (
            O => \N__27098\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__27093\,
            I => \N__27090\
        );

    \I__4265\ : InMux
    port map (
            O => \N__27090\,
            I => \N__27085\
        );

    \I__4264\ : InMux
    port map (
            O => \N__27089\,
            I => \N__27082\
        );

    \I__4263\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27079\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__27085\,
            I => \N__27074\
        );

    \I__4261\ : LocalMux
    port map (
            O => \N__27082\,
            I => \N__27074\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__27079\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4259\ : Odrv4
    port map (
            O => \N__27074\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\
        );

    \I__4258\ : InMux
    port map (
            O => \N__27069\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\
        );

    \I__4257\ : InMux
    port map (
            O => \N__27066\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\
        );

    \I__4256\ : CEMux
    port map (
            O => \N__27063\,
            I => \N__27056\
        );

    \I__4255\ : CEMux
    port map (
            O => \N__27062\,
            I => \N__27053\
        );

    \I__4254\ : CEMux
    port map (
            O => \N__27061\,
            I => \N__27050\
        );

    \I__4253\ : CEMux
    port map (
            O => \N__27060\,
            I => \N__27047\
        );

    \I__4252\ : CEMux
    port map (
            O => \N__27059\,
            I => \N__27044\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__27056\,
            I => \N__27041\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__27053\,
            I => \N__27038\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__27050\,
            I => \N__27035\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__27047\,
            I => \N__27032\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__27044\,
            I => \N__27029\
        );

    \I__4246\ : Span4Mux_v
    port map (
            O => \N__27041\,
            I => \N__27026\
        );

    \I__4245\ : Span4Mux_v
    port map (
            O => \N__27038\,
            I => \N__27023\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__27035\,
            I => \N__27020\
        );

    \I__4243\ : Span4Mux_v
    port map (
            O => \N__27032\,
            I => \N__27015\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__27029\,
            I => \N__27015\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__27026\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__27023\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__27020\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__4238\ : Odrv4
    port map (
            O => \N__27015\,
            I => \delay_measurement_inst.delay_tr_timer.N_165_i\
        );

    \I__4237\ : InMux
    port map (
            O => \N__27006\,
            I => \N__26991\
        );

    \I__4236\ : InMux
    port map (
            O => \N__27005\,
            I => \N__26991\
        );

    \I__4235\ : InMux
    port map (
            O => \N__27004\,
            I => \N__26991\
        );

    \I__4234\ : InMux
    port map (
            O => \N__27003\,
            I => \N__26991\
        );

    \I__4233\ : InMux
    port map (
            O => \N__27002\,
            I => \N__26991\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__26991\,
            I => \N__26985\
        );

    \I__4231\ : InMux
    port map (
            O => \N__26990\,
            I => \N__26980\
        );

    \I__4230\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26977\
        );

    \I__4229\ : InMux
    port map (
            O => \N__26988\,
            I => \N__26974\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__26985\,
            I => \N__26971\
        );

    \I__4227\ : InMux
    port map (
            O => \N__26984\,
            I => \N__26966\
        );

    \I__4226\ : InMux
    port map (
            O => \N__26983\,
            I => \N__26966\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__26980\,
            I => \N__26963\
        );

    \I__4224\ : LocalMux
    port map (
            O => \N__26977\,
            I => \N__26960\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__26974\,
            I => \N__26957\
        );

    \I__4222\ : Span4Mux_v
    port map (
            O => \N__26971\,
            I => \N__26952\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__26966\,
            I => \N__26952\
        );

    \I__4220\ : Span12Mux_h
    port map (
            O => \N__26963\,
            I => \N__26949\
        );

    \I__4219\ : Span4Mux_v
    port map (
            O => \N__26960\,
            I => \N__26944\
        );

    \I__4218\ : Span4Mux_h
    port map (
            O => \N__26957\,
            I => \N__26944\
        );

    \I__4217\ : Span4Mux_h
    port map (
            O => \N__26952\,
            I => \N__26941\
        );

    \I__4216\ : Odrv12
    port map (
            O => \N__26949\,
            I => \pwm_generator_inst.N_16\
        );

    \I__4215\ : Odrv4
    port map (
            O => \N__26944\,
            I => \pwm_generator_inst.N_16\
        );

    \I__4214\ : Odrv4
    port map (
            O => \N__26941\,
            I => \pwm_generator_inst.N_16\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26934\,
            I => \N__26931\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26931\,
            I => \N__26928\
        );

    \I__4211\ : Span4Mux_v
    port map (
            O => \N__26928\,
            I => \N__26925\
        );

    \I__4210\ : Span4Mux_h
    port map (
            O => \N__26925\,
            I => \N__26922\
        );

    \I__4209\ : Odrv4
    port map (
            O => \N__26922\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26919\,
            I => \N__26908\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26918\,
            I => \N__26903\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26917\,
            I => \N__26903\
        );

    \I__4205\ : InMux
    port map (
            O => \N__26916\,
            I => \N__26900\
        );

    \I__4204\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26889\
        );

    \I__4203\ : InMux
    port map (
            O => \N__26914\,
            I => \N__26889\
        );

    \I__4202\ : InMux
    port map (
            O => \N__26913\,
            I => \N__26889\
        );

    \I__4201\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26889\
        );

    \I__4200\ : InMux
    port map (
            O => \N__26911\,
            I => \N__26889\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__26908\,
            I => \N__26884\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__26903\,
            I => \N__26884\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26900\,
            I => \N__26879\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__26889\,
            I => \N__26879\
        );

    \I__4195\ : Span4Mux_v
    port map (
            O => \N__26884\,
            I => \N__26875\
        );

    \I__4194\ : Span4Mux_v
    port map (
            O => \N__26879\,
            I => \N__26872\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26878\,
            I => \N__26869\
        );

    \I__4192\ : Sp12to4
    port map (
            O => \N__26875\,
            I => \N__26862\
        );

    \I__4191\ : Sp12to4
    port map (
            O => \N__26872\,
            I => \N__26862\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26869\,
            I => \N__26862\
        );

    \I__4189\ : Odrv12
    port map (
            O => \N__26862\,
            I => \pwm_generator_inst.N_17\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__26859\,
            I => \N__26856\
        );

    \I__4187\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__26853\,
            I => \pwm_generator_inst.threshold_0\
        );

    \I__4185\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__26847\,
            I => \pwm_generator_inst.counter_i_0\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__26844\,
            I => \N__26841\
        );

    \I__4182\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26838\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__4180\ : Odrv4
    port map (
            O => \N__26835\,
            I => \pwm_generator_inst.threshold_1\
        );

    \I__4179\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__26829\,
            I => \pwm_generator_inst.counter_i_1\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__26826\,
            I => \N__26823\
        );

    \I__4176\ : InMux
    port map (
            O => \N__26823\,
            I => \N__26820\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__26820\,
            I => \N__26817\
        );

    \I__4174\ : Odrv12
    port map (
            O => \N__26817\,
            I => \pwm_generator_inst.threshold_2\
        );

    \I__4173\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26811\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26811\,
            I => \pwm_generator_inst.counter_i_2\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__26808\,
            I => \N__26805\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26805\,
            I => \N__26800\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26804\,
            I => \N__26797\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26803\,
            I => \N__26794\
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__26800\,
            I => \N__26789\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__26797\,
            I => \N__26789\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__26794\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__4164\ : Odrv4
    port map (
            O => \N__26789\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26784\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26781\,
            I => \N__26774\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26780\,
            I => \N__26774\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26771\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__26774\,
            I => \N__26768\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__26771\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__4157\ : Odrv4
    port map (
            O => \N__26768\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\
        );

    \I__4156\ : InMux
    port map (
            O => \N__26763\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\
        );

    \I__4155\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26753\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26759\,
            I => \N__26753\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26758\,
            I => \N__26750\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__26753\,
            I => \N__26747\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__26750\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__26747\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\
        );

    \I__4149\ : InMux
    port map (
            O => \N__26742\,
            I => \N__26737\
        );

    \I__4148\ : InMux
    port map (
            O => \N__26741\,
            I => \N__26732\
        );

    \I__4147\ : InMux
    port map (
            O => \N__26740\,
            I => \N__26732\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__26737\,
            I => \N__26728\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26725\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26722\
        );

    \I__4143\ : Sp12to4
    port map (
            O => \N__26728\,
            I => \N__26715\
        );

    \I__4142\ : Span12Mux_s3_v
    port map (
            O => \N__26725\,
            I => \N__26715\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__26722\,
            I => \N__26715\
        );

    \I__4140\ : Odrv12
    port map (
            O => \N__26715\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\
        );

    \I__4139\ : InMux
    port map (
            O => \N__26712\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__26709\,
            I => \N__26705\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26708\,
            I => \N__26702\
        );

    \I__4136\ : InMux
    port map (
            O => \N__26705\,
            I => \N__26699\
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__26702\,
            I => \N__26693\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__26699\,
            I => \N__26693\
        );

    \I__4133\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26690\
        );

    \I__4132\ : Span4Mux_h
    port map (
            O => \N__26693\,
            I => \N__26687\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__26690\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__26687\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\
        );

    \I__4129\ : CascadeMux
    port map (
            O => \N__26682\,
            I => \N__26678\
        );

    \I__4128\ : InMux
    port map (
            O => \N__26681\,
            I => \N__26673\
        );

    \I__4127\ : InMux
    port map (
            O => \N__26678\,
            I => \N__26670\
        );

    \I__4126\ : InMux
    port map (
            O => \N__26677\,
            I => \N__26667\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26676\,
            I => \N__26664\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__26673\,
            I => \N__26661\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26670\,
            I => \N__26654\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__26667\,
            I => \N__26654\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26664\,
            I => \N__26654\
        );

    \I__4120\ : Span4Mux_h
    port map (
            O => \N__26661\,
            I => \N__26649\
        );

    \I__4119\ : Span4Mux_v
    port map (
            O => \N__26654\,
            I => \N__26649\
        );

    \I__4118\ : Odrv4
    port map (
            O => \N__26649\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26646\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__26643\,
            I => \N__26639\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__26642\,
            I => \N__26636\
        );

    \I__4114\ : InMux
    port map (
            O => \N__26639\,
            I => \N__26631\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26636\,
            I => \N__26631\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__26631\,
            I => \N__26627\
        );

    \I__4111\ : InMux
    port map (
            O => \N__26630\,
            I => \N__26624\
        );

    \I__4110\ : Span4Mux_h
    port map (
            O => \N__26627\,
            I => \N__26621\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__26624\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__4108\ : Odrv4
    port map (
            O => \N__26621\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\
        );

    \I__4107\ : InMux
    port map (
            O => \N__26616\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__26613\,
            I => \N__26609\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__26612\,
            I => \N__26606\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26600\
        );

    \I__4103\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26600\
        );

    \I__4102\ : InMux
    port map (
            O => \N__26605\,
            I => \N__26597\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__26600\,
            I => \N__26594\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26597\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__4099\ : Odrv4
    port map (
            O => \N__26594\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\
        );

    \I__4098\ : InMux
    port map (
            O => \N__26589\,
            I => \N__26584\
        );

    \I__4097\ : InMux
    port map (
            O => \N__26588\,
            I => \N__26579\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26579\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__26584\,
            I => \N__26575\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26579\,
            I => \N__26572\
        );

    \I__4093\ : InMux
    port map (
            O => \N__26578\,
            I => \N__26569\
        );

    \I__4092\ : Sp12to4
    port map (
            O => \N__26575\,
            I => \N__26562\
        );

    \I__4091\ : Span12Mux_s6_v
    port map (
            O => \N__26572\,
            I => \N__26562\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__26569\,
            I => \N__26562\
        );

    \I__4089\ : Odrv12
    port map (
            O => \N__26562\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\
        );

    \I__4088\ : InMux
    port map (
            O => \N__26559\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__26556\,
            I => \N__26553\
        );

    \I__4086\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26549\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26546\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26540\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__26546\,
            I => \N__26540\
        );

    \I__4082\ : InMux
    port map (
            O => \N__26545\,
            I => \N__26537\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__26540\,
            I => \N__26534\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__26537\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__26534\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\
        );

    \I__4078\ : InMux
    port map (
            O => \N__26529\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__26526\,
            I => \N__26523\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26523\,
            I => \N__26518\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26522\,
            I => \N__26515\
        );

    \I__4074\ : InMux
    port map (
            O => \N__26521\,
            I => \N__26512\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26518\,
            I => \N__26507\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26515\,
            I => \N__26507\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__26512\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__26507\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\
        );

    \I__4069\ : InMux
    port map (
            O => \N__26502\,
            I => \bfn_8_14_0_\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__26499\,
            I => \N__26496\
        );

    \I__4067\ : InMux
    port map (
            O => \N__26496\,
            I => \N__26493\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__26493\,
            I => \N__26488\
        );

    \I__4065\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26485\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26491\,
            I => \N__26482\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__26488\,
            I => \N__26479\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26485\,
            I => \N__26476\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__26482\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26479\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__26476\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\
        );

    \I__4058\ : InMux
    port map (
            O => \N__26469\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\
        );

    \I__4057\ : CascadeMux
    port map (
            O => \N__26466\,
            I => \N__26463\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26463\,
            I => \N__26458\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26462\,
            I => \N__26455\
        );

    \I__4054\ : InMux
    port map (
            O => \N__26461\,
            I => \N__26452\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26458\,
            I => \N__26447\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__26455\,
            I => \N__26447\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__26452\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__4050\ : Odrv4
    port map (
            O => \N__26447\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\
        );

    \I__4049\ : InMux
    port map (
            O => \N__26442\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\
        );

    \I__4048\ : InMux
    port map (
            O => \N__26439\,
            I => \N__26433\
        );

    \I__4047\ : InMux
    port map (
            O => \N__26438\,
            I => \N__26433\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__26433\,
            I => \N__26429\
        );

    \I__4045\ : InMux
    port map (
            O => \N__26432\,
            I => \N__26426\
        );

    \I__4044\ : Span4Mux_v
    port map (
            O => \N__26429\,
            I => \N__26423\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__26426\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__26423\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26418\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\
        );

    \I__4040\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26408\
        );

    \I__4039\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26408\
        );

    \I__4038\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26405\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__26408\,
            I => \N__26402\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__26405\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__26402\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\
        );

    \I__4034\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26393\
        );

    \I__4033\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26390\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__26393\,
            I => \N__26386\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26383\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26380\
        );

    \I__4029\ : Span4Mux_h
    port map (
            O => \N__26386\,
            I => \N__26376\
        );

    \I__4028\ : Span4Mux_s3_v
    port map (
            O => \N__26383\,
            I => \N__26371\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__26380\,
            I => \N__26371\
        );

    \I__4026\ : InMux
    port map (
            O => \N__26379\,
            I => \N__26368\
        );

    \I__4025\ : Span4Mux_v
    port map (
            O => \N__26376\,
            I => \N__26365\
        );

    \I__4024\ : Span4Mux_v
    port map (
            O => \N__26371\,
            I => \N__26360\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__26368\,
            I => \N__26360\
        );

    \I__4022\ : Odrv4
    port map (
            O => \N__26365\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__4021\ : Odrv4
    port map (
            O => \N__26360\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\
        );

    \I__4020\ : InMux
    port map (
            O => \N__26355\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__26352\,
            I => \N__26348\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__26351\,
            I => \N__26345\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26339\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26345\,
            I => \N__26339\
        );

    \I__4015\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26336\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26333\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__26336\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__26333\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\
        );

    \I__4011\ : InMux
    port map (
            O => \N__26328\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__26325\,
            I => \N__26321\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__26324\,
            I => \N__26318\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26313\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26318\,
            I => \N__26313\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26313\,
            I => \N__26309\
        );

    \I__4005\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26306\
        );

    \I__4004\ : Span4Mux_h
    port map (
            O => \N__26309\,
            I => \N__26303\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__26306\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__26303\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\
        );

    \I__4001\ : InMux
    port map (
            O => \N__26298\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__26295\,
            I => \N__26292\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26287\
        );

    \I__3998\ : InMux
    port map (
            O => \N__26291\,
            I => \N__26284\
        );

    \I__3997\ : InMux
    port map (
            O => \N__26290\,
            I => \N__26281\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__26287\,
            I => \N__26276\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__26284\,
            I => \N__26276\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__26281\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__26276\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26271\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__26268\,
            I => \N__26265\
        );

    \I__3990\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26260\
        );

    \I__3989\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26257\
        );

    \I__3988\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26254\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__26260\,
            I => \N__26249\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__26257\,
            I => \N__26249\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__26254\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__26249\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\
        );

    \I__3983\ : InMux
    port map (
            O => \N__26244\,
            I => \bfn_8_13_0_\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__26241\,
            I => \N__26237\
        );

    \I__3981\ : InMux
    port map (
            O => \N__26240\,
            I => \N__26234\
        );

    \I__3980\ : InMux
    port map (
            O => \N__26237\,
            I => \N__26231\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__26234\,
            I => \N__26225\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__26231\,
            I => \N__26225\
        );

    \I__3977\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26222\
        );

    \I__3976\ : Span4Mux_h
    port map (
            O => \N__26225\,
            I => \N__26219\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__26222\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3974\ : Odrv4
    port map (
            O => \N__26219\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26214\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\
        );

    \I__3972\ : InMux
    port map (
            O => \N__26211\,
            I => \N__26205\
        );

    \I__3971\ : InMux
    port map (
            O => \N__26210\,
            I => \N__26205\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__26205\,
            I => \N__26201\
        );

    \I__3969\ : InMux
    port map (
            O => \N__26204\,
            I => \N__26198\
        );

    \I__3968\ : Span4Mux_v
    port map (
            O => \N__26201\,
            I => \N__26195\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__26198\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3966\ : Odrv4
    port map (
            O => \N__26195\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\
        );

    \I__3965\ : InMux
    port map (
            O => \N__26190\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\
        );

    \I__3964\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26180\
        );

    \I__3963\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26180\
        );

    \I__3962\ : InMux
    port map (
            O => \N__26185\,
            I => \N__26177\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__26180\,
            I => \N__26174\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__26177\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__26174\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26169\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\
        );

    \I__3957\ : CascadeMux
    port map (
            O => \N__26166\,
            I => \N__26162\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__26165\,
            I => \N__26159\
        );

    \I__3955\ : InMux
    port map (
            O => \N__26162\,
            I => \N__26153\
        );

    \I__3954\ : InMux
    port map (
            O => \N__26159\,
            I => \N__26153\
        );

    \I__3953\ : InMux
    port map (
            O => \N__26158\,
            I => \N__26150\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__26153\,
            I => \N__26147\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__26150\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3950\ : Odrv4
    port map (
            O => \N__26147\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\
        );

    \I__3949\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26137\
        );

    \I__3948\ : InMux
    port map (
            O => \N__26141\,
            I => \N__26134\
        );

    \I__3947\ : InMux
    port map (
            O => \N__26140\,
            I => \N__26131\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__26137\,
            I => \N__26126\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__26134\,
            I => \N__26126\
        );

    \I__3944\ : LocalMux
    port map (
            O => \N__26131\,
            I => \N__26122\
        );

    \I__3943\ : Sp12to4
    port map (
            O => \N__26126\,
            I => \N__26119\
        );

    \I__3942\ : InMux
    port map (
            O => \N__26125\,
            I => \N__26116\
        );

    \I__3941\ : Odrv4
    port map (
            O => \N__26122\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__3940\ : Odrv12
    port map (
            O => \N__26119\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__26116\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\
        );

    \I__3938\ : InMux
    port map (
            O => \N__26109\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\
        );

    \I__3937\ : CascadeMux
    port map (
            O => \N__26106\,
            I => \N__26102\
        );

    \I__3936\ : CascadeMux
    port map (
            O => \N__26105\,
            I => \N__26099\
        );

    \I__3935\ : InMux
    port map (
            O => \N__26102\,
            I => \N__26093\
        );

    \I__3934\ : InMux
    port map (
            O => \N__26099\,
            I => \N__26093\
        );

    \I__3933\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26090\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26087\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__26090\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3930\ : Odrv4
    port map (
            O => \N__26087\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\
        );

    \I__3929\ : InMux
    port map (
            O => \N__26082\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__26079\,
            I => \N__26076\
        );

    \I__3927\ : InMux
    port map (
            O => \N__26076\,
            I => \N__26071\
        );

    \I__3926\ : InMux
    port map (
            O => \N__26075\,
            I => \N__26068\
        );

    \I__3925\ : InMux
    port map (
            O => \N__26074\,
            I => \N__26065\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__26071\,
            I => \N__26060\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__26068\,
            I => \N__26060\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__26065\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__26060\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26055\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\
        );

    \I__3919\ : CascadeMux
    port map (
            O => \N__26052\,
            I => \N__26049\
        );

    \I__3918\ : InMux
    port map (
            O => \N__26049\,
            I => \N__26045\
        );

    \I__3917\ : InMux
    port map (
            O => \N__26048\,
            I => \N__26042\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__26045\,
            I => \N__26036\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__26042\,
            I => \N__26036\
        );

    \I__3914\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26033\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__26036\,
            I => \N__26030\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__26033\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__26030\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\
        );

    \I__3910\ : InMux
    port map (
            O => \N__26025\,
            I => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__26022\,
            I => \N__26019\
        );

    \I__3908\ : InMux
    port map (
            O => \N__26019\,
            I => \N__26014\
        );

    \I__3907\ : InMux
    port map (
            O => \N__26018\,
            I => \N__26011\
        );

    \I__3906\ : InMux
    port map (
            O => \N__26017\,
            I => \N__26008\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__26014\,
            I => \N__26003\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26011\,
            I => \N__26003\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__26008\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__26003\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\
        );

    \I__3901\ : InMux
    port map (
            O => \N__25998\,
            I => \N__25995\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__25995\,
            I => \N__25990\
        );

    \I__3899\ : InMux
    port map (
            O => \N__25994\,
            I => \N__25987\
        );

    \I__3898\ : InMux
    port map (
            O => \N__25993\,
            I => \N__25983\
        );

    \I__3897\ : Span4Mux_h
    port map (
            O => \N__25990\,
            I => \N__25980\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__25987\,
            I => \N__25977\
        );

    \I__3895\ : InMux
    port map (
            O => \N__25986\,
            I => \N__25974\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25971\
        );

    \I__3893\ : Span4Mux_v
    port map (
            O => \N__25980\,
            I => \N__25968\
        );

    \I__3892\ : Sp12to4
    port map (
            O => \N__25977\,
            I => \N__25963\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__25974\,
            I => \N__25963\
        );

    \I__3890\ : Odrv4
    port map (
            O => \N__25971\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__3889\ : Odrv4
    port map (
            O => \N__25968\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__3888\ : Odrv12
    port map (
            O => \N__25963\,
            I => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\
        );

    \I__3887\ : InMux
    port map (
            O => \N__25956\,
            I => \bfn_8_12_0_\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__25953\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__25950\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\
        );

    \I__3884\ : InMux
    port map (
            O => \N__25947\,
            I => \N__25944\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__25944\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__25941\,
            I => \N__25938\
        );

    \I__3881\ : InMux
    port map (
            O => \N__25938\,
            I => \N__25935\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__25935\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__25932\,
            I => \N__25928\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25925\
        );

    \I__3877\ : InMux
    port map (
            O => \N__25928\,
            I => \N__25922\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25925\,
            I => \N__25916\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__25922\,
            I => \N__25916\
        );

    \I__3874\ : InMux
    port map (
            O => \N__25921\,
            I => \N__25913\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__25916\,
            I => \N__25910\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25913\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__25910\,
            I => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\
        );

    \I__3870\ : InMux
    port map (
            O => \N__25905\,
            I => \N__25902\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__25902\,
            I => \N__25899\
        );

    \I__3868\ : Span4Mux_s3_v
    port map (
            O => \N__25899\,
            I => \N__25896\
        );

    \I__3867\ : Odrv4
    port map (
            O => \N__25896\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__25893\,
            I => \N__25890\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25890\,
            I => \N__25884\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25884\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__25884\,
            I => \N__25881\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__25881\,
            I => \N__25878\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__25878\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\
        );

    \I__3860\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25870\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25867\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25864\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__25870\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25867\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__25864\,
            I => \elapsed_time_ns_1_RNI1CPBB_0_23\
        );

    \I__3854\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25854\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25851\
        );

    \I__3852\ : Odrv4
    port map (
            O => \N__25851\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\
        );

    \I__3851\ : CascadeMux
    port map (
            O => \N__25848\,
            I => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\
        );

    \I__3850\ : InMux
    port map (
            O => \N__25845\,
            I => \N__25839\
        );

    \I__3849\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25839\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25839\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\
        );

    \I__3847\ : InMux
    port map (
            O => \N__25836\,
            I => \N__25833\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__25833\,
            I => \N__25830\
        );

    \I__3845\ : Odrv12
    port map (
            O => \N__25830\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__25827\,
            I => \N__25824\
        );

    \I__3843\ : InMux
    port map (
            O => \N__25824\,
            I => \N__25821\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25821\,
            I => \N__25818\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__25818\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt26\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25815\,
            I => \N__25812\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__25812\,
            I => \N__25809\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__25809\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__25806\,
            I => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__25803\,
            I => \N__25800\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25800\,
            I => \N__25794\
        );

    \I__3834\ : InMux
    port map (
            O => \N__25799\,
            I => \N__25794\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__25794\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\
        );

    \I__3832\ : InMux
    port map (
            O => \N__25791\,
            I => \N__25785\
        );

    \I__3831\ : InMux
    port map (
            O => \N__25790\,
            I => \N__25785\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__25785\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\
        );

    \I__3829\ : InMux
    port map (
            O => \N__25782\,
            I => \N__25779\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__25779\,
            I => \N__25776\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__25776\,
            I => \N__25772\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25769\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__25772\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__25769\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__25764\,
            I => \N__25760\
        );

    \I__3822\ : CascadeMux
    port map (
            O => \N__25763\,
            I => \N__25757\
        );

    \I__3821\ : InMux
    port map (
            O => \N__25760\,
            I => \N__25754\
        );

    \I__3820\ : InMux
    port map (
            O => \N__25757\,
            I => \N__25751\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__25754\,
            I => \N__25748\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__25751\,
            I => \N__25745\
        );

    \I__3817\ : Span4Mux_v
    port map (
            O => \N__25748\,
            I => \N__25742\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__25745\,
            I => \N__25739\
        );

    \I__3815\ : Odrv4
    port map (
            O => \N__25742\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__25739\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\
        );

    \I__3813\ : InMux
    port map (
            O => \N__25734\,
            I => \N__25731\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__25731\,
            I => \N__25728\
        );

    \I__3811\ : Span4Mux_s3_v
    port map (
            O => \N__25728\,
            I => \N__25725\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__25725\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\
        );

    \I__3809\ : InMux
    port map (
            O => \N__25722\,
            I => \N__25719\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__25719\,
            I => \N__25716\
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__25716\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\
        );

    \I__3806\ : InMux
    port map (
            O => \N__25713\,
            I => \N__25710\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__25710\,
            I => \N__25707\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__25707\,
            I => \N__25703\
        );

    \I__3803\ : InMux
    port map (
            O => \N__25706\,
            I => \N__25700\
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__25703\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__25700\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__25695\,
            I => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25692\,
            I => \N__25686\
        );

    \I__3798\ : InMux
    port map (
            O => \N__25691\,
            I => \N__25686\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__25686\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__25683\,
            I => \N__25679\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__25682\,
            I => \N__25676\
        );

    \I__3794\ : InMux
    port map (
            O => \N__25679\,
            I => \N__25671\
        );

    \I__3793\ : InMux
    port map (
            O => \N__25676\,
            I => \N__25671\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__25671\,
            I => \N__25668\
        );

    \I__3791\ : Span4Mux_h
    port map (
            O => \N__25668\,
            I => \N__25665\
        );

    \I__3790\ : Odrv4
    port map (
            O => \N__25665\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\
        );

    \I__3789\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25659\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__25659\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25656\,
            I => \N__25653\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__25653\,
            I => \N__25650\
        );

    \I__3785\ : Odrv12
    port map (
            O => \N__25650\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__3783\ : InMux
    port map (
            O => \N__25644\,
            I => \N__25641\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__25638\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt24\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25632\,
            I => \N__25629\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__25629\,
            I => \N__25625\
        );

    \I__3777\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25622\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__25625\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__25622\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25\
        );

    \I__3774\ : CascadeMux
    port map (
            O => \N__25617\,
            I => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__25614\,
            I => \N__25610\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__25613\,
            I => \N__25607\
        );

    \I__3771\ : InMux
    port map (
            O => \N__25610\,
            I => \N__25602\
        );

    \I__3770\ : InMux
    port map (
            O => \N__25607\,
            I => \N__25602\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__25602\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\
        );

    \I__3768\ : InMux
    port map (
            O => \N__25599\,
            I => \N__25596\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__25596\,
            I => \N__25593\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__25593\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\
        );

    \I__3765\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__25587\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__25584\,
            I => \N__25581\
        );

    \I__3762\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25578\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__25578\,
            I => \N__25575\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__25575\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt18\
        );

    \I__3759\ : InMux
    port map (
            O => \N__25572\,
            I => \N__25569\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25566\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__25566\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__25563\,
            I => \N__25560\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25557\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__25557\,
            I => \N__25554\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__25554\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt20\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__25551\,
            I => \N__25548\
        );

    \I__3751\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25545\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__25545\,
            I => \N__25542\
        );

    \I__3749\ : Span12Mux_s5_v
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__3748\ : Odrv12
    port map (
            O => \N__25539\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt30\
        );

    \I__3747\ : InMux
    port map (
            O => \N__25536\,
            I => \phase_controller_inst1.stoper_tr.un4_running_cry_30\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__25533\,
            I => \N__25530\
        );

    \I__3745\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25527\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__25527\,
            I => \phase_controller_inst1.stoper_tr.un4_running_lt22\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__25524\,
            I => \N__25521\
        );

    \I__3742\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25518\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__25518\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__25515\,
            I => \N__25512\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25512\,
            I => \N__25509\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__25509\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\
        );

    \I__3737\ : InMux
    port map (
            O => \N__25506\,
            I => \N__25503\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25503\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__25500\,
            I => \N__25497\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25494\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__25494\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__25491\,
            I => \N__25488\
        );

    \I__3731\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25485\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__25485\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__25482\,
            I => \N__25479\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25476\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25476\,
            I => \N__25473\
        );

    \I__3726\ : Odrv4
    port map (
            O => \N__25473\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__25470\,
            I => \N__25467\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25464\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__25464\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__25461\,
            I => \N__25458\
        );

    \I__3721\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25455\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__25455\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25452\,
            I => \N__25449\
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__25449\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\
        );

    \I__3717\ : InMux
    port map (
            O => \N__25446\,
            I => \pwm_generator_inst.counter_cry_8\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__25443\,
            I => \N__25440\
        );

    \I__3715\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25437\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__25437\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\
        );

    \I__3713\ : InMux
    port map (
            O => \N__25434\,
            I => \N__25431\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__25431\,
            I => \N__25428\
        );

    \I__3711\ : Span4Mux_s1_v
    port map (
            O => \N__25428\,
            I => \N__25425\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__25425\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25416\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__3705\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__25407\,
            I => \N__25404\
        );

    \I__3703\ : Odrv4
    port map (
            O => \N__25404\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\
        );

    \I__3702\ : CascadeMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__3701\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25395\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__25395\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25389\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__25389\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__25386\,
            I => \N__25383\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25383\,
            I => \N__25380\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__25380\,
            I => \N__25377\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__25377\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__25374\,
            I => \N__25371\
        );

    \I__3692\ : InMux
    port map (
            O => \N__25371\,
            I => \N__25368\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__25368\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\
        );

    \I__3690\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25362\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__25362\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__25359\,
            I => \N__25356\
        );

    \I__3687\ : InMux
    port map (
            O => \N__25356\,
            I => \N__25353\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__25353\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__25350\,
            I => \N__25347\
        );

    \I__3684\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25344\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__25344\,
            I => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25341\,
            I => \bfn_7_26_0_\
        );

    \I__3681\ : InMux
    port map (
            O => \N__25338\,
            I => \pwm_generator_inst.counter_cry_0\
        );

    \I__3680\ : InMux
    port map (
            O => \N__25335\,
            I => \pwm_generator_inst.counter_cry_1\
        );

    \I__3679\ : InMux
    port map (
            O => \N__25332\,
            I => \pwm_generator_inst.counter_cry_2\
        );

    \I__3678\ : InMux
    port map (
            O => \N__25329\,
            I => \pwm_generator_inst.counter_cry_3\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25326\,
            I => \pwm_generator_inst.counter_cry_4\
        );

    \I__3676\ : InMux
    port map (
            O => \N__25323\,
            I => \pwm_generator_inst.counter_cry_5\
        );

    \I__3675\ : InMux
    port map (
            O => \N__25320\,
            I => \pwm_generator_inst.counter_cry_6\
        );

    \I__3674\ : InMux
    port map (
            O => \N__25317\,
            I => \bfn_7_27_0_\
        );

    \I__3673\ : InMux
    port map (
            O => \N__25314\,
            I => \N__25308\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25313\,
            I => \N__25301\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25312\,
            I => \N__25301\
        );

    \I__3670\ : InMux
    port map (
            O => \N__25311\,
            I => \N__25301\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25308\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__25301\,
            I => \delay_measurement_inst.delay_tr_timer.runningZ0\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__25296\,
            I => \N__25293\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25286\
        );

    \I__3665\ : InMux
    port map (
            O => \N__25292\,
            I => \N__25286\
        );

    \I__3664\ : InMux
    port map (
            O => \N__25291\,
            I => \N__25283\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__25286\,
            I => \N__25280\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__25283\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__25280\,
            I => \delay_measurement_inst.stop_timer_trZ0\
        );

    \I__3660\ : InMux
    port map (
            O => \N__25275\,
            I => \N__25269\
        );

    \I__3659\ : InMux
    port map (
            O => \N__25274\,
            I => \N__25266\
        );

    \I__3658\ : InMux
    port map (
            O => \N__25273\,
            I => \N__25263\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25260\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__25269\,
            I => \N__25255\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__25266\,
            I => \N__25255\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__25263\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__25260\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3652\ : Odrv4
    port map (
            O => \N__25255\,
            I => \delay_measurement_inst.start_timer_trZ0\
        );

    \I__3651\ : ClkMux
    port map (
            O => \N__25248\,
            I => \N__25242\
        );

    \I__3650\ : ClkMux
    port map (
            O => \N__25247\,
            I => \N__25242\
        );

    \I__3649\ : GlobalMux
    port map (
            O => \N__25242\,
            I => \N__25239\
        );

    \I__3648\ : gio2CtrlBuf
    port map (
            O => \N__25239\,
            I => delay_tr_input_c_g
        );

    \I__3647\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25233\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__25233\,
            I => \N__25230\
        );

    \I__3645\ : Odrv12
    port map (
            O => \N__25230\,
            I => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25227\,
            I => \N__25224\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__25224\,
            I => \N__25221\
        );

    \I__3642\ : Odrv12
    port map (
            O => \N__25221\,
            I => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\
        );

    \I__3641\ : InMux
    port map (
            O => \N__25218\,
            I => \N__25215\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__25215\,
            I => \N__25212\
        );

    \I__3639\ : Odrv12
    port map (
            O => \N__25212\,
            I => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__25209\,
            I => \N__25206\
        );

    \I__3637\ : InMux
    port map (
            O => \N__25206\,
            I => \N__25203\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25203\,
            I => \N__25200\
        );

    \I__3635\ : Odrv12
    port map (
            O => \N__25200\,
            I => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25197\,
            I => \N__25194\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__25194\,
            I => \N__25191\
        );

    \I__3632\ : Odrv12
    port map (
            O => \N__25191\,
            I => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\
        );

    \I__3631\ : InMux
    port map (
            O => \N__25188\,
            I => \N__25185\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__25185\,
            I => \N__25182\
        );

    \I__3629\ : Odrv12
    port map (
            O => \N__25182\,
            I => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\
        );

    \I__3628\ : InMux
    port map (
            O => \N__25179\,
            I => \bfn_7_16_0_\
        );

    \I__3627\ : InMux
    port map (
            O => \N__25176\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_24\
        );

    \I__3626\ : InMux
    port map (
            O => \N__25173\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_25\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25170\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_26\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25167\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_27\
        );

    \I__3623\ : InMux
    port map (
            O => \N__25164\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_28\
        );

    \I__3622\ : CEMux
    port map (
            O => \N__25161\,
            I => \N__25156\
        );

    \I__3621\ : CEMux
    port map (
            O => \N__25160\,
            I => \N__25153\
        );

    \I__3620\ : CEMux
    port map (
            O => \N__25159\,
            I => \N__25150\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__25156\,
            I => \N__25146\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__25153\,
            I => \N__25141\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__25150\,
            I => \N__25141\
        );

    \I__3616\ : CEMux
    port map (
            O => \N__25149\,
            I => \N__25138\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__25146\,
            I => \N__25135\
        );

    \I__3614\ : Span4Mux_v
    port map (
            O => \N__25141\,
            I => \N__25132\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__25138\,
            I => \N__25129\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__25135\,
            I => \delay_measurement_inst.delay_tr_timer.N_166_i\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__25132\,
            I => \delay_measurement_inst.delay_tr_timer.N_166_i\
        );

    \I__3610\ : Odrv12
    port map (
            O => \N__25129\,
            I => \delay_measurement_inst.delay_tr_timer.N_166_i\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25084\
        );

    \I__3608\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25084\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25120\,
            I => \N__25084\
        );

    \I__3606\ : InMux
    port map (
            O => \N__25119\,
            I => \N__25084\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25075\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25117\,
            I => \N__25075\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25116\,
            I => \N__25075\
        );

    \I__3602\ : InMux
    port map (
            O => \N__25115\,
            I => \N__25075\
        );

    \I__3601\ : InMux
    port map (
            O => \N__25114\,
            I => \N__25066\
        );

    \I__3600\ : InMux
    port map (
            O => \N__25113\,
            I => \N__25066\
        );

    \I__3599\ : InMux
    port map (
            O => \N__25112\,
            I => \N__25066\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25111\,
            I => \N__25066\
        );

    \I__3597\ : InMux
    port map (
            O => \N__25110\,
            I => \N__25057\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25109\,
            I => \N__25057\
        );

    \I__3595\ : InMux
    port map (
            O => \N__25108\,
            I => \N__25057\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25107\,
            I => \N__25057\
        );

    \I__3593\ : InMux
    port map (
            O => \N__25106\,
            I => \N__25048\
        );

    \I__3592\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25048\
        );

    \I__3591\ : InMux
    port map (
            O => \N__25104\,
            I => \N__25048\
        );

    \I__3590\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25048\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25039\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25039\
        );

    \I__3587\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25039\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25039\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25098\,
            I => \N__25034\
        );

    \I__3584\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25034\
        );

    \I__3583\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25025\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25095\,
            I => \N__25025\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25025\
        );

    \I__3580\ : InMux
    port map (
            O => \N__25093\,
            I => \N__25025\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__25084\,
            I => \N__25012\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__25075\,
            I => \N__25012\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__25066\,
            I => \N__25012\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__25057\,
            I => \N__25012\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__25048\,
            I => \N__25012\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__25039\,
            I => \N__25012\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__25034\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25025\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3571\ : Odrv12
    port map (
            O => \N__25012\,
            I => \delay_measurement_inst.delay_tr_timer.running_i\
        );

    \I__3570\ : InMux
    port map (
            O => \N__25005\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_14\
        );

    \I__3569\ : InMux
    port map (
            O => \N__25002\,
            I => \bfn_7_15_0_\
        );

    \I__3568\ : InMux
    port map (
            O => \N__24999\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_16\
        );

    \I__3567\ : InMux
    port map (
            O => \N__24996\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_17\
        );

    \I__3566\ : InMux
    port map (
            O => \N__24993\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_18\
        );

    \I__3565\ : InMux
    port map (
            O => \N__24990\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_19\
        );

    \I__3564\ : InMux
    port map (
            O => \N__24987\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_20\
        );

    \I__3563\ : InMux
    port map (
            O => \N__24984\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_21\
        );

    \I__3562\ : InMux
    port map (
            O => \N__24981\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_22\
        );

    \I__3561\ : InMux
    port map (
            O => \N__24978\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_5\
        );

    \I__3560\ : InMux
    port map (
            O => \N__24975\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_6\
        );

    \I__3559\ : InMux
    port map (
            O => \N__24972\,
            I => \bfn_7_14_0_\
        );

    \I__3558\ : InMux
    port map (
            O => \N__24969\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_8\
        );

    \I__3557\ : InMux
    port map (
            O => \N__24966\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_9\
        );

    \I__3556\ : InMux
    port map (
            O => \N__24963\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_10\
        );

    \I__3555\ : InMux
    port map (
            O => \N__24960\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_11\
        );

    \I__3554\ : InMux
    port map (
            O => \N__24957\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_12\
        );

    \I__3553\ : InMux
    port map (
            O => \N__24954\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_13\
        );

    \I__3552\ : InMux
    port map (
            O => \N__24951\,
            I => \bfn_7_13_0_\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24948\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_0\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24945\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_1\
        );

    \I__3549\ : InMux
    port map (
            O => \N__24942\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_2\
        );

    \I__3548\ : InMux
    port map (
            O => \N__24939\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_3\
        );

    \I__3547\ : InMux
    port map (
            O => \N__24936\,
            I => \delay_measurement_inst.delay_tr_timer.counter_cry_4\
        );

    \I__3546\ : InMux
    port map (
            O => \N__24933\,
            I => \N__24927\
        );

    \I__3545\ : InMux
    port map (
            O => \N__24932\,
            I => \N__24927\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__24927\,
            I => \N__24924\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__24924\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\
        );

    \I__3542\ : InMux
    port map (
            O => \N__24921\,
            I => \N__24918\
        );

    \I__3541\ : LocalMux
    port map (
            O => \N__24918\,
            I => \N__24914\
        );

    \I__3540\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24910\
        );

    \I__3539\ : Span4Mux_v
    port map (
            O => \N__24914\,
            I => \N__24907\
        );

    \I__3538\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24904\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24910\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__3536\ : Odrv4
    port map (
            O => \N__24907\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__24904\,
            I => \elapsed_time_ns_1_RNIJI91B_0_7\
        );

    \I__3534\ : InMux
    port map (
            O => \N__24897\,
            I => \N__24892\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24896\,
            I => \N__24889\
        );

    \I__3532\ : InMux
    port map (
            O => \N__24895\,
            I => \N__24886\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__24892\,
            I => \N__24883\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__24889\,
            I => \N__24880\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__24886\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__3528\ : Odrv12
    port map (
            O => \N__24883\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__24880\,
            I => \elapsed_time_ns_1_RNIU7OBB_0_11\
        );

    \I__3526\ : InMux
    port map (
            O => \N__24873\,
            I => \N__24867\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24872\,
            I => \N__24867\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__24867\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__24864\,
            I => \N__24860\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24863\,
            I => \N__24855\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24855\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24855\,
            I => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\
        );

    \I__3519\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24844\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24848\,
            I => \N__24841\
        );

    \I__3516\ : InMux
    port map (
            O => \N__24847\,
            I => \N__24838\
        );

    \I__3515\ : Span4Mux_h
    port map (
            O => \N__24844\,
            I => \N__24835\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__24841\,
            I => \N__24832\
        );

    \I__3513\ : LocalMux
    port map (
            O => \N__24838\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__24835\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__24832\,
            I => \elapsed_time_ns_1_RNI2COBB_0_15\
        );

    \I__3510\ : InMux
    port map (
            O => \N__24825\,
            I => \N__24821\
        );

    \I__3509\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24818\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__24821\,
            I => \N__24813\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__24818\,
            I => \N__24813\
        );

    \I__3506\ : Odrv4
    port map (
            O => \N__24813\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__24810\,
            I => \N__24806\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__24809\,
            I => \N__24803\
        );

    \I__3503\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24800\
        );

    \I__3502\ : InMux
    port map (
            O => \N__24803\,
            I => \N__24797\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__24800\,
            I => \N__24792\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__24797\,
            I => \N__24792\
        );

    \I__3499\ : Odrv12
    port map (
            O => \N__24792\,
            I => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\
        );

    \I__3498\ : InMux
    port map (
            O => \N__24789\,
            I => \N__24786\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24786\,
            I => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24783\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_14\
        );

    \I__3495\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24777\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__24777\,
            I => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\
        );

    \I__3493\ : InMux
    port map (
            O => \N__24774\,
            I => \bfn_5_25_0_\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__24771\,
            I => \N__24767\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24770\,
            I => \N__24761\
        );

    \I__3490\ : InMux
    port map (
            O => \N__24767\,
            I => \N__24758\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__24766\,
            I => \N__24752\
        );

    \I__3488\ : CascadeMux
    port map (
            O => \N__24765\,
            I => \N__24749\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__24764\,
            I => \N__24746\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__24761\,
            I => \N__24742\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24758\,
            I => \N__24739\
        );

    \I__3484\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24733\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24730\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24755\,
            I => \N__24721\
        );

    \I__3481\ : InMux
    port map (
            O => \N__24752\,
            I => \N__24721\
        );

    \I__3480\ : InMux
    port map (
            O => \N__24749\,
            I => \N__24721\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24746\,
            I => \N__24721\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24718\
        );

    \I__3477\ : Span4Mux_v
    port map (
            O => \N__24742\,
            I => \N__24713\
        );

    \I__3476\ : Span4Mux_v
    port map (
            O => \N__24739\,
            I => \N__24713\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24738\,
            I => \N__24706\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24737\,
            I => \N__24706\
        );

    \I__3473\ : InMux
    port map (
            O => \N__24736\,
            I => \N__24706\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24733\,
            I => \N__24697\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__24730\,
            I => \N__24697\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__24721\,
            I => \N__24697\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24718\,
            I => \N__24697\
        );

    \I__3468\ : Odrv4
    port map (
            O => \N__24713\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__24706\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3466\ : Odrv12
    port map (
            O => \N__24697\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24687\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24684\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__24684\,
            I => \N__24681\
        );

    \I__3462\ : Span4Mux_h
    port map (
            O => \N__24681\,
            I => \N__24678\
        );

    \I__3461\ : Odrv4
    port map (
            O => \N__24678\,
            I => \pwm_generator_inst.un2_threshold_1_22\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__24675\,
            I => \N__24672\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24672\,
            I => \N__24669\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__24669\,
            I => \N__24666\
        );

    \I__3457\ : Span12Mux_h
    port map (
            O => \N__24666\,
            I => \N__24663\
        );

    \I__3456\ : Odrv12
    port map (
            O => \N__24663\,
            I => \pwm_generator_inst.un2_threshold_2_7\
        );

    \I__3455\ : InMux
    port map (
            O => \N__24660\,
            I => \N__24657\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__24657\,
            I => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\
        );

    \I__3453\ : InMux
    port map (
            O => \N__24654\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_6\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24651\,
            I => \N__24648\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24645\
        );

    \I__3450\ : Span4Mux_h
    port map (
            O => \N__24645\,
            I => \N__24642\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__24642\,
            I => \N__24639\
        );

    \I__3448\ : Odrv4
    port map (
            O => \N__24639\,
            I => \pwm_generator_inst.un2_threshold_1_23\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__3446\ : InMux
    port map (
            O => \N__24633\,
            I => \N__24630\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__24630\,
            I => \N__24627\
        );

    \I__3444\ : Span4Mux_h
    port map (
            O => \N__24627\,
            I => \N__24624\
        );

    \I__3443\ : Sp12to4
    port map (
            O => \N__24624\,
            I => \N__24621\
        );

    \I__3442\ : Span12Mux_h
    port map (
            O => \N__24621\,
            I => \N__24618\
        );

    \I__3441\ : Odrv12
    port map (
            O => \N__24618\,
            I => \pwm_generator_inst.un2_threshold_2_8\
        );

    \I__3440\ : InMux
    port map (
            O => \N__24615\,
            I => \N__24612\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__24612\,
            I => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\
        );

    \I__3438\ : InMux
    port map (
            O => \N__24609\,
            I => \bfn_5_24_0_\
        );

    \I__3437\ : InMux
    port map (
            O => \N__24606\,
            I => \N__24603\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__24603\,
            I => \N__24600\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__24600\,
            I => \N__24597\
        );

    \I__3434\ : Span4Mux_h
    port map (
            O => \N__24597\,
            I => \N__24594\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__24594\,
            I => \pwm_generator_inst.un2_threshold_1_24\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__24591\,
            I => \N__24588\
        );

    \I__3431\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24582\
        );

    \I__3429\ : Span4Mux_h
    port map (
            O => \N__24582\,
            I => \N__24579\
        );

    \I__3428\ : Sp12to4
    port map (
            O => \N__24579\,
            I => \N__24576\
        );

    \I__3427\ : Span12Mux_h
    port map (
            O => \N__24576\,
            I => \N__24573\
        );

    \I__3426\ : Odrv12
    port map (
            O => \N__24573\,
            I => \pwm_generator_inst.un2_threshold_2_9\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24570\,
            I => \N__24567\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24567\,
            I => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\
        );

    \I__3423\ : InMux
    port map (
            O => \N__24564\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_8\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__24561\,
            I => \N__24558\
        );

    \I__3421\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24555\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__24555\,
            I => \N__24552\
        );

    \I__3419\ : Span4Mux_h
    port map (
            O => \N__24552\,
            I => \N__24549\
        );

    \I__3418\ : Sp12to4
    port map (
            O => \N__24549\,
            I => \N__24546\
        );

    \I__3417\ : Span12Mux_h
    port map (
            O => \N__24546\,
            I => \N__24543\
        );

    \I__3416\ : Odrv12
    port map (
            O => \N__24543\,
            I => \pwm_generator_inst.un2_threshold_2_10\
        );

    \I__3415\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24537\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__24537\,
            I => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24534\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_9\
        );

    \I__3412\ : InMux
    port map (
            O => \N__24531\,
            I => \N__24528\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__24528\,
            I => \N__24525\
        );

    \I__3410\ : Span12Mux_s6_h
    port map (
            O => \N__24525\,
            I => \N__24522\
        );

    \I__3409\ : Span12Mux_h
    port map (
            O => \N__24522\,
            I => \N__24519\
        );

    \I__3408\ : Odrv12
    port map (
            O => \N__24519\,
            I => \pwm_generator_inst.un2_threshold_2_11\
        );

    \I__3407\ : InMux
    port map (
            O => \N__24516\,
            I => \N__24513\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__24513\,
            I => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\
        );

    \I__3405\ : InMux
    port map (
            O => \N__24510\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_10\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__24507\,
            I => \N__24504\
        );

    \I__3403\ : InMux
    port map (
            O => \N__24504\,
            I => \N__24501\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__24501\,
            I => \N__24498\
        );

    \I__3401\ : Span12Mux_h
    port map (
            O => \N__24498\,
            I => \N__24495\
        );

    \I__3400\ : Odrv12
    port map (
            O => \N__24495\,
            I => \pwm_generator_inst.un2_threshold_2_12\
        );

    \I__3399\ : InMux
    port map (
            O => \N__24492\,
            I => \N__24489\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__24489\,
            I => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\
        );

    \I__3397\ : InMux
    port map (
            O => \N__24486\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_11\
        );

    \I__3396\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24480\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__24480\,
            I => \N__24477\
        );

    \I__3394\ : Span12Mux_h
    port map (
            O => \N__24477\,
            I => \N__24474\
        );

    \I__3393\ : Odrv12
    port map (
            O => \N__24474\,
            I => \pwm_generator_inst.un2_threshold_2_13\
        );

    \I__3392\ : InMux
    port map (
            O => \N__24471\,
            I => \N__24468\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__24468\,
            I => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\
        );

    \I__3390\ : InMux
    port map (
            O => \N__24465\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_12\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__24462\,
            I => \N__24459\
        );

    \I__3388\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24453\
        );

    \I__3386\ : Sp12to4
    port map (
            O => \N__24453\,
            I => \N__24450\
        );

    \I__3385\ : Span12Mux_s11_h
    port map (
            O => \N__24450\,
            I => \N__24447\
        );

    \I__3384\ : Span12Mux_h
    port map (
            O => \N__24447\,
            I => \N__24444\
        );

    \I__3383\ : Odrv12
    port map (
            O => \N__24444\,
            I => \pwm_generator_inst.un2_threshold_2_14\
        );

    \I__3382\ : InMux
    port map (
            O => \N__24441\,
            I => \N__24438\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__24438\,
            I => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24435\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_13\
        );

    \I__3379\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24429\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24429\,
            I => \N__24426\
        );

    \I__3377\ : Span12Mux_s9_h
    port map (
            O => \N__24426\,
            I => \N__24423\
        );

    \I__3376\ : Span12Mux_h
    port map (
            O => \N__24423\,
            I => \N__24420\
        );

    \I__3375\ : Odrv12
    port map (
            O => \N__24420\,
            I => \pwm_generator_inst.un2_threshold_2_0\
        );

    \I__3374\ : CascadeMux
    port map (
            O => \N__24417\,
            I => \N__24414\
        );

    \I__3373\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24411\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__24411\,
            I => \N__24408\
        );

    \I__3371\ : Span4Mux_h
    port map (
            O => \N__24408\,
            I => \N__24405\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__24402\,
            I => \pwm_generator_inst.un2_threshold_1_15\
        );

    \I__3368\ : InMux
    port map (
            O => \N__24399\,
            I => \N__24396\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__24396\,
            I => \pwm_generator_inst.un3_threshold_axbZ0Z_4\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24390\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__24390\,
            I => \N__24387\
        );

    \I__3364\ : Span4Mux_h
    port map (
            O => \N__24387\,
            I => \N__24384\
        );

    \I__3363\ : Sp12to4
    port map (
            O => \N__24384\,
            I => \N__24381\
        );

    \I__3362\ : Span12Mux_h
    port map (
            O => \N__24381\,
            I => \N__24378\
        );

    \I__3361\ : Odrv12
    port map (
            O => \N__24378\,
            I => \pwm_generator_inst.un2_threshold_2_1\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__24375\,
            I => \N__24372\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24369\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24366\
        );

    \I__3357\ : Span4Mux_h
    port map (
            O => \N__24366\,
            I => \N__24363\
        );

    \I__3356\ : Span4Mux_h
    port map (
            O => \N__24363\,
            I => \N__24360\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__24360\,
            I => \pwm_generator_inst.un2_threshold_1_16\
        );

    \I__3354\ : InMux
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24354\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\
        );

    \I__3352\ : InMux
    port map (
            O => \N__24351\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_0\
        );

    \I__3351\ : InMux
    port map (
            O => \N__24348\,
            I => \N__24345\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__3349\ : Span12Mux_s7_h
    port map (
            O => \N__24342\,
            I => \N__24339\
        );

    \I__3348\ : Span12Mux_h
    port map (
            O => \N__24339\,
            I => \N__24336\
        );

    \I__3347\ : Odrv12
    port map (
            O => \N__24336\,
            I => \pwm_generator_inst.un2_threshold_2_2\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__24333\,
            I => \N__24330\
        );

    \I__3345\ : InMux
    port map (
            O => \N__24330\,
            I => \N__24327\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__24327\,
            I => \N__24324\
        );

    \I__3343\ : Span4Mux_h
    port map (
            O => \N__24324\,
            I => \N__24321\
        );

    \I__3342\ : Span4Mux_h
    port map (
            O => \N__24321\,
            I => \N__24318\
        );

    \I__3341\ : Odrv4
    port map (
            O => \N__24318\,
            I => \pwm_generator_inst.un2_threshold_1_17\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__24315\,
            I => \N__24312\
        );

    \I__3339\ : InMux
    port map (
            O => \N__24312\,
            I => \N__24309\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__24309\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\
        );

    \I__3337\ : InMux
    port map (
            O => \N__24306\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_1\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24300\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24297\
        );

    \I__3334\ : Span12Mux_s6_h
    port map (
            O => \N__24297\,
            I => \N__24294\
        );

    \I__3333\ : Span12Mux_h
    port map (
            O => \N__24294\,
            I => \N__24291\
        );

    \I__3332\ : Odrv12
    port map (
            O => \N__24291\,
            I => \pwm_generator_inst.un2_threshold_2_3\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__24288\,
            I => \N__24285\
        );

    \I__3330\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24282\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__24282\,
            I => \N__24279\
        );

    \I__3328\ : Span12Mux_h
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__3327\ : Odrv12
    port map (
            O => \N__24276\,
            I => \pwm_generator_inst.un2_threshold_1_18\
        );

    \I__3326\ : InMux
    port map (
            O => \N__24273\,
            I => \N__24270\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__24270\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\
        );

    \I__3324\ : InMux
    port map (
            O => \N__24267\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_2\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24261\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__24261\,
            I => \N__24258\
        );

    \I__3321\ : Span12Mux_v
    port map (
            O => \N__24258\,
            I => \N__24255\
        );

    \I__3320\ : Odrv12
    port map (
            O => \N__24255\,
            I => \pwm_generator_inst.un2_threshold_1_19\
        );

    \I__3319\ : CascadeMux
    port map (
            O => \N__24252\,
            I => \N__24249\
        );

    \I__3318\ : InMux
    port map (
            O => \N__24249\,
            I => \N__24246\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__24246\,
            I => \N__24243\
        );

    \I__3316\ : Span12Mux_h
    port map (
            O => \N__24243\,
            I => \N__24240\
        );

    \I__3315\ : Odrv12
    port map (
            O => \N__24240\,
            I => \pwm_generator_inst.un2_threshold_2_4\
        );

    \I__3314\ : InMux
    port map (
            O => \N__24237\,
            I => \N__24234\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__24234\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\
        );

    \I__3312\ : InMux
    port map (
            O => \N__24231\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_3\
        );

    \I__3311\ : InMux
    port map (
            O => \N__24228\,
            I => \N__24225\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__24225\,
            I => \N__24222\
        );

    \I__3309\ : Span12Mux_h
    port map (
            O => \N__24222\,
            I => \N__24219\
        );

    \I__3308\ : Odrv12
    port map (
            O => \N__24219\,
            I => \pwm_generator_inst.un2_threshold_2_5\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__24216\,
            I => \N__24213\
        );

    \I__3306\ : InMux
    port map (
            O => \N__24213\,
            I => \N__24210\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__24210\,
            I => \N__24207\
        );

    \I__3304\ : Span4Mux_h
    port map (
            O => \N__24207\,
            I => \N__24204\
        );

    \I__3303\ : Span4Mux_h
    port map (
            O => \N__24204\,
            I => \N__24201\
        );

    \I__3302\ : Odrv4
    port map (
            O => \N__24201\,
            I => \pwm_generator_inst.un2_threshold_1_20\
        );

    \I__3301\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24195\
        );

    \I__3300\ : LocalMux
    port map (
            O => \N__24195\,
            I => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\
        );

    \I__3299\ : InMux
    port map (
            O => \N__24192\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_4\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24186\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24186\,
            I => \N__24183\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__24183\,
            I => \N__24180\
        );

    \I__3295\ : Span4Mux_h
    port map (
            O => \N__24180\,
            I => \N__24177\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__24177\,
            I => \pwm_generator_inst.un2_threshold_1_21\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__24174\,
            I => \N__24171\
        );

    \I__3292\ : InMux
    port map (
            O => \N__24171\,
            I => \N__24168\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__24168\,
            I => \N__24165\
        );

    \I__3290\ : Span12Mux_h
    port map (
            O => \N__24165\,
            I => \N__24162\
        );

    \I__3289\ : Odrv12
    port map (
            O => \N__24162\,
            I => \pwm_generator_inst.un2_threshold_2_6\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24156\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__24156\,
            I => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\
        );

    \I__3286\ : InMux
    port map (
            O => \N__24153\,
            I => \pwm_generator_inst.un2_threshold_add_1_cry_5\
        );

    \I__3285\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24147\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__24147\,
            I => \N__24143\
        );

    \I__3283\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24140\
        );

    \I__3282\ : Odrv12
    port map (
            O => \N__24143\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__24140\,
            I => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\
        );

    \I__3280\ : CascadeMux
    port map (
            O => \N__24135\,
            I => \N__24132\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24129\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__24129\,
            I => \N__24126\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__24126\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24118\
        );

    \I__3275\ : InMux
    port map (
            O => \N__24122\,
            I => \N__24115\
        );

    \I__3274\ : InMux
    port map (
            O => \N__24121\,
            I => \N__24112\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__24118\,
            I => \N__24109\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24115\,
            I => \N__24106\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__24112\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__24109\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__24106\,
            I => \pwm_generator_inst.un15_threshold_1_axb_14\
        );

    \I__3268\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24096\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__24096\,
            I => \pwm_generator_inst.un19_threshold_axb_4\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24093\,
            I => \N__24089\
        );

    \I__3265\ : InMux
    port map (
            O => \N__24092\,
            I => \N__24086\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__24089\,
            I => \N__24083\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__24086\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__24083\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13\
        );

    \I__3261\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24075\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__24072\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__24072\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__24069\,
            I => \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__24066\,
            I => \N__24062\
        );

    \I__3256\ : InMux
    port map (
            O => \N__24065\,
            I => \N__24057\
        );

    \I__3255\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24057\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24054\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__24054\,
            I => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\
        );

    \I__3252\ : InMux
    port map (
            O => \N__24051\,
            I => \N__24048\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__24048\,
            I => \pwm_generator_inst.un19_threshold_axb_3\
        );

    \I__3250\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24042\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__24042\,
            I => \N__24039\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__24039\,
            I => \N__24036\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__24036\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\
        );

    \I__3246\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24030\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__24030\,
            I => \N__24027\
        );

    \I__3244\ : Span4Mux_v
    port map (
            O => \N__24027\,
            I => \N__24024\
        );

    \I__3243\ : Span4Mux_h
    port map (
            O => \N__24024\,
            I => \N__24021\
        );

    \I__3242\ : Odrv4
    port map (
            O => \N__24021\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\
        );

    \I__3241\ : InMux
    port map (
            O => \N__24018\,
            I => \N__24015\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24015\,
            I => \N__24012\
        );

    \I__3239\ : Span4Mux_h
    port map (
            O => \N__24012\,
            I => \N__24009\
        );

    \I__3238\ : Odrv4
    port map (
            O => \N__24009\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24006\,
            I => \pwm_generator_inst.un3_threshold_cry_19\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24003\,
            I => \N__24000\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__24000\,
            I => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\
        );

    \I__3234\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23994\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__23994\,
            I => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__23991\,
            I => \N__23988\
        );

    \I__3231\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23985\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__23985\,
            I => \N__23982\
        );

    \I__3229\ : Odrv4
    port map (
            O => \N__23982\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\
        );

    \I__3228\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23976\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__23976\,
            I => \N__23973\
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__23973\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__23970\,
            I => \N__23967\
        );

    \I__3224\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23962\
        );

    \I__3223\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23959\
        );

    \I__3222\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23956\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__23962\,
            I => \N__23953\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23950\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__23956\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__23953\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__23950\,
            I => \pwm_generator_inst.un15_threshold_1_axb_12\
        );

    \I__3216\ : InMux
    port map (
            O => \N__23943\,
            I => \N__23940\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__23940\,
            I => \N__23936\
        );

    \I__3214\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23933\
        );

    \I__3213\ : Odrv12
    port map (
            O => \N__23936\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__23933\,
            I => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\
        );

    \I__3211\ : InMux
    port map (
            O => \N__23928\,
            I => \N__23925\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__23925\,
            I => \pwm_generator_inst.un19_threshold_axb_2\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23919\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__23919\,
            I => \N__23916\
        );

    \I__3207\ : Span4Mux_h
    port map (
            O => \N__23916\,
            I => \N__23912\
        );

    \I__3206\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23909\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__23912\,
            I => \pwm_generator_inst.O_10\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__23909\,
            I => \pwm_generator_inst.O_10\
        );

    \I__3203\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23901\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__23901\,
            I => \N__23898\
        );

    \I__3201\ : Span4Mux_v
    port map (
            O => \N__23898\,
            I => \N__23894\
        );

    \I__3200\ : InMux
    port map (
            O => \N__23897\,
            I => \N__23890\
        );

    \I__3199\ : Span4Mux_h
    port map (
            O => \N__23894\,
            I => \N__23887\
        );

    \I__3198\ : InMux
    port map (
            O => \N__23893\,
            I => \N__23884\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__23890\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3196\ : Odrv4
    port map (
            O => \N__23887\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__23884\,
            I => \pwm_generator_inst.un15_threshold_1_axb_10\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__23877\,
            I => \N__23874\
        );

    \I__3193\ : InMux
    port map (
            O => \N__23874\,
            I => \N__23871\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__23871\,
            I => \N__23868\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__23868\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\
        );

    \I__3190\ : InMux
    port map (
            O => \N__23865\,
            I => \N__23862\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__23862\,
            I => \pwm_generator_inst.un19_threshold_axb_0\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__23859\,
            I => \N__23856\
        );

    \I__3187\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23853\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__23853\,
            I => \N__23850\
        );

    \I__3185\ : Span4Mux_h
    port map (
            O => \N__23850\,
            I => \N__23847\
        );

    \I__3184\ : Odrv4
    port map (
            O => \N__23847\,
            I => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\
        );

    \I__3183\ : InMux
    port map (
            O => \N__23844\,
            I => \bfn_4_23_0_\
        );

    \I__3182\ : InMux
    port map (
            O => \N__23841\,
            I => \N__23837\
        );

    \I__3181\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23834\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__23837\,
            I => \N__23831\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__23834\,
            I => \N__23828\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__23831\,
            I => \N__23825\
        );

    \I__3177\ : Span4Mux_v
    port map (
            O => \N__23828\,
            I => \N__23822\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__23825\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__23822\,
            I => \pwm_generator_inst.un3_threshold\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23817\,
            I => \N__23814\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__23814\,
            I => \N__23811\
        );

    \I__3172\ : Span4Mux_h
    port map (
            O => \N__23811\,
            I => \N__23808\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__23808\,
            I => \pwm_generator_inst.O_12\
        );

    \I__3170\ : InMux
    port map (
            O => \N__23805\,
            I => \pwm_generator_inst.un3_threshold_cry_0\
        );

    \I__3169\ : InMux
    port map (
            O => \N__23802\,
            I => \N__23799\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__23799\,
            I => \N__23796\
        );

    \I__3167\ : Span4Mux_v
    port map (
            O => \N__23796\,
            I => \N__23793\
        );

    \I__3166\ : Odrv4
    port map (
            O => \N__23793\,
            I => \pwm_generator_inst.O_13\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23790\,
            I => \pwm_generator_inst.un3_threshold_cry_1\
        );

    \I__3164\ : InMux
    port map (
            O => \N__23787\,
            I => \N__23784\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23781\
        );

    \I__3162\ : Span4Mux_h
    port map (
            O => \N__23781\,
            I => \N__23778\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__23778\,
            I => \pwm_generator_inst.O_14\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23775\,
            I => \pwm_generator_inst.un3_threshold_cry_2\
        );

    \I__3159\ : InMux
    port map (
            O => \N__23772\,
            I => \N__23769\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23766\
        );

    \I__3157\ : Span4Mux_h
    port map (
            O => \N__23766\,
            I => \N__23762\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23765\,
            I => \N__23759\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__23762\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__23759\,
            I => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\
        );

    \I__3153\ : InMux
    port map (
            O => \N__23754\,
            I => \pwm_generator_inst.un3_threshold_cry_3\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__23751\,
            I => \N__23747\
        );

    \I__3151\ : InMux
    port map (
            O => \N__23750\,
            I => \N__23742\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23742\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23742\,
            I => \N__23739\
        );

    \I__3148\ : Odrv4
    port map (
            O => \N__23739\,
            I => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\
        );

    \I__3147\ : InMux
    port map (
            O => \N__23736\,
            I => \pwm_generator_inst.un3_threshold_cry_4\
        );

    \I__3146\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23730\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__23730\,
            I => \N__23726\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23723\
        );

    \I__3143\ : Odrv4
    port map (
            O => \N__23726\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__23723\,
            I => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23718\,
            I => \pwm_generator_inst.un3_threshold_cry_5\
        );

    \I__3140\ : InMux
    port map (
            O => \N__23715\,
            I => \N__23711\
        );

    \I__3139\ : InMux
    port map (
            O => \N__23714\,
            I => \N__23708\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__23711\,
            I => \N__23705\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23708\,
            I => \N__23702\
        );

    \I__3136\ : Span4Mux_v
    port map (
            O => \N__23705\,
            I => \N__23699\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__23702\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__23699\,
            I => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23694\,
            I => \pwm_generator_inst.un3_threshold_cry_6\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__23691\,
            I => \N__23688\
        );

    \I__3131\ : InMux
    port map (
            O => \N__23688\,
            I => \N__23685\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23685\,
            I => \N__23682\
        );

    \I__3129\ : Odrv4
    port map (
            O => \N__23682\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23679\,
            I => \N__23676\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__23676\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\
        );

    \I__3126\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23670\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23670\,
            I => \N__23667\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__23667\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\
        );

    \I__3123\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23661\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__23661\,
            I => \N__23658\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__23658\,
            I => \N__23655\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__23655\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\
        );

    \I__3119\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23649\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23649\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\
        );

    \I__3117\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__23643\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23637\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__23637\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__23634\,
            I => \N__23631\
        );

    \I__3112\ : InMux
    port map (
            O => \N__23631\,
            I => \N__23628\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23628\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\
        );

    \I__3110\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__23622\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23619\,
            I => \N__23616\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__3106\ : Span4Mux_v
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__23610\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23604\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__23604\,
            I => \N__23601\
        );

    \I__3102\ : Odrv4
    port map (
            O => \N__23601\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23594\
        );

    \I__3100\ : InMux
    port map (
            O => \N__23597\,
            I => \N__23575\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__23594\,
            I => \N__23572\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23593\,
            I => \N__23567\
        );

    \I__3097\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23567\
        );

    \I__3096\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23564\
        );

    \I__3095\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23561\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23589\,
            I => \N__23556\
        );

    \I__3093\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23556\
        );

    \I__3092\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23553\
        );

    \I__3091\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23549\
        );

    \I__3090\ : InMux
    port map (
            O => \N__23585\,
            I => \N__23534\
        );

    \I__3089\ : InMux
    port map (
            O => \N__23584\,
            I => \N__23534\
        );

    \I__3088\ : InMux
    port map (
            O => \N__23583\,
            I => \N__23534\
        );

    \I__3087\ : InMux
    port map (
            O => \N__23582\,
            I => \N__23534\
        );

    \I__3086\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23534\
        );

    \I__3085\ : InMux
    port map (
            O => \N__23580\,
            I => \N__23534\
        );

    \I__3084\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23534\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23531\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23575\,
            I => \N__23510\
        );

    \I__3081\ : Span4Mux_h
    port map (
            O => \N__23572\,
            I => \N__23510\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__23567\,
            I => \N__23510\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__23564\,
            I => \N__23510\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23507\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23556\,
            I => \N__23501\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__23553\,
            I => \N__23501\
        );

    \I__3075\ : InMux
    port map (
            O => \N__23552\,
            I => \N__23498\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__23549\,
            I => \N__23491\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23491\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__23531\,
            I => \N__23491\
        );

    \I__3071\ : InMux
    port map (
            O => \N__23530\,
            I => \N__23488\
        );

    \I__3070\ : InMux
    port map (
            O => \N__23529\,
            I => \N__23477\
        );

    \I__3069\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23477\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23477\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23526\,
            I => \N__23477\
        );

    \I__3066\ : InMux
    port map (
            O => \N__23525\,
            I => \N__23477\
        );

    \I__3065\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23474\
        );

    \I__3064\ : InMux
    port map (
            O => \N__23523\,
            I => \N__23463\
        );

    \I__3063\ : InMux
    port map (
            O => \N__23522\,
            I => \N__23463\
        );

    \I__3062\ : InMux
    port map (
            O => \N__23521\,
            I => \N__23463\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23463\
        );

    \I__3060\ : InMux
    port map (
            O => \N__23519\,
            I => \N__23463\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__23510\,
            I => \N__23458\
        );

    \I__3058\ : Span4Mux_v
    port map (
            O => \N__23507\,
            I => \N__23458\
        );

    \I__3057\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23455\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__23501\,
            I => \N__23450\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__23498\,
            I => \N__23450\
        );

    \I__3054\ : Span4Mux_v
    port map (
            O => \N__23491\,
            I => \N__23445\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__23488\,
            I => \N__23445\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__23477\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23474\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__23463\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3049\ : Odrv4
    port map (
            O => \N__23458\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__23455\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3047\ : Odrv4
    port map (
            O => \N__23450\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__23445\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_31\
        );

    \I__3045\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23412\
        );

    \I__3044\ : InMux
    port map (
            O => \N__23429\,
            I => \N__23412\
        );

    \I__3043\ : InMux
    port map (
            O => \N__23428\,
            I => \N__23409\
        );

    \I__3042\ : InMux
    port map (
            O => \N__23427\,
            I => \N__23406\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23426\,
            I => \N__23391\
        );

    \I__3040\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23391\
        );

    \I__3039\ : InMux
    port map (
            O => \N__23424\,
            I => \N__23391\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23423\,
            I => \N__23391\
        );

    \I__3037\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23391\
        );

    \I__3036\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23391\
        );

    \I__3035\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23391\
        );

    \I__3034\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23382\
        );

    \I__3033\ : InMux
    port map (
            O => \N__23418\,
            I => \N__23382\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__23417\,
            I => \N__23375\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__23412\,
            I => \N__23366\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23359\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__23406\,
            I => \N__23359\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23359\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23390\,
            I => \N__23352\
        );

    \I__3026\ : InMux
    port map (
            O => \N__23389\,
            I => \N__23352\
        );

    \I__3025\ : InMux
    port map (
            O => \N__23388\,
            I => \N__23352\
        );

    \I__3024\ : InMux
    port map (
            O => \N__23387\,
            I => \N__23349\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__23382\,
            I => \N__23346\
        );

    \I__3022\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23341\
        );

    \I__3021\ : InMux
    port map (
            O => \N__23380\,
            I => \N__23341\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__23379\,
            I => \N__23335\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__23378\,
            I => \N__23332\
        );

    \I__3018\ : InMux
    port map (
            O => \N__23375\,
            I => \N__23329\
        );

    \I__3017\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23318\
        );

    \I__3016\ : InMux
    port map (
            O => \N__23373\,
            I => \N__23318\
        );

    \I__3015\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23318\
        );

    \I__3014\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23318\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23318\
        );

    \I__3012\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23315\
        );

    \I__3011\ : Span4Mux_h
    port map (
            O => \N__23366\,
            I => \N__23312\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__23359\,
            I => \N__23305\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__23352\,
            I => \N__23305\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23305\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__23346\,
            I => \N__23300\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__23341\,
            I => \N__23300\
        );

    \I__3005\ : InMux
    port map (
            O => \N__23340\,
            I => \N__23289\
        );

    \I__3004\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23289\
        );

    \I__3003\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23289\
        );

    \I__3002\ : InMux
    port map (
            O => \N__23335\,
            I => \N__23289\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23332\,
            I => \N__23289\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__23329\,
            I => \N__23284\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23284\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23279\
        );

    \I__2997\ : Span4Mux_v
    port map (
            O => \N__23312\,
            I => \N__23279\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__23305\,
            I => \N__23276\
        );

    \I__2995\ : Span4Mux_v
    port map (
            O => \N__23300\,
            I => \N__23273\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__23289\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__23284\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__23279\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__23276\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__23273\,
            I => \current_shift_inst.PI_CTRL.N_47\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__2988\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23256\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__2986\ : Span4Mux_h
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__23250\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__23247\,
            I => \N__23234\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__23246\,
            I => \N__23231\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__23245\,
            I => \N__23227\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__23244\,
            I => \N__23224\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__23243\,
            I => \N__23218\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__23242\,
            I => \N__23214\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__23241\,
            I => \N__23209\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__23240\,
            I => \N__23197\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__23239\,
            I => \N__23193\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__23238\,
            I => \N__23190\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__23237\,
            I => \N__23187\
        );

    \I__2973\ : InMux
    port map (
            O => \N__23234\,
            I => \N__23182\
        );

    \I__2972\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23182\
        );

    \I__2971\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23179\
        );

    \I__2970\ : InMux
    port map (
            O => \N__23227\,
            I => \N__23172\
        );

    \I__2969\ : InMux
    port map (
            O => \N__23224\,
            I => \N__23172\
        );

    \I__2968\ : InMux
    port map (
            O => \N__23223\,
            I => \N__23172\
        );

    \I__2967\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23167\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23221\,
            I => \N__23167\
        );

    \I__2965\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23164\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23159\
        );

    \I__2963\ : InMux
    port map (
            O => \N__23214\,
            I => \N__23159\
        );

    \I__2962\ : InMux
    port map (
            O => \N__23213\,
            I => \N__23152\
        );

    \I__2961\ : InMux
    port map (
            O => \N__23212\,
            I => \N__23152\
        );

    \I__2960\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23152\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__23208\,
            I => \N__23146\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__23207\,
            I => \N__23143\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__23206\,
            I => \N__23140\
        );

    \I__2956\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23137\
        );

    \I__2955\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23126\
        );

    \I__2954\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23126\
        );

    \I__2953\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23126\
        );

    \I__2952\ : InMux
    port map (
            O => \N__23201\,
            I => \N__23126\
        );

    \I__2951\ : InMux
    port map (
            O => \N__23200\,
            I => \N__23126\
        );

    \I__2950\ : InMux
    port map (
            O => \N__23197\,
            I => \N__23123\
        );

    \I__2949\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23114\
        );

    \I__2948\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23114\
        );

    \I__2947\ : InMux
    port map (
            O => \N__23190\,
            I => \N__23114\
        );

    \I__2946\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23114\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__23182\,
            I => \N__23111\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__23179\,
            I => \N__23108\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23105\
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__23167\,
            I => \N__23096\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__23164\,
            I => \N__23096\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__23159\,
            I => \N__23096\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__23152\,
            I => \N__23096\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23151\,
            I => \N__23093\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23150\,
            I => \N__23082\
        );

    \I__2936\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23082\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23146\,
            I => \N__23082\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23143\,
            I => \N__23082\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23082\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23137\,
            I => \N__23079\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__23076\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__23123\,
            I => \N__23067\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__23114\,
            I => \N__23067\
        );

    \I__2928\ : Span4Mux_h
    port map (
            O => \N__23111\,
            I => \N__23067\
        );

    \I__2927\ : Span4Mux_s3_h
    port map (
            O => \N__23108\,
            I => \N__23067\
        );

    \I__2926\ : Span4Mux_s3_h
    port map (
            O => \N__23105\,
            I => \N__23062\
        );

    \I__2925\ : Span4Mux_v
    port map (
            O => \N__23096\,
            I => \N__23062\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__23093\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__23082\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__23079\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__23076\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__23067\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__23062\,
            I => \current_shift_inst.PI_CTRL.N_46\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23046\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__23046\,
            I => \N__23043\
        );

    \I__2916\ : Odrv4
    port map (
            O => \N__23043\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\
        );

    \I__2915\ : InMux
    port map (
            O => \N__23040\,
            I => \N__23037\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__23037\,
            I => \N__23034\
        );

    \I__2913\ : Span4Mux_v
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__2912\ : Odrv4
    port map (
            O => \N__23031\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\
        );

    \I__2911\ : InMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__23025\,
            I => \N__23022\
        );

    \I__2909\ : Span4Mux_v
    port map (
            O => \N__23022\,
            I => \N__23019\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__23019\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__23016\,
            I => \N__23013\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23009\
        );

    \I__2905\ : InMux
    port map (
            O => \N__23012\,
            I => \N__23004\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23001\
        );

    \I__2903\ : InMux
    port map (
            O => \N__23008\,
            I => \N__22998\
        );

    \I__2902\ : InMux
    port map (
            O => \N__23007\,
            I => \N__22995\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__23004\,
            I => \N__22992\
        );

    \I__2900\ : Span4Mux_v
    port map (
            O => \N__23001\,
            I => \N__22987\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__22998\,
            I => \N__22987\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__22995\,
            I => \N__22984\
        );

    \I__2897\ : Odrv4
    port map (
            O => \N__22992\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__22987\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__22984\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_15\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__22977\,
            I => \N__22974\
        );

    \I__2893\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22970\
        );

    \I__2892\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22966\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__22970\,
            I => \N__22962\
        );

    \I__2890\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22959\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22956\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22965\,
            I => \N__22953\
        );

    \I__2887\ : Span4Mux_v
    port map (
            O => \N__22962\,
            I => \N__22946\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__22959\,
            I => \N__22946\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__22956\,
            I => \N__22946\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__22953\,
            I => \N__22943\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__22946\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2882\ : Odrv12
    port map (
            O => \N__22943\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_13\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__2880\ : InMux
    port map (
            O => \N__22935\,
            I => \N__22930\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__22934\,
            I => \N__22927\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__22933\,
            I => \N__22924\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22921\
        );

    \I__2876\ : InMux
    port map (
            O => \N__22927\,
            I => \N__22918\
        );

    \I__2875\ : InMux
    port map (
            O => \N__22924\,
            I => \N__22914\
        );

    \I__2874\ : Span12Mux_s3_h
    port map (
            O => \N__22921\,
            I => \N__22909\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__22918\,
            I => \N__22909\
        );

    \I__2872\ : InMux
    port map (
            O => \N__22917\,
            I => \N__22906\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__22914\,
            I => \N__22903\
        );

    \I__2870\ : Span12Mux_v
    port map (
            O => \N__22909\,
            I => \N__22900\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__22906\,
            I => \N__22897\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__22903\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2867\ : Odrv12
    port map (
            O => \N__22900\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2866\ : Odrv4
    port map (
            O => \N__22897\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_10\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__22884\,
            I => \N__22878\
        );

    \I__2862\ : InMux
    port map (
            O => \N__22883\,
            I => \N__22875\
        );

    \I__2861\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22872\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22881\,
            I => \N__22869\
        );

    \I__2859\ : Span4Mux_h
    port map (
            O => \N__22878\,
            I => \N__22864\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22864\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__22872\,
            I => \N__22861\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22869\,
            I => \N__22858\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__22864\,
            I => \N__22853\
        );

    \I__2854\ : Span4Mux_v
    port map (
            O => \N__22861\,
            I => \N__22853\
        );

    \I__2853\ : Odrv4
    port map (
            O => \N__22858\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__22853\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_16\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22848\,
            I => \N__22845\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__22845\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\
        );

    \I__2849\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22839\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__22839\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22836\,
            I => \N__22833\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22833\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\
        );

    \I__2845\ : InMux
    port map (
            O => \N__22830\,
            I => \bfn_3_25_0_\
        );

    \I__2844\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22824\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__22824\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\
        );

    \I__2842\ : InMux
    port map (
            O => \N__22821\,
            I => \pwm_generator_inst.un19_threshold_cry_8\
        );

    \I__2841\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22815\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__22815\,
            I => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\
        );

    \I__2839\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22805\
        );

    \I__2838\ : InMux
    port map (
            O => \N__22811\,
            I => \N__22805\
        );

    \I__2837\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22802\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__22805\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__22802\,
            I => \pwm_generator_inst.un15_threshold_1_axb_16\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22794\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__22794\,
            I => \pwm_generator_inst.un19_threshold_axb_6\
        );

    \I__2832\ : InMux
    port map (
            O => \N__22791\,
            I => \N__22788\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__22788\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\
        );

    \I__2830\ : InMux
    port map (
            O => \N__22785\,
            I => \N__22780\
        );

    \I__2829\ : InMux
    port map (
            O => \N__22784\,
            I => \N__22777\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22774\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__22780\,
            I => \N__22769\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22777\,
            I => \N__22769\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__22774\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2824\ : Odrv4
    port map (
            O => \N__22769\,
            I => \pwm_generator_inst.un15_threshold_1_axb_15\
        );

    \I__2823\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22761\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22761\,
            I => \pwm_generator_inst.un19_threshold_axb_5\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22758\,
            I => \N__22751\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22757\,
            I => \N__22751\
        );

    \I__2819\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22748\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22751\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__22748\,
            I => \pwm_generator_inst.un15_threshold_1_axb_18\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__22743\,
            I => \N__22740\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22737\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__22737\,
            I => \N__22734\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__22734\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\
        );

    \I__2812\ : InMux
    port map (
            O => \N__22731\,
            I => \N__22728\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__22728\,
            I => \pwm_generator_inst.un19_threshold_axb_8\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22722\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22722\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\
        );

    \I__2808\ : InMux
    port map (
            O => \N__22719\,
            I => \N__22714\
        );

    \I__2807\ : InMux
    port map (
            O => \N__22718\,
            I => \N__22711\
        );

    \I__2806\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22708\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__22714\,
            I => \N__22705\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__22711\,
            I => \N__22702\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__22708\,
            I => \N__22697\
        );

    \I__2802\ : Span4Mux_v
    port map (
            O => \N__22705\,
            I => \N__22697\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__22702\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__22697\,
            I => \pwm_generator_inst.un15_threshold_1_axb_17\
        );

    \I__2799\ : InMux
    port map (
            O => \N__22692\,
            I => \N__22689\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__22689\,
            I => \pwm_generator_inst.un19_threshold_axb_7\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22686\,
            I => \N__22683\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__22680\,
            I => \N__22677\
        );

    \I__2794\ : Span4Mux_h
    port map (
            O => \N__22677\,
            I => \N__22674\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__22674\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__22671\,
            I => \N__22665\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__22670\,
            I => \N__22662\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22669\,
            I => \N__22659\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22668\,
            I => \N__22656\
        );

    \I__2788\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22653\
        );

    \I__2787\ : InMux
    port map (
            O => \N__22662\,
            I => \N__22650\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22659\,
            I => \N__22643\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22643\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22643\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__22650\,
            I => \N__22640\
        );

    \I__2782\ : Span4Mux_v
    port map (
            O => \N__22643\,
            I => \N__22637\
        );

    \I__2781\ : Span4Mux_v
    port map (
            O => \N__22640\,
            I => \N__22634\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__22637\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__22634\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_5\
        );

    \I__2778\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__22626\,
            I => \pwm_generator_inst.un19_threshold_axb_1\
        );

    \I__2776\ : InMux
    port map (
            O => \N__22623\,
            I => \pwm_generator_inst.un19_threshold_cry_0\
        );

    \I__2775\ : InMux
    port map (
            O => \N__22620\,
            I => \pwm_generator_inst.un19_threshold_cry_1\
        );

    \I__2774\ : InMux
    port map (
            O => \N__22617\,
            I => \pwm_generator_inst.un19_threshold_cry_2\
        );

    \I__2773\ : InMux
    port map (
            O => \N__22614\,
            I => \pwm_generator_inst.un19_threshold_cry_3\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22611\,
            I => \pwm_generator_inst.un19_threshold_cry_4\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22608\,
            I => \pwm_generator_inst.un19_threshold_cry_5\
        );

    \I__2770\ : InMux
    port map (
            O => \N__22605\,
            I => \pwm_generator_inst.un19_threshold_cry_6\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__2768\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__22596\,
            I => \N__22591\
        );

    \I__2766\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22587\
        );

    \I__2765\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22584\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__22591\,
            I => \N__22581\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22590\,
            I => \N__22578\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__22587\,
            I => \N__22575\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22572\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__22581\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__22578\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2758\ : Odrv12
    port map (
            O => \N__22575\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2757\ : Odrv4
    port map (
            O => \N__22572\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_30\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__22563\,
            I => \N__22559\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__22562\,
            I => \N__22556\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22551\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22551\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__22551\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\
        );

    \I__2751\ : InMux
    port map (
            O => \N__22548\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\
        );

    \I__2750\ : InMux
    port map (
            O => \N__22545\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\
        );

    \I__2749\ : InMux
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__22539\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\
        );

    \I__2747\ : InMux
    port map (
            O => \N__22536\,
            I => \N__22533\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22530\
        );

    \I__2745\ : Odrv12
    port map (
            O => \N__22530\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\
        );

    \I__2744\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22524\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__22524\,
            I => \N__22521\
        );

    \I__2742\ : Span4Mux_s3_h
    port map (
            O => \N__22521\,
            I => \N__22518\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__22518\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__22515\,
            I => \N__22512\
        );

    \I__2739\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22508\
        );

    \I__2738\ : InMux
    port map (
            O => \N__22511\,
            I => \N__22505\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__22508\,
            I => \N__22501\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__22505\,
            I => \N__22498\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22495\
        );

    \I__2734\ : Span12Mux_s3_h
    port map (
            O => \N__22501\,
            I => \N__22488\
        );

    \I__2733\ : Sp12to4
    port map (
            O => \N__22498\,
            I => \N__22488\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__22495\,
            I => \N__22488\
        );

    \I__2731\ : Odrv12
    port map (
            O => \N__22488\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22485\,
            I => \N__22481\
        );

    \I__2729\ : InMux
    port map (
            O => \N__22484\,
            I => \N__22477\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__22481\,
            I => \N__22474\
        );

    \I__2727\ : InMux
    port map (
            O => \N__22480\,
            I => \N__22471\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__22477\,
            I => \N__22468\
        );

    \I__2725\ : Span4Mux_h
    port map (
            O => \N__22474\,
            I => \N__22463\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22463\
        );

    \I__2723\ : Span4Mux_v
    port map (
            O => \N__22468\,
            I => \N__22458\
        );

    \I__2722\ : Span4Mux_v
    port map (
            O => \N__22463\,
            I => \N__22458\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__22458\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__22455\,
            I => \N__22452\
        );

    \I__2719\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22449\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__22449\,
            I => \N__22444\
        );

    \I__2717\ : InMux
    port map (
            O => \N__22448\,
            I => \N__22441\
        );

    \I__2716\ : InMux
    port map (
            O => \N__22447\,
            I => \N__22438\
        );

    \I__2715\ : Span4Mux_v
    port map (
            O => \N__22444\,
            I => \N__22433\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22433\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__22438\,
            I => \N__22430\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__22433\,
            I => \N__22427\
        );

    \I__2711\ : Odrv12
    port map (
            O => \N__22430\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__22427\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__22422\,
            I => \N__22419\
        );

    \I__2708\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22416\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22416\,
            I => \N__22411\
        );

    \I__2706\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22408\
        );

    \I__2705\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22405\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__22411\,
            I => \N__22400\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22400\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__22405\,
            I => \N__22397\
        );

    \I__2701\ : Span4Mux_v
    port map (
            O => \N__22400\,
            I => \N__22394\
        );

    \I__2700\ : Odrv12
    port map (
            O => \N__22397\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2699\ : Odrv4
    port map (
            O => \N__22394\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__22389\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22379\
        );

    \I__2695\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22376\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__22379\,
            I => \N__22372\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22369\
        );

    \I__2692\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22366\
        );

    \I__2691\ : Span4Mux_v
    port map (
            O => \N__22372\,
            I => \N__22363\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__22369\,
            I => \N__22358\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__22366\,
            I => \N__22358\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__22363\,
            I => \N__22355\
        );

    \I__2687\ : Span4Mux_v
    port map (
            O => \N__22358\,
            I => \N__22352\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__22355\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__22352\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__22347\,
            I => \N__22344\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22337\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22334\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__22337\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__22334\,
            I => \current_shift_inst.PI_CTRL.N_27\
        );

    \I__2678\ : InMux
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__2676\ : Odrv12
    port map (
            O => \N__22323\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__22320\,
            I => \N__22317\
        );

    \I__2674\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22312\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__22316\,
            I => \N__22309\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__22315\,
            I => \N__22306\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__22312\,
            I => \N__22303\
        );

    \I__2670\ : InMux
    port map (
            O => \N__22309\,
            I => \N__22299\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22296\
        );

    \I__2668\ : Span4Mux_v
    port map (
            O => \N__22303\,
            I => \N__22293\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22290\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__22299\,
            I => \N__22287\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22284\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__22293\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__22290\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2662\ : Odrv4
    port map (
            O => \N__22287\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2661\ : Odrv12
    port map (
            O => \N__22284\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_22\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__22275\,
            I => \N__22272\
        );

    \I__2659\ : InMux
    port map (
            O => \N__22272\,
            I => \N__22269\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__22269\,
            I => \N__22266\
        );

    \I__2657\ : Span4Mux_v
    port map (
            O => \N__22266\,
            I => \N__22262\
        );

    \I__2656\ : InMux
    port map (
            O => \N__22265\,
            I => \N__22259\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__22262\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__22259\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\
        );

    \I__2653\ : InMux
    port map (
            O => \N__22254\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\
        );

    \I__2652\ : CascadeMux
    port map (
            O => \N__22251\,
            I => \N__22248\
        );

    \I__2651\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22244\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__22247\,
            I => \N__22241\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22244\,
            I => \N__22236\
        );

    \I__2648\ : InMux
    port map (
            O => \N__22241\,
            I => \N__22233\
        );

    \I__2647\ : InMux
    port map (
            O => \N__22240\,
            I => \N__22230\
        );

    \I__2646\ : InMux
    port map (
            O => \N__22239\,
            I => \N__22227\
        );

    \I__2645\ : Span4Mux_v
    port map (
            O => \N__22236\,
            I => \N__22224\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__22233\,
            I => \N__22219\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__22230\,
            I => \N__22219\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22216\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__22224\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__22219\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2639\ : Odrv12
    port map (
            O => \N__22216\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_23\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__22209\,
            I => \N__22205\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__22208\,
            I => \N__22202\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22197\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22197\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__22197\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\
        );

    \I__2633\ : InMux
    port map (
            O => \N__22194\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22187\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__22190\,
            I => \N__22183\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22179\
        );

    \I__2629\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22176\
        );

    \I__2628\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22173\
        );

    \I__2627\ : InMux
    port map (
            O => \N__22182\,
            I => \N__22170\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__22179\,
            I => \N__22165\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__22176\,
            I => \N__22165\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__22173\,
            I => \N__22162\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__22170\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__22165\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__22162\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_24\
        );

    \I__2620\ : InMux
    port map (
            O => \N__22155\,
            I => \N__22149\
        );

    \I__2619\ : InMux
    port map (
            O => \N__22154\,
            I => \N__22149\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__22149\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\
        );

    \I__2617\ : InMux
    port map (
            O => \N__22146\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__22143\,
            I => \N__22140\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22140\,
            I => \N__22137\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__22137\,
            I => \N__22132\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__22136\,
            I => \N__22129\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22125\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__22132\,
            I => \N__22122\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22119\
        );

    \I__2609\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22116\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__22125\,
            I => \N__22113\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__22122\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__22119\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__22116\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2604\ : Odrv12
    port map (
            O => \N__22113\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_25\
        );

    \I__2603\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22101\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22101\,
            I => \N__22097\
        );

    \I__2601\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22094\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__22097\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__22094\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\
        );

    \I__2598\ : InMux
    port map (
            O => \N__22089\,
            I => \bfn_3_20_0_\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__22086\,
            I => \N__22083\
        );

    \I__2596\ : InMux
    port map (
            O => \N__22083\,
            I => \N__22080\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22077\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__22077\,
            I => \N__22072\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22069\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22075\,
            I => \N__22065\
        );

    \I__2591\ : Sp12to4
    port map (
            O => \N__22072\,
            I => \N__22060\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__22069\,
            I => \N__22060\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22068\,
            I => \N__22057\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__22065\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2587\ : Odrv12
    port map (
            O => \N__22060\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__22057\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_26\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22050\,
            I => \N__22046\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__22049\,
            I => \N__22043\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__22046\,
            I => \N__22040\
        );

    \I__2582\ : InMux
    port map (
            O => \N__22043\,
            I => \N__22037\
        );

    \I__2581\ : Odrv4
    port map (
            O => \N__22040\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__22037\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22032\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__22029\,
            I => \N__22026\
        );

    \I__2577\ : InMux
    port map (
            O => \N__22026\,
            I => \N__22023\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__22023\,
            I => \N__22020\
        );

    \I__2575\ : Span4Mux_h
    port map (
            O => \N__22020\,
            I => \N__22014\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22019\,
            I => \N__22011\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22018\,
            I => \N__22008\
        );

    \I__2572\ : InMux
    port map (
            O => \N__22017\,
            I => \N__22005\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__22014\,
            I => \N__22000\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__22011\,
            I => \N__22000\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__21997\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__22005\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__22000\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__21997\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_27\
        );

    \I__2565\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21984\
        );

    \I__2564\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21984\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__21984\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\
        );

    \I__2562\ : InMux
    port map (
            O => \N__21981\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\
        );

    \I__2561\ : CascadeMux
    port map (
            O => \N__21978\,
            I => \N__21975\
        );

    \I__2560\ : InMux
    port map (
            O => \N__21975\,
            I => \N__21971\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__21974\,
            I => \N__21967\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__21971\,
            I => \N__21964\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__21970\,
            I => \N__21960\
        );

    \I__2556\ : InMux
    port map (
            O => \N__21967\,
            I => \N__21957\
        );

    \I__2555\ : Span4Mux_v
    port map (
            O => \N__21964\,
            I => \N__21954\
        );

    \I__2554\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21951\
        );

    \I__2553\ : InMux
    port map (
            O => \N__21960\,
            I => \N__21948\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__21957\,
            I => \N__21945\
        );

    \I__2551\ : Odrv4
    port map (
            O => \N__21954\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__21951\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__21948\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__21945\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_28\
        );

    \I__2547\ : InMux
    port map (
            O => \N__21936\,
            I => \N__21932\
        );

    \I__2546\ : InMux
    port map (
            O => \N__21935\,
            I => \N__21929\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__21932\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__21929\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\
        );

    \I__2543\ : InMux
    port map (
            O => \N__21924\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__21921\,
            I => \N__21918\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21915\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21912\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__21912\,
            I => \N__21909\
        );

    \I__2538\ : Span4Mux_v
    port map (
            O => \N__21909\,
            I => \N__21903\
        );

    \I__2537\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21900\
        );

    \I__2536\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21895\
        );

    \I__2535\ : InMux
    port map (
            O => \N__21906\,
            I => \N__21895\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__21903\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__21900\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__21895\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_29\
        );

    \I__2531\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21882\
        );

    \I__2530\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21882\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21882\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\
        );

    \I__2528\ : InMux
    port map (
            O => \N__21879\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__2526\ : InMux
    port map (
            O => \N__21873\,
            I => \N__21869\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21872\,
            I => \N__21865\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21869\,
            I => \N__21862\
        );

    \I__2523\ : InMux
    port map (
            O => \N__21868\,
            I => \N__21859\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__21865\,
            I => \N__21853\
        );

    \I__2521\ : Span4Mux_v
    port map (
            O => \N__21862\,
            I => \N__21853\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__21859\,
            I => \N__21850\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21858\,
            I => \N__21847\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__21853\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__21850\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__21847\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_14\
        );

    \I__2515\ : InMux
    port map (
            O => \N__21840\,
            I => \N__21834\
        );

    \I__2514\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21834\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21834\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\
        );

    \I__2512\ : InMux
    port map (
            O => \N__21831\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21828\,
            I => \N__21825\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__21825\,
            I => \N__21822\
        );

    \I__2509\ : Span4Mux_s3_h
    port map (
            O => \N__21822\,
            I => \N__21818\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21821\,
            I => \N__21815\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__21818\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__21815\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\
        );

    \I__2505\ : InMux
    port map (
            O => \N__21810\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\
        );

    \I__2504\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21804\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21801\
        );

    \I__2502\ : Span4Mux_s3_h
    port map (
            O => \N__21801\,
            I => \N__21797\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21800\,
            I => \N__21794\
        );

    \I__2500\ : Odrv4
    port map (
            O => \N__21797\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21794\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\
        );

    \I__2498\ : InMux
    port map (
            O => \N__21789\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__21786\,
            I => \N__21783\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21783\,
            I => \N__21780\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21780\,
            I => \N__21775\
        );

    \I__2494\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21771\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21768\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__21775\,
            I => \N__21765\
        );

    \I__2491\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21762\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__21771\,
            I => \N__21757\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__21768\,
            I => \N__21757\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__21765\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__21762\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2486\ : Odrv12
    port map (
            O => \N__21757\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_17\
        );

    \I__2485\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21744\
        );

    \I__2484\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21744\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__21744\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21741\,
            I => \bfn_3_19_0_\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21735\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__21732\,
            I => \N__21729\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__21729\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__21726\,
            I => \N__21723\
        );

    \I__2476\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21720\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__21720\,
            I => \N__21714\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21711\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21708\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21705\
        );

    \I__2471\ : Span4Mux_v
    port map (
            O => \N__21714\,
            I => \N__21700\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21711\,
            I => \N__21700\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21708\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__21705\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__21700\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_18\
        );

    \I__2466\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21689\
        );

    \I__2465\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21686\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__21689\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__21686\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\
        );

    \I__2462\ : InMux
    port map (
            O => \N__21681\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__21678\,
            I => \N__21675\
        );

    \I__2460\ : InMux
    port map (
            O => \N__21675\,
            I => \N__21671\
        );

    \I__2459\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21667\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21664\
        );

    \I__2457\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21660\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__21667\,
            I => \N__21657\
        );

    \I__2455\ : Span4Mux_v
    port map (
            O => \N__21664\,
            I => \N__21654\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21651\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__21660\,
            I => \N__21646\
        );

    \I__2452\ : Span4Mux_v
    port map (
            O => \N__21657\,
            I => \N__21646\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__21654\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__21651\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__21646\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_19\
        );

    \I__2448\ : InMux
    port map (
            O => \N__21639\,
            I => \N__21635\
        );

    \I__2447\ : InMux
    port map (
            O => \N__21638\,
            I => \N__21632\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__21635\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__21632\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\
        );

    \I__2444\ : InMux
    port map (
            O => \N__21627\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\
        );

    \I__2443\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21621\,
            I => \N__21615\
        );

    \I__2441\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21612\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__21619\,
            I => \N__21609\
        );

    \I__2439\ : InMux
    port map (
            O => \N__21618\,
            I => \N__21606\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__21615\,
            I => \N__21601\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__21612\,
            I => \N__21601\
        );

    \I__2436\ : InMux
    port map (
            O => \N__21609\,
            I => \N__21598\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__21606\,
            I => \N__21595\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__21601\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__21598\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2432\ : Odrv12
    port map (
            O => \N__21595\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_20\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__21588\,
            I => \N__21585\
        );

    \I__2430\ : InMux
    port map (
            O => \N__21585\,
            I => \N__21581\
        );

    \I__2429\ : InMux
    port map (
            O => \N__21584\,
            I => \N__21578\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__21581\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__21578\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\
        );

    \I__2426\ : InMux
    port map (
            O => \N__21573\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__21570\,
            I => \N__21567\
        );

    \I__2424\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21563\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__21566\,
            I => \N__21560\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__21563\,
            I => \N__21555\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21552\
        );

    \I__2420\ : InMux
    port map (
            O => \N__21559\,
            I => \N__21549\
        );

    \I__2419\ : InMux
    port map (
            O => \N__21558\,
            I => \N__21546\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__21555\,
            I => \N__21541\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__21552\,
            I => \N__21541\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__21549\,
            I => \N__21538\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__21546\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__21541\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__21538\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_21\
        );

    \I__2412\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21525\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21525\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__21525\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\
        );

    \I__2409\ : InMux
    port map (
            O => \N__21522\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\
        );

    \I__2408\ : InMux
    port map (
            O => \N__21519\,
            I => \N__21516\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__21516\,
            I => \N__21513\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__21513\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__21510\,
            I => \N__21505\
        );

    \I__2404\ : InMux
    port map (
            O => \N__21509\,
            I => \N__21502\
        );

    \I__2403\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21499\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21505\,
            I => \N__21496\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__21502\,
            I => \N__21492\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21499\,
            I => \N__21487\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__21496\,
            I => \N__21487\
        );

    \I__2398\ : InMux
    port map (
            O => \N__21495\,
            I => \N__21484\
        );

    \I__2397\ : Span4Mux_s3_h
    port map (
            O => \N__21492\,
            I => \N__21481\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__21487\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__21484\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2394\ : Odrv4
    port map (
            O => \N__21481\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_6\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21474\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__21471\,
            I => \N__21466\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__21470\,
            I => \N__21463\
        );

    \I__2390\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21460\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21466\,
            I => \N__21457\
        );

    \I__2388\ : InMux
    port map (
            O => \N__21463\,
            I => \N__21454\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__21460\,
            I => \N__21446\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21457\,
            I => \N__21446\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__21454\,
            I => \N__21446\
        );

    \I__2384\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21443\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__21446\,
            I => \N__21440\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21443\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__21440\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_7\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21435\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21427\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \N__21424\
        );

    \I__2377\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21420\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21417\
        );

    \I__2375\ : InMux
    port map (
            O => \N__21424\,
            I => \N__21414\
        );

    \I__2374\ : InMux
    port map (
            O => \N__21423\,
            I => \N__21411\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21408\
        );

    \I__2372\ : Sp12to4
    port map (
            O => \N__21417\,
            I => \N__21401\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__21414\,
            I => \N__21401\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21401\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__21408\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2368\ : Odrv12
    port map (
            O => \N__21401\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_8\
        );

    \I__2367\ : InMux
    port map (
            O => \N__21396\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\
        );

    \I__2366\ : InMux
    port map (
            O => \N__21393\,
            I => \N__21390\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__21390\,
            I => \N__21387\
        );

    \I__2364\ : Odrv12
    port map (
            O => \N__21387\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__2362\ : InMux
    port map (
            O => \N__21381\,
            I => \N__21377\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21380\,
            I => \N__21373\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__21377\,
            I => \N__21370\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21367\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21373\,
            I => \N__21361\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__21370\,
            I => \N__21361\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__21367\,
            I => \N__21358\
        );

    \I__2355\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21355\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__21361\,
            I => \N__21350\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__21358\,
            I => \N__21350\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__21355\,
            I => \N__21347\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__21350\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__21347\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_9\
        );

    \I__2349\ : InMux
    port map (
            O => \N__21342\,
            I => \bfn_3_18_0_\
        );

    \I__2348\ : InMux
    port map (
            O => \N__21339\,
            I => \N__21336\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__21336\,
            I => \N__21333\
        );

    \I__2346\ : Odrv12
    port map (
            O => \N__21333\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__21330\,
            I => \N__21326\
        );

    \I__2344\ : InMux
    port map (
            O => \N__21329\,
            I => \N__21321\
        );

    \I__2343\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21321\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__21321\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\
        );

    \I__2341\ : InMux
    port map (
            O => \N__21318\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__21315\,
            I => \N__21312\
        );

    \I__2339\ : InMux
    port map (
            O => \N__21312\,
            I => \N__21308\
        );

    \I__2338\ : InMux
    port map (
            O => \N__21311\,
            I => \N__21303\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21300\
        );

    \I__2336\ : InMux
    port map (
            O => \N__21307\,
            I => \N__21297\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21306\,
            I => \N__21294\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21289\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__21300\,
            I => \N__21289\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21286\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__21294\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__21289\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__21286\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_11\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21279\,
            I => \N__21273\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21273\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__21273\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\
        );

    \I__2325\ : InMux
    port map (
            O => \N__21270\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\
        );

    \I__2324\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21264\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__21264\,
            I => \N__21261\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__21261\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__21258\,
            I => \N__21254\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21250\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21246\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21243\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__21250\,
            I => \N__21240\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__21249\,
            I => \N__21237\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__21246\,
            I => \N__21234\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__21243\,
            I => \N__21231\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__21240\,
            I => \N__21228\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21237\,
            I => \N__21225\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__21234\,
            I => \N__21222\
        );

    \I__2310\ : Span4Mux_s2_h
    port map (
            O => \N__21231\,
            I => \N__21219\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__21228\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21225\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__21222\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__21219\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_12\
        );

    \I__2305\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21206\
        );

    \I__2304\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21203\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__21206\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__21203\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\
        );

    \I__2301\ : InMux
    port map (
            O => \N__21198\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\
        );

    \I__2300\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21189\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21189\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__21189\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\
        );

    \I__2297\ : InMux
    port map (
            O => \N__21186\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__21183\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\
        );

    \I__2295\ : InMux
    port map (
            O => \N__21180\,
            I => \N__21177\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__21177\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__21171\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__21168\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21162\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__21156\,
            I => \N__21152\
        );

    \I__2286\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21149\
        );

    \I__2285\ : Span4Mux_h
    port map (
            O => \N__21152\,
            I => \N__21146\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__21149\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2283\ : Odrv4
    port map (
            O => \N__21146\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\
        );

    \I__2282\ : CascadeMux
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21138\,
            I => \N__21133\
        );

    \I__2280\ : InMux
    port map (
            O => \N__21137\,
            I => \N__21130\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21136\,
            I => \N__21127\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21133\,
            I => \N__21124\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__21130\,
            I => \N__21120\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__21127\,
            I => \N__21117\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__21124\,
            I => \N__21114\
        );

    \I__2274\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21110\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__21120\,
            I => \N__21107\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__21117\,
            I => \N__21104\
        );

    \I__2271\ : Span4Mux_s3_h
    port map (
            O => \N__21114\,
            I => \N__21101\
        );

    \I__2270\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21098\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__21110\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__21107\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__21104\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__21101\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__21098\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_1\
        );

    \I__2264\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21084\,
            I => \N__21081\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__21081\,
            I => \N__21078\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__21078\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__21075\,
            I => \N__21071\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__21074\,
            I => \N__21068\
        );

    \I__2258\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21064\
        );

    \I__2257\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21061\
        );

    \I__2256\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21058\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21064\,
            I => \N__21053\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__21061\,
            I => \N__21053\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__21058\,
            I => \N__21050\
        );

    \I__2252\ : Span4Mux_v
    port map (
            O => \N__21053\,
            I => \N__21047\
        );

    \I__2251\ : Span4Mux_s2_h
    port map (
            O => \N__21050\,
            I => \N__21044\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__21047\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__21044\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_2\
        );

    \I__2248\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21036\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__21036\,
            I => \N__21033\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__21033\,
            I => \N__21030\
        );

    \I__2245\ : Span4Mux_v
    port map (
            O => \N__21030\,
            I => \N__21027\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__21027\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\
        );

    \I__2243\ : InMux
    port map (
            O => \N__21024\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\
        );

    \I__2242\ : InMux
    port map (
            O => \N__21021\,
            I => \N__21018\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__21018\,
            I => \N__21013\
        );

    \I__2240\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21007\
        );

    \I__2239\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21007\
        );

    \I__2238\ : Span4Mux_v
    port map (
            O => \N__21013\,
            I => \N__21004\
        );

    \I__2237\ : InMux
    port map (
            O => \N__21012\,
            I => \N__21001\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__21007\,
            I => \N__20998\
        );

    \I__2235\ : Odrv4
    port map (
            O => \N__21004\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__21001\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2233\ : Odrv12
    port map (
            O => \N__20998\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_3\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__20991\,
            I => \N__20988\
        );

    \I__2231\ : InMux
    port map (
            O => \N__20988\,
            I => \N__20985\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__20985\,
            I => \N__20982\
        );

    \I__2229\ : Odrv12
    port map (
            O => \N__20982\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\
        );

    \I__2228\ : InMux
    port map (
            O => \N__20979\,
            I => \N__20976\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__20976\,
            I => \N__20971\
        );

    \I__2226\ : InMux
    port map (
            O => \N__20975\,
            I => \N__20968\
        );

    \I__2225\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20965\
        );

    \I__2224\ : Span4Mux_s3_h
    port map (
            O => \N__20971\,
            I => \N__20962\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__20968\,
            I => \N__20957\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__20965\,
            I => \N__20957\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__20962\,
            I => \N__20954\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__20957\,
            I => \N__20951\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__20954\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2218\ : Odrv4
    port map (
            O => \N__20951\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto3\
        );

    \I__2217\ : InMux
    port map (
            O => \N__20946\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\
        );

    \I__2216\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20940\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__20940\,
            I => \N__20937\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__20937\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__20934\,
            I => \N__20931\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20925\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__20930\,
            I => \N__20922\
        );

    \I__2210\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20917\
        );

    \I__2209\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20917\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__20925\,
            I => \N__20914\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20922\,
            I => \N__20911\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__20917\,
            I => \N__20908\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__20914\,
            I => \N__20905\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__20911\,
            I => \N__20902\
        );

    \I__2203\ : Odrv4
    port map (
            O => \N__20908\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__20905\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2201\ : Odrv4
    port map (
            O => \N__20902\,
            I => \current_shift_inst.PI_CTRL.integratorZ0Z_4\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20891\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__20894\,
            I => \N__20886\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20883\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20890\,
            I => \N__20880\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20889\,
            I => \N__20875\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20875\
        );

    \I__2194\ : Span4Mux_s3_h
    port map (
            O => \N__20883\,
            I => \N__20872\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20867\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__20875\,
            I => \N__20867\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__20872\,
            I => \N__20864\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__20867\,
            I => \N__20861\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__20864\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__20861\,
            I => \current_shift_inst.PI_CTRL.un7_enablelto4\
        );

    \I__2187\ : InMux
    port map (
            O => \N__20856\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20850\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20847\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__20847\,
            I => \N__20844\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__20844\,
            I => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20841\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20838\,
            I => \N__20835\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20835\,
            I => \N__20832\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__20832\,
            I => \N__20829\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__20829\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__20826\,
            I => \N__20823\
        );

    \I__2176\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20820\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20820\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__20817\,
            I => \N__20814\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20814\,
            I => \N__20811\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__20811\,
            I => \N__20808\
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__20808\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__20805\,
            I => \N__20802\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20799\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__20796\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\
        );

    \I__2166\ : InMux
    port map (
            O => \N__20793\,
            I => \N__20790\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20790\,
            I => \N__20787\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__20787\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\
        );

    \I__2163\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20781\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20781\,
            I => \N__20778\
        );

    \I__2161\ : Span4Mux_h
    port map (
            O => \N__20778\,
            I => \N__20775\
        );

    \I__2160\ : Odrv4
    port map (
            O => \N__20775\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\
        );

    \I__2159\ : InMux
    port map (
            O => \N__20772\,
            I => \pwm_generator_inst.un15_threshold_1_cry_13\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20769\,
            I => \pwm_generator_inst.un15_threshold_1_cry_14\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20766\,
            I => \bfn_2_26_0_\
        );

    \I__2156\ : InMux
    port map (
            O => \N__20763\,
            I => \pwm_generator_inst.un15_threshold_1_cry_16\
        );

    \I__2155\ : InMux
    port map (
            O => \N__20760\,
            I => \pwm_generator_inst.un15_threshold_1_cry_17\
        );

    \I__2154\ : InMux
    port map (
            O => \N__20757\,
            I => \pwm_generator_inst.un15_threshold_1_cry_18\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20751\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__20751\,
            I => \N__20748\
        );

    \I__2151\ : Odrv4
    port map (
            O => \N__20748\,
            I => \N_88_i_i\
        );

    \I__2150\ : InMux
    port map (
            O => \N__20745\,
            I => \N__20742\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__20742\,
            I => \N__20739\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__20739\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\
        );

    \I__2147\ : InMux
    port map (
            O => \N__20736\,
            I => \N__20733\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__20733\,
            I => \N__20730\
        );

    \I__2145\ : Span4Mux_v
    port map (
            O => \N__20730\,
            I => \N__20727\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__20727\,
            I => \pwm_generator_inst.O_5\
        );

    \I__2143\ : InMux
    port map (
            O => \N__20724\,
            I => \N__20721\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__20721\,
            I => \pwm_generator_inst.un15_threshold_1_axb_5\
        );

    \I__2141\ : InMux
    port map (
            O => \N__20718\,
            I => \N__20715\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__20715\,
            I => \N__20712\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__20712\,
            I => \N__20709\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__20709\,
            I => \pwm_generator_inst.O_6\
        );

    \I__2137\ : InMux
    port map (
            O => \N__20706\,
            I => \N__20703\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__20703\,
            I => \pwm_generator_inst.un15_threshold_1_axb_6\
        );

    \I__2135\ : InMux
    port map (
            O => \N__20700\,
            I => \N__20697\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__20697\,
            I => \N__20694\
        );

    \I__2133\ : Span4Mux_h
    port map (
            O => \N__20694\,
            I => \N__20691\
        );

    \I__2132\ : Odrv4
    port map (
            O => \N__20691\,
            I => \pwm_generator_inst.O_7\
        );

    \I__2131\ : InMux
    port map (
            O => \N__20688\,
            I => \N__20685\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20685\,
            I => \pwm_generator_inst.un15_threshold_1_axb_7\
        );

    \I__2129\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__20679\,
            I => \N__20676\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__20676\,
            I => \N__20673\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__20673\,
            I => \pwm_generator_inst.O_8\
        );

    \I__2125\ : InMux
    port map (
            O => \N__20670\,
            I => \N__20667\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__20667\,
            I => \pwm_generator_inst.un15_threshold_1_axb_8\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20661\,
            I => \N__20658\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__20658\,
            I => \N__20655\
        );

    \I__2120\ : Odrv4
    port map (
            O => \N__20655\,
            I => \pwm_generator_inst.O_9\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20649\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20649\,
            I => \pwm_generator_inst.un15_threshold_1_axb_9\
        );

    \I__2117\ : InMux
    port map (
            O => \N__20646\,
            I => \pwm_generator_inst.un15_threshold_1_cry_9\
        );

    \I__2116\ : InMux
    port map (
            O => \N__20643\,
            I => \pwm_generator_inst.un15_threshold_1_cry_10\
        );

    \I__2115\ : InMux
    port map (
            O => \N__20640\,
            I => \pwm_generator_inst.un15_threshold_1_cry_11\
        );

    \I__2114\ : InMux
    port map (
            O => \N__20637\,
            I => \pwm_generator_inst.un15_threshold_1_cry_12\
        );

    \I__2113\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20629\
        );

    \I__2112\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20626\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20623\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__20629\,
            I => \N__20620\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__20626\,
            I => pwm_duty_input_9
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20623\,
            I => pwm_duty_input_9
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__20620\,
            I => pwm_duty_input_9
        );

    \I__2106\ : InMux
    port map (
            O => \N__20613\,
            I => \N__20609\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20612\,
            I => \N__20605\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20609\,
            I => \N__20602\
        );

    \I__2103\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20599\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__20605\,
            I => \N__20594\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__20602\,
            I => \N__20594\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20599\,
            I => pwm_duty_input_6
        );

    \I__2099\ : Odrv4
    port map (
            O => \N__20594\,
            I => pwm_duty_input_6
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__20589\,
            I => \N__20585\
        );

    \I__2097\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20581\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20585\,
            I => \N__20578\
        );

    \I__2095\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20575\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20572\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__20578\,
            I => pwm_duty_input_7
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__20575\,
            I => pwm_duty_input_7
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__20572\,
            I => pwm_duty_input_7
        );

    \I__2090\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20562\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__20562\,
            I => \N__20557\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20552\
        );

    \I__2087\ : InMux
    port map (
            O => \N__20560\,
            I => \N__20552\
        );

    \I__2086\ : Span4Mux_s1_h
    port map (
            O => \N__20557\,
            I => \N__20549\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__20552\,
            I => pwm_duty_input_8
        );

    \I__2084\ : Odrv4
    port map (
            O => \N__20549\,
            I => pwm_duty_input_8
        );

    \I__2083\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20539\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20543\,
            I => \N__20534\
        );

    \I__2081\ : InMux
    port map (
            O => \N__20542\,
            I => \N__20534\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__20539\,
            I => \N__20531\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20534\,
            I => pwm_duty_input_3
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__20531\,
            I => pwm_duty_input_3
        );

    \I__2077\ : InMux
    port map (
            O => \N__20526\,
            I => \N__20521\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20525\,
            I => \N__20516\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20524\,
            I => \N__20516\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__20521\,
            I => \N__20513\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20516\,
            I => pwm_duty_input_4
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__20513\,
            I => pwm_duty_input_4
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__20508\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__20505\,
            I => \N__20501\
        );

    \I__2069\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20498\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20501\,
            I => \N__20494\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20491\
        );

    \I__2066\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20488\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__20494\,
            I => \N__20483\
        );

    \I__2064\ : Span4Mux_v
    port map (
            O => \N__20491\,
            I => \N__20483\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__20488\,
            I => pwm_duty_input_5
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__20483\,
            I => pwm_duty_input_5
        );

    \I__2061\ : InMux
    port map (
            O => \N__20478\,
            I => \N__20475\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__20475\,
            I => \N__20472\
        );

    \I__2059\ : Span4Mux_h
    port map (
            O => \N__20472\,
            I => \N__20469\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__20469\,
            I => \pwm_generator_inst.O_0\
        );

    \I__2057\ : InMux
    port map (
            O => \N__20466\,
            I => \N__20463\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20463\,
            I => \pwm_generator_inst.un15_threshold_1_axb_0\
        );

    \I__2055\ : InMux
    port map (
            O => \N__20460\,
            I => \N__20457\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__20457\,
            I => \N__20454\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__20454\,
            I => \N__20451\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__20451\,
            I => \pwm_generator_inst.O_1\
        );

    \I__2051\ : InMux
    port map (
            O => \N__20448\,
            I => \N__20445\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__20445\,
            I => \pwm_generator_inst.un15_threshold_1_axb_1\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20442\,
            I => \N__20439\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__20436\,
            I => \N__20433\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__20433\,
            I => \pwm_generator_inst.O_2\
        );

    \I__2045\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__20427\,
            I => \pwm_generator_inst.un15_threshold_1_axb_2\
        );

    \I__2043\ : InMux
    port map (
            O => \N__20424\,
            I => \N__20421\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__20421\,
            I => \N__20418\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__20418\,
            I => \N__20415\
        );

    \I__2040\ : Odrv4
    port map (
            O => \N__20415\,
            I => \pwm_generator_inst.O_3\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20412\,
            I => \N__20409\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__20409\,
            I => \pwm_generator_inst.un15_threshold_1_axb_3\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20403\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20403\,
            I => \N__20400\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__20400\,
            I => \N__20397\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__20397\,
            I => \pwm_generator_inst.O_4\
        );

    \I__2033\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20391\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__20391\,
            I => \pwm_generator_inst.un15_threshold_1_axb_4\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__20388\,
            I => \current_shift_inst.PI_CTRL.N_31_cascade_\
        );

    \I__2030\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20382\,
            I => \current_shift_inst.PI_CTRL.N_91\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__20379\,
            I => \current_shift_inst.PI_CTRL.N_98_cascade_\
        );

    \I__2027\ : InMux
    port map (
            O => \N__20376\,
            I => \N__20357\
        );

    \I__2026\ : InMux
    port map (
            O => \N__20375\,
            I => \N__20357\
        );

    \I__2025\ : InMux
    port map (
            O => \N__20374\,
            I => \N__20357\
        );

    \I__2024\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20357\
        );

    \I__2023\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20357\
        );

    \I__2022\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20357\
        );

    \I__2021\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20354\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__20357\,
            I => \N__20351\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__20354\,
            I => \N__20348\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__20351\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__20348\,
            I => \current_shift_inst.PI_CTRL.N_158\
        );

    \I__2016\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20340\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__20340\,
            I => \current_shift_inst.PI_CTRL.N_96\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__20337\,
            I => \current_shift_inst.PI_CTRL.N_96_cascade_\
        );

    \I__2013\ : InMux
    port map (
            O => \N__20334\,
            I => \N__20325\
        );

    \I__2012\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20325\
        );

    \I__2011\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20325\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__20325\,
            I => \current_shift_inst.PI_CTRL.N_160\
        );

    \I__2009\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20318\
        );

    \I__2008\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20315\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__20318\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__20315\,
            I => \current_shift_inst.PI_CTRL.N_94\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20304\
        );

    \I__2004\ : InMux
    port map (
            O => \N__20309\,
            I => \N__20304\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__20304\,
            I => \current_shift_inst.PI_CTRL.N_31\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__20301\,
            I => \N__20296\
        );

    \I__2001\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20289\
        );

    \I__2000\ : InMux
    port map (
            O => \N__20299\,
            I => \N__20289\
        );

    \I__1999\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20282\
        );

    \I__1998\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20282\
        );

    \I__1997\ : InMux
    port map (
            O => \N__20294\,
            I => \N__20282\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20275\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__20282\,
            I => \N__20275\
        );

    \I__1994\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20269\
        );

    \I__1993\ : InMux
    port map (
            O => \N__20280\,
            I => \N__20269\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__20275\,
            I => \N__20266\
        );

    \I__1991\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20263\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__20269\,
            I => \N__20260\
        );

    \I__1989\ : Odrv4
    port map (
            O => \N__20266\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__20263\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__20260\,
            I => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\
        );

    \I__1986\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20250\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__20250\,
            I => \current_shift_inst.PI_CTRL.N_97\
        );

    \I__1984\ : InMux
    port map (
            O => \N__20247\,
            I => \N__20243\
        );

    \I__1983\ : InMux
    port map (
            O => \N__20246\,
            I => \N__20240\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20237\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__20240\,
            I => pwm_duty_input_1
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__20237\,
            I => pwm_duty_input_1
        );

    \I__1979\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20228\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__20231\,
            I => \N__20225\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__20228\,
            I => \N__20222\
        );

    \I__1976\ : InMux
    port map (
            O => \N__20225\,
            I => \N__20219\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__20222\,
            I => \N__20216\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__20219\,
            I => pwm_duty_input_2
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__20216\,
            I => pwm_duty_input_2
        );

    \I__1972\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20207\
        );

    \I__1971\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20204\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__20207\,
            I => \N__20201\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__20204\,
            I => pwm_duty_input_0
        );

    \I__1968\ : Odrv4
    port map (
            O => \N__20201\,
            I => pwm_duty_input_0
        );

    \I__1967\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20193\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__20193\,
            I => \pwm_generator_inst.un2_duty_input_0_o3_1Z0Z_0\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__20190\,
            I => \pwm_generator_inst.N_7_cascade_\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\
        );

    \I__1963\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20181\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__20181\,
            I => \N__20178\
        );

    \I__1961\ : Odrv4
    port map (
            O => \N__20178\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\
        );

    \I__1960\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20172\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__20172\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\
        );

    \I__1958\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20166\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20166\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__20163\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\
        );

    \I__1955\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20157\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__20157\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\
        );

    \I__1953\ : InMux
    port map (
            O => \N__20154\,
            I => \N__20151\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__20151\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\
        );

    \I__1951\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20145\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__20145\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__20142\,
            I => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__20139\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\
        );

    \I__1947\ : InMux
    port map (
            O => \N__20136\,
            I => \N__20133\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__20133\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\
        );

    \I__1945\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20127\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__20127\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\
        );

    \I__1943\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20121\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__20121\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\
        );

    \I__1941\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20115\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__20115\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__20112\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20106\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__20106\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20100\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__20100\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__20097\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\
        );

    \I__1933\ : InMux
    port map (
            O => \N__20094\,
            I => \N__20091\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20091\,
            I => \current_shift_inst.PI_CTRL.N_44\
        );

    \I__1931\ : InMux
    port map (
            O => \N__20088\,
            I => \N__20085\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__20085\,
            I => \current_shift_inst.PI_CTRL.N_77\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__20082\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\
        );

    \I__1928\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20076\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__20076\,
            I => \N__20073\
        );

    \I__1926\ : Odrv4
    port map (
            O => \N__20073\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\
        );

    \I__1925\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20067\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__20067\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__20064\,
            I => \current_shift_inst.PI_CTRL.N_43_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20058\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__20058\,
            I => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__20055\,
            I => \N__20052\
        );

    \I__1919\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20049\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__20049\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__20046\,
            I => \N__20043\
        );

    \I__1916\ : InMux
    port map (
            O => \N__20043\,
            I => \N__20040\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__20040\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\
        );

    \I__1914\ : InMux
    port map (
            O => \N__20037\,
            I => \N__20034\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__20034\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20028\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__20028\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__1909\ : InMux
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20019\,
            I => \N__20016\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__20016\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\
        );

    \I__1906\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20010\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20004\,
            I => \N__20001\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__20001\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\
        );

    \I__1901\ : InMux
    port map (
            O => \N__19998\,
            I => \N__19995\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__19995\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\
        );

    \I__1899\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19989\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__19989\,
            I => un7_start_stop
        );

    \I__1897\ : InMux
    port map (
            O => \N__19986\,
            I => \N__19983\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__19983\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__19980\,
            I => \N__19976\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__19979\,
            I => \N__19973\
        );

    \I__1893\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19970\
        );

    \I__1892\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19967\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__19970\,
            I => \N__19962\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__19967\,
            I => \N__19962\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__19962\,
            I => \N__19959\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__19959\,
            I => \N__19956\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__19956\,
            I => \current_shift_inst.PI_CTRL.un1_integrator\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19950\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__19950\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\
        );

    \I__1884\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19944\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__19944\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\
        );

    \I__1882\ : InMux
    port map (
            O => \N__19941\,
            I => \N__19938\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19938\,
            I => \N__19935\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__19935\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\
        );

    \I__1879\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19929\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__19929\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\
        );

    \I__1877\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19923\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__19923\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\
        );

    \I__1875\ : InMux
    port map (
            O => \N__19920\,
            I => \N__19917\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19917\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\
        );

    \I__1873\ : InMux
    port map (
            O => \N__19914\,
            I => \N__19911\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__19911\,
            I => \N__19908\
        );

    \I__1871\ : Odrv12
    port map (
            O => \N__19908\,
            I => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__19905\,
            I => \N__19902\
        );

    \I__1869\ : InMux
    port map (
            O => \N__19902\,
            I => \N__19899\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__19899\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\
        );

    \I__1867\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19893\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__19893\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__19890\,
            I => \N__19887\
        );

    \I__1864\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19884\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__19884\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__19881\,
            I => \N__19878\
        );

    \I__1861\ : InMux
    port map (
            O => \N__19878\,
            I => \N__19875\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__19875\,
            I => \N__19872\
        );

    \I__1859\ : Odrv12
    port map (
            O => \N__19872\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\
        );

    \I__1858\ : InMux
    port map (
            O => \N__19869\,
            I => \N__19866\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__19866\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__19863\,
            I => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__1854\ : InMux
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19851\
        );

    \I__1852\ : Odrv12
    port map (
            O => \N__19851\,
            I => \current_shift_inst.PI_CTRL.integrator_1_26\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19848\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__19845\,
            I => \N__19842\
        );

    \I__1849\ : InMux
    port map (
            O => \N__19842\,
            I => \N__19839\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__19839\,
            I => \N__19836\
        );

    \I__1847\ : Span4Mux_v
    port map (
            O => \N__19836\,
            I => \N__19833\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__19833\,
            I => \current_shift_inst.PI_CTRL.integrator_1_27\
        );

    \I__1845\ : InMux
    port map (
            O => \N__19830\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__19827\,
            I => \N__19824\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19821\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__19821\,
            I => \N__19818\
        );

    \I__1841\ : Span4Mux_v
    port map (
            O => \N__19818\,
            I => \N__19815\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__19815\,
            I => \current_shift_inst.PI_CTRL.integrator_1_28\
        );

    \I__1839\ : InMux
    port map (
            O => \N__19812\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__19809\,
            I => \N__19806\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19803\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19803\,
            I => \N__19800\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__19800\,
            I => \N__19797\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__19797\,
            I => \current_shift_inst.PI_CTRL.integrator_1_29\
        );

    \I__1833\ : InMux
    port map (
            O => \N__19794\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__19791\,
            I => \N__19788\
        );

    \I__1831\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19785\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__19785\,
            I => \N__19782\
        );

    \I__1829\ : Span4Mux_v
    port map (
            O => \N__19782\,
            I => \N__19779\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__19779\,
            I => \current_shift_inst.PI_CTRL.integrator_1_30\
        );

    \I__1827\ : InMux
    port map (
            O => \N__19776\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\
        );

    \I__1826\ : InMux
    port map (
            O => \N__19773\,
            I => \N__19770\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__19770\,
            I => \N__19767\
        );

    \I__1824\ : Odrv12
    port map (
            O => \N__19767\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__19764\,
            I => \N__19761\
        );

    \I__1822\ : InMux
    port map (
            O => \N__19761\,
            I => \N__19758\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__19758\,
            I => \N__19755\
        );

    \I__1820\ : Odrv12
    port map (
            O => \N__19755\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\
        );

    \I__1819\ : InMux
    port map (
            O => \N__19752\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\
        );

    \I__1818\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19746\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__19746\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__19743\,
            I => \N__19740\
        );

    \I__1815\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__19737\,
            I => \N__19734\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__19734\,
            I => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\
        );

    \I__1812\ : InMux
    port map (
            O => \N__19731\,
            I => \bfn_1_14_0_\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__19728\,
            I => \N__19725\
        );

    \I__1810\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19722\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__19722\,
            I => \N__19719\
        );

    \I__1808\ : Span4Mux_v
    port map (
            O => \N__19719\,
            I => \N__19716\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__19716\,
            I => \current_shift_inst.PI_CTRL.integrator_1_18\
        );

    \I__1806\ : InMux
    port map (
            O => \N__19713\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__19710\,
            I => \N__19707\
        );

    \I__1804\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19704\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__19704\,
            I => \N__19701\
        );

    \I__1802\ : Span4Mux_v
    port map (
            O => \N__19701\,
            I => \N__19698\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__19698\,
            I => \current_shift_inst.PI_CTRL.integrator_1_19\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19695\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19689\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__19689\,
            I => \N__19686\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__19686\,
            I => \N__19683\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__19683\,
            I => \current_shift_inst.PI_CTRL.integrator_1_20\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19680\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__19677\,
            I => \N__19674\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19674\,
            I => \N__19671\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__19671\,
            I => \N__19668\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__19668\,
            I => \N__19665\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__19665\,
            I => \current_shift_inst.PI_CTRL.integrator_1_21\
        );

    \I__1789\ : InMux
    port map (
            O => \N__19662\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__19659\,
            I => \N__19656\
        );

    \I__1787\ : InMux
    port map (
            O => \N__19656\,
            I => \N__19653\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19653\,
            I => \N__19650\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__19650\,
            I => \N__19647\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__19647\,
            I => \current_shift_inst.PI_CTRL.integrator_1_22\
        );

    \I__1783\ : InMux
    port map (
            O => \N__19644\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\
        );

    \I__1782\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19638\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__19638\,
            I => \N__19635\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__19635\,
            I => \current_shift_inst.PI_CTRL.integrator_1_23\
        );

    \I__1779\ : InMux
    port map (
            O => \N__19632\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__19629\,
            I => \N__19626\
        );

    \I__1777\ : InMux
    port map (
            O => \N__19626\,
            I => \N__19623\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__19623\,
            I => \N__19620\
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__19620\,
            I => \current_shift_inst.PI_CTRL.integrator_1_24\
        );

    \I__1774\ : InMux
    port map (
            O => \N__19617\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\
        );

    \I__1773\ : InMux
    port map (
            O => \N__19614\,
            I => \N__19611\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__19611\,
            I => \N__19608\
        );

    \I__1771\ : Span4Mux_v
    port map (
            O => \N__19608\,
            I => \N__19605\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__19605\,
            I => \current_shift_inst.PI_CTRL.integrator_1_25\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19602\,
            I => \bfn_1_15_0_\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__19599\,
            I => \N__19596\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19593\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__1765\ : Span4Mux_v
    port map (
            O => \N__19590\,
            I => \N__19587\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__19587\,
            I => \N__19584\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__19584\,
            I => \current_shift_inst.PI_CTRL.integrator_1_9\
        );

    \I__1762\ : InMux
    port map (
            O => \N__19581\,
            I => \bfn_1_13_0_\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__19578\,
            I => \N__19575\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19572\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19572\,
            I => \N__19569\
        );

    \I__1758\ : Span4Mux_v
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__1757\ : Span4Mux_v
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__19563\,
            I => \current_shift_inst.PI_CTRL.integrator_1_10\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19560\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__19545\,
            I => \current_shift_inst.PI_CTRL.integrator_1_11\
        );

    \I__1749\ : InMux
    port map (
            O => \N__19542\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__19539\,
            I => \N__19536\
        );

    \I__1747\ : InMux
    port map (
            O => \N__19536\,
            I => \N__19533\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19530\
        );

    \I__1745\ : Span4Mux_v
    port map (
            O => \N__19530\,
            I => \N__19527\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__19527\,
            I => \current_shift_inst.PI_CTRL.integrator_1_12\
        );

    \I__1743\ : InMux
    port map (
            O => \N__19524\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__19521\,
            I => \N__19518\
        );

    \I__1741\ : InMux
    port map (
            O => \N__19518\,
            I => \N__19515\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__19515\,
            I => \N__19512\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__19512\,
            I => \N__19509\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__19509\,
            I => \current_shift_inst.PI_CTRL.integrator_1_13\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19506\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \N__19500\
        );

    \I__1735\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19497\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19494\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__19494\,
            I => \N__19491\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__19491\,
            I => \current_shift_inst.PI_CTRL.integrator_1_14\
        );

    \I__1731\ : InMux
    port map (
            O => \N__19488\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__19485\,
            I => \N__19482\
        );

    \I__1729\ : InMux
    port map (
            O => \N__19482\,
            I => \N__19479\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19479\,
            I => \N__19476\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__19476\,
            I => \N__19473\
        );

    \I__1726\ : Odrv4
    port map (
            O => \N__19473\,
            I => \current_shift_inst.PI_CTRL.integrator_1_15\
        );

    \I__1725\ : InMux
    port map (
            O => \N__19470\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19464\,
            I => \N__19461\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19458\
        );

    \I__1721\ : Odrv12
    port map (
            O => \N__19458\,
            I => \current_shift_inst.PI_CTRL.integrator_1_16\
        );

    \I__1720\ : InMux
    port map (
            O => \N__19455\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__19452\,
            I => \N__19449\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19446\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__19446\,
            I => \N__19443\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__19443\,
            I => \N__19440\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__19440\,
            I => \current_shift_inst.PI_CTRL.integrator_1_17\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__19437\,
            I => \N__19434\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19431\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__19431\,
            I => \N__19428\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__19428\,
            I => \N__19425\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__19422\,
            I => \current_shift_inst.PI_CTRL.integrator_1_2\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19419\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__19416\,
            I => \N__19413\
        );

    \I__1706\ : InMux
    port map (
            O => \N__19413\,
            I => \N__19410\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__19410\,
            I => \N__19407\
        );

    \I__1704\ : Span4Mux_v
    port map (
            O => \N__19407\,
            I => \N__19404\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__19404\,
            I => \current_shift_inst.PI_CTRL.integrator_1_3\
        );

    \I__1702\ : InMux
    port map (
            O => \N__19401\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\
        );

    \I__1701\ : InMux
    port map (
            O => \N__19398\,
            I => \N__19395\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__19395\,
            I => \N__19392\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__19392\,
            I => \N__19389\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__19389\,
            I => \current_shift_inst.PI_CTRL.integrator_1_4\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19386\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19383\,
            I => \N__19380\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__19380\,
            I => \N__19377\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__19377\,
            I => \N__19374\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__19374\,
            I => \current_shift_inst.PI_CTRL.integrator_1_5\
        );

    \I__1692\ : InMux
    port map (
            O => \N__19371\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\
        );

    \I__1691\ : CascadeMux
    port map (
            O => \N__19368\,
            I => \N__19365\
        );

    \I__1690\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19362\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__19362\,
            I => \N__19359\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__19359\,
            I => \N__19356\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__19356\,
            I => \current_shift_inst.PI_CTRL.integrator_1_6\
        );

    \I__1686\ : InMux
    port map (
            O => \N__19353\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__19350\,
            I => \N__19347\
        );

    \I__1684\ : InMux
    port map (
            O => \N__19347\,
            I => \N__19344\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__19344\,
            I => \N__19341\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__19341\,
            I => \N__19338\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__19338\,
            I => \current_shift_inst.PI_CTRL.integrator_1_7\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19335\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__19332\,
            I => \N__19329\
        );

    \I__1678\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19326\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__19326\,
            I => \N__19323\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__19323\,
            I => \N__19320\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__19320\,
            I => \current_shift_inst.PI_CTRL.integrator_1_8\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19317\,
            I => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19311\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19311\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_8\
        );

    \I__1671\ : InMux
    port map (
            O => \N__19308\,
            I => \bfn_1_10_0_\
        );

    \I__1670\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__19302\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_9\
        );

    \I__1668\ : InMux
    port map (
            O => \N__19299\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19293\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19293\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_10\
        );

    \I__1665\ : InMux
    port map (
            O => \N__19290\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19284\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__19284\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_11\
        );

    \I__1662\ : InMux
    port map (
            O => \N__19281\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\
        );

    \I__1661\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__19275\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_12\
        );

    \I__1659\ : InMux
    port map (
            O => \N__19272\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\
        );

    \I__1658\ : InMux
    port map (
            O => \N__19269\,
            I => \N__19266\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__19266\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_13\
        );

    \I__1656\ : InMux
    port map (
            O => \N__19263\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19257\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__19257\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_14\
        );

    \I__1653\ : InMux
    port map (
            O => \N__19254\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\
        );

    \I__1652\ : InMux
    port map (
            O => \N__19251\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__19245\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_15\
        );

    \I__1649\ : InMux
    port map (
            O => \N__19242\,
            I => \N__19228\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__19241\,
            I => \N__19225\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__19240\,
            I => \N__19222\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__19239\,
            I => \N__19219\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__19238\,
            I => \N__19216\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__19237\,
            I => \N__19213\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__19236\,
            I => \N__19210\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__19235\,
            I => \N__19207\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__19234\,
            I => \N__19204\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__19233\,
            I => \N__19201\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__19232\,
            I => \N__19198\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__19231\,
            I => \N__19195\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__19228\,
            I => \N__19192\
        );

    \I__1636\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19185\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19222\,
            I => \N__19185\
        );

    \I__1634\ : InMux
    port map (
            O => \N__19219\,
            I => \N__19185\
        );

    \I__1633\ : InMux
    port map (
            O => \N__19216\,
            I => \N__19176\
        );

    \I__1632\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19176\
        );

    \I__1631\ : InMux
    port map (
            O => \N__19210\,
            I => \N__19176\
        );

    \I__1630\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19176\
        );

    \I__1629\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19171\
        );

    \I__1628\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19171\
        );

    \I__1627\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19166\
        );

    \I__1626\ : InMux
    port map (
            O => \N__19195\,
            I => \N__19166\
        );

    \I__1625\ : Span4Mux_v
    port map (
            O => \N__19192\,
            I => \N__19155\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19155\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__19176\,
            I => \N__19155\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__19171\,
            I => \N__19155\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__19166\,
            I => \N__19155\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__19155\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_19\
        );

    \I__1619\ : InMux
    port map (
            O => \N__19152\,
            I => \N__19149\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__19149\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_0\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__19146\,
            I => \N__19143\
        );

    \I__1616\ : InMux
    port map (
            O => \N__19143\,
            I => \N__19140\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19137\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__19137\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_15\
        );

    \I__1613\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19131\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__19131\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_1\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__19128\,
            I => \N__19125\
        );

    \I__1610\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19122\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__19122\,
            I => \N__19119\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__19119\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_16\
        );

    \I__1607\ : InMux
    port map (
            O => \N__19116\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\
        );

    \I__1606\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19110\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__19110\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_2\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__19107\,
            I => \N__19104\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19101\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__19101\,
            I => \N__19098\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__19098\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_17\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19095\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\
        );

    \I__1599\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19089\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__19089\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_3\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__19086\,
            I => \N__19083\
        );

    \I__1596\ : InMux
    port map (
            O => \N__19083\,
            I => \N__19080\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__19080\,
            I => \N__19077\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__19077\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_1_18\
        );

    \I__1593\ : InMux
    port map (
            O => \N__19074\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\
        );

    \I__1592\ : InMux
    port map (
            O => \N__19071\,
            I => \N__19068\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__19068\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_4\
        );

    \I__1590\ : InMux
    port map (
            O => \N__19065\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\
        );

    \I__1589\ : InMux
    port map (
            O => \N__19062\,
            I => \N__19059\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__19059\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_5\
        );

    \I__1587\ : InMux
    port map (
            O => \N__19056\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\
        );

    \I__1586\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19050\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__19050\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_6\
        );

    \I__1584\ : InMux
    port map (
            O => \N__19047\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\
        );

    \I__1583\ : InMux
    port map (
            O => \N__19044\,
            I => \N__19041\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__19041\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_2_7\
        );

    \I__1581\ : InMux
    port map (
            O => \N__19038\,
            I => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\
        );

    \I__1580\ : IoInMux
    port map (
            O => \N__19035\,
            I => \N__19032\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__19032\,
            I => \N__19029\
        );

    \I__1578\ : Span4Mux_s3_v
    port map (
            O => \N__19029\,
            I => \N__19026\
        );

    \I__1577\ : Span4Mux_h
    port map (
            O => \N__19026\,
            I => \N__19023\
        );

    \I__1576\ : Sp12to4
    port map (
            O => \N__19023\,
            I => \N__19020\
        );

    \I__1575\ : Span12Mux_v
    port map (
            O => \N__19020\,
            I => \N__19017\
        );

    \I__1574\ : Span12Mux_v
    port map (
            O => \N__19017\,
            I => \N__19014\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__19014\,
            I => delay_tr_input_ibuf_gb_io_gb_input
        );

    \I__1572\ : IoInMux
    port map (
            O => \N__19011\,
            I => \N__19008\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__19008\,
            I => \N__19005\
        );

    \I__1570\ : IoSpan4Mux
    port map (
            O => \N__19005\,
            I => \N__19002\
        );

    \I__1569\ : IoSpan4Mux
    port map (
            O => \N__19002\,
            I => \N__18999\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__18999\,
            I => delay_hc_input_ibuf_gb_io_gb_input
        );

    \IN_MUX_bfv_4_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_22_0_\
        );

    \IN_MUX_bfv_4_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_7\,
            carryinitout => \bfn_4_23_0_\
        );

    \IN_MUX_bfv_4_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un3_threshold_cry_15\,
            carryinitout => \bfn_4_24_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_17_8_0_\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s1\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s1\,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_13_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s1\,
            carryinitout => \bfn_13_19_0_\
        );

    \IN_MUX_bfv_14_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_13_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_7_s0\,
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_15_s0\,
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un38_control_input_cry_23_s0\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_15_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_21_0_\
        );

    \IN_MUX_bfv_15_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_7\,
            carryinitout => \bfn_15_22_0_\
        );

    \IN_MUX_bfv_15_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_15\,
            carryinitout => \bfn_15_23_0_\
        );

    \IN_MUX_bfv_15_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un10_control_input_cry_23\,
            carryinitout => \bfn_15_24_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_3_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_17_0_\
        );

    \IN_MUX_bfv_3_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            carryinitout => \bfn_3_18_0_\
        );

    \IN_MUX_bfv_3_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            carryinitout => \bfn_3_19_0_\
        );

    \IN_MUX_bfv_3_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            carryinitout => \bfn_3_20_0_\
        );

    \IN_MUX_bfv_5_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_23_0_\
        );

    \IN_MUX_bfv_5_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            carryinitout => \bfn_5_24_0_\
        );

    \IN_MUX_bfv_5_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            carryinitout => \bfn_5_25_0_\
        );

    \IN_MUX_bfv_3_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_24_0_\
        );

    \IN_MUX_bfv_3_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un19_threshold_cry_7\,
            carryinitout => \bfn_3_25_0_\
        );

    \IN_MUX_bfv_2_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_24_0_\
        );

    \IN_MUX_bfv_2_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_7\,
            carryinitout => \bfn_2_25_0_\
        );

    \IN_MUX_bfv_2_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un15_threshold_1_cry_15\,
            carryinitout => \bfn_2_26_0_\
        );

    \IN_MUX_bfv_8_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_24_0_\
        );

    \IN_MUX_bfv_8_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.un14_counter_cry_7\,
            carryinitout => \bfn_8_25_0_\
        );

    \IN_MUX_bfv_7_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_26_0_\
        );

    \IN_MUX_bfv_7_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \pwm_generator_inst.counter_cry_7\,
            carryinitout => \bfn_7_27_0_\
        );

    \IN_MUX_bfv_10_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_8_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_16_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_7_0_\
        );

    \IN_MUX_bfv_16_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_16_8_0_\
        );

    \IN_MUX_bfv_16_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_16_9_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_8_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_11_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_8_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_16_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_12_0_\
        );

    \IN_MUX_bfv_16_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_13_0_\
        );

    \IN_MUX_bfv_18_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_11_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_7\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_15\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.control_input_cry_23\,
            carryinitout => \bfn_11_16_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_16_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            carryinitout => \bfn_16_20_0_\
        );

    \IN_MUX_bfv_16_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            carryinitout => \bfn_16_21_0_\
        );

    \IN_MUX_bfv_16_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            carryinitout => \bfn_16_22_0_\
        );

    \IN_MUX_bfv_17_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_15_0_\
        );

    \IN_MUX_bfv_17_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_8\,
            carryinitout => \bfn_17_16_0_\
        );

    \IN_MUX_bfv_17_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_16\,
            carryinitout => \bfn_17_17_0_\
        );

    \IN_MUX_bfv_17_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.un4_control_input_1_cry_24\,
            carryinitout => \bfn_17_18_0_\
        );

    \IN_MUX_bfv_17_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_23_0_\
        );

    \IN_MUX_bfv_17_24_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_7\,
            carryinitout => \bfn_17_24_0_\
        );

    \IN_MUX_bfv_17_25_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_15\,
            carryinitout => \bfn_17_25_0_\
        );

    \IN_MUX_bfv_17_26_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.timer_s1.counter_cry_23\,
            carryinitout => \bfn_17_26_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_9_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            carryinitout => \bfn_9_16_0_\
        );

    \delay_tr_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19035\,
            GLOBALBUFFEROUTPUT => delay_tr_input_c_g
        );

    \delay_hc_input_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19011\,
            GLOBALBUFFEROUTPUT => delay_hc_input_c_g
        );

    \current_shift_inst.timer_s1.running_RNII51H_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34794\,
            GLOBALBUFFEROUTPUT => \current_shift_inst.timer_s1.N_161_i_g\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__33684\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_tr.un1_start_g\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__41286\,
            GLOBALBUFFEROUTPUT => \phase_controller_inst2.stoper_hc.un1_start_g\
        );

    \osc\ : SB_HFOSC
    generic map (
            CLKHF_DIV => "0b10"
        )
    port map (
            CLKHFPU => \N__38678\,
            CLKHFEN => \N__38680\,
            CLKHF => clk_12mhz
        );

    \rgb_drv\ : SB_RGBA_DRV
    generic map (
            RGB2_CURRENT => "0b111111",
            CURRENT_MODE => "0b0",
            RGB0_CURRENT => "0b111111",
            RGB1_CURRENT => "0b111111"
        )
    port map (
            RGBLEDEN => \N__38679\,
            RGB2PWM => \N__20754\,
            RGB1 => rgb_g_wire,
            CURREN => \N__38848\,
            RGB2 => rgb_b_wire,
            RGB1PWM => \N__19992\,
            RGB0PWM => \N__49479\,
            RGB0 => rgb_r_wire
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19152\,
            in2 => \N__19146\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_16\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_s_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19134\,
            in2 => \N__19128\,
            in3 => \N__19116\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_s_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19113\,
            in2 => \N__19107\,
            in3 => \N__19095\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_s_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19092\,
            in2 => \N__19086\,
            in3 => \N__19074\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_s_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19071\,
            in2 => \N__19231\,
            in3 => \N__19065\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_s_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19062\,
            in2 => \N__19233\,
            in3 => \N__19056\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_s_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19053\,
            in2 => \N__19232\,
            in3 => \N__19047\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_s_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19044\,
            in2 => \N__19234\,
            in3 => \N__19038\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_s_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19314\,
            in2 => \N__19235\,
            in3 => \N__19308\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_24\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_s_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19305\,
            in2 => \N__19239\,
            in3 => \N__19299\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_s_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19296\,
            in2 => \N__19236\,
            in3 => \N__19290\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_s_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19287\,
            in2 => \N__19240\,
            in3 => \N__19281\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_s_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19278\,
            in2 => \N__19237\,
            in3 => \N__19272\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_s_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19269\,
            in2 => \N__19241\,
            in3 => \N__19263\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_s_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19260\,
            in2 => \N__19238\,
            in3 => \N__19254\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19251\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19248\,
            in2 => \_gnd_net_\,
            in3 => \N__19242\,
            lcout => \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.un1_integrator_cry_1_c_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21113\,
            in2 => \N__19979\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_2_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21067\,
            in2 => \N__19437\,
            in3 => \N__19419\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_3_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21012\,
            in2 => \N__19416\,
            in3 => \N__19401\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19398\,
            in2 => \N__20930\,
            in3 => \N__19386\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19383\,
            in2 => \N__22670\,
            in3 => \N__19371\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21509\,
            in2 => \N__19368\,
            in3 => \N__19353\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21453\,
            in2 => \N__19350\,
            in3 => \N__19335\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21430\,
            in2 => \N__19332\,
            in3 => \N__19317\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21376\,
            in2 => \N__19599\,
            in3 => \N__19581\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22917\,
            in2 => \N__19578\,
            in3 => \N__19560\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21307\,
            in2 => \N__19557\,
            in3 => \N__19542\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21253\,
            in2 => \N__19539\,
            in3 => \N__19524\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22965\,
            in2 => \N__19521\,
            in3 => \N__19506\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21858\,
            in2 => \N__19503\,
            in3 => \N__19488\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23007\,
            in2 => \N__19485\,
            in3 => \N__19470\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22882\,
            in2 => \N__19467\,
            in3 => \N__19455\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21774\,
            in2 => \N__19452\,
            in3 => \N__19731\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21718\,
            in2 => \N__19728\,
            in3 => \N__19713\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21663\,
            in2 => \N__19710\,
            in3 => \N__19695\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19692\,
            in2 => \N__21619\,
            in3 => \N__19680\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21558\,
            in2 => \N__19677\,
            in3 => \N__19662\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22302\,
            in2 => \N__19659\,
            in3 => \N__19644\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19641\,
            in2 => \N__22247\,
            in3 => \N__19632\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22182\,
            in2 => \N__19629\,
            in3 => \N__19617\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19614\,
            in2 => \N__22136\,
            in3 => \N__19602\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22075\,
            in2 => \N__19860\,
            in3 => \N__19848\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22017\,
            in2 => \N__19845\,
            in3 => \N__19830\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21963\,
            in2 => \N__19827\,
            in3 => \N__19812\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21908\,
            in2 => \N__19809\,
            in3 => \N__19794\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22590\,
            in2 => \N__19791\,
            in3 => \N__19776\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.un1_integrator_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.un1_integrator_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNO_0_31_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__19773\,
            in1 => \N__23506\,
            in2 => \N__19764\,
            in3 => \N__19752\,
            lcout => \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_27_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23519\,
            in1 => \N__23203\,
            in2 => \N__23378\,
            in3 => \N__19749\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.integrator_29_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23201\,
            in1 => \N__23522\,
            in2 => \N__19743\,
            in3 => \N__23339\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.integrator_31_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23202\,
            in1 => \N__23523\,
            in2 => \N__19905\,
            in3 => \N__23340\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.integrator_30_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000100010"
        )
    port map (
            in0 => \N__23520\,
            in1 => \N__23204\,
            in2 => \N__23379\,
            in3 => \N__19896\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.integrator_26_LC_1_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010011100100"
        )
    port map (
            in0 => \N__23200\,
            in1 => \N__23521\,
            in2 => \N__19890\,
            in3 => \N__23338\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49901\,
            ce => 'H',
            sr => \N__49438\
        );

    \current_shift_inst.PI_CTRL.integrator_12_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23524\,
            in1 => \N__23369\,
            in2 => \N__19881\,
            in3 => \N__23230\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49888\,
            ce => 'H',
            sr => \N__49441\
        );

    \current_shift_inst.PI_CTRL.prop_term_1_LC_1_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28734\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => 'H',
            sr => \N__49444\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_LC_1_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21155\,
            in2 => \_gnd_net_\,
            in3 => \N__21137\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49878\,
            ce => 'H',
            sr => \N__49444\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIRN52_15_LC_1_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21807\,
            in2 => \_gnd_net_\,
            in3 => \N__21828\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI3EH5_22_LC_1_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22104\,
            in1 => \N__19869\,
            in2 => \N__22275\,
            in3 => \N__22050\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_11_LC_1_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20118\,
            in1 => \N__20148\,
            in2 => \N__19863\,
            in3 => \N__20103\,
            lcout => \current_shift_inst.PI_CTRL.N_158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_5_LC_1_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__29782\,
            in1 => \N__20371\,
            in2 => \N__22386\,
            in3 => \N__20299\,
            lcout => pwm_duty_input_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_6_LC_1_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000011111100"
        )
    port map (
            in0 => \N__20372\,
            in1 => \N__20294\,
            in2 => \N__22515\,
            in3 => \N__29783\,
            lcout => pwm_duty_input_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_7_LC_1_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111010000"
        )
    port map (
            in0 => \N__29784\,
            in1 => \N__20373\,
            in2 => \N__22422\,
            in3 => \N__20300\,
            lcout => pwm_duty_input_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_3_LC_1_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__20979\,
            in1 => \N__20343\,
            in2 => \_gnd_net_\,
            in3 => \N__20322\,
            lcout => pwm_duty_input_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_9_LC_1_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110101010000"
        )
    port map (
            in0 => \N__29786\,
            in1 => \N__20375\,
            in2 => \N__20301\,
            in3 => \N__22484\,
            lcout => pwm_duty_input_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_8_LC_1_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110110000"
        )
    port map (
            in0 => \N__20374\,
            in1 => \N__29785\,
            in2 => \N__22455\,
            in3 => \N__20295\,
            lcout => pwm_duty_input_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_4_LC_1_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__20376\,
            in1 => \N__20895\,
            in2 => \N__22347\,
            in3 => \N__20385\,
            lcout => pwm_duty_input_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49832\,
            ce => 'H',
            sr => \N__49453\
        );

    \current_shift_inst.PI_CTRL.control_out_2_LC_1_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21039\,
            in2 => \_gnd_net_\,
            in3 => \N__20334\,
            lcout => pwm_duty_input_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49825\,
            ce => 'H',
            sr => \N__49454\
        );

    \current_shift_inst.PI_CTRL.control_out_1_LC_1_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20333\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19914\,
            lcout => pwm_duty_input_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49825\,
            ce => 'H',
            sr => \N__49454\
        );

    \current_shift_inst.PI_CTRL.control_out_0_LC_1_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22527\,
            in2 => \_gnd_net_\,
            in3 => \N__20332\,
            lcout => pwm_duty_input_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49825\,
            ce => 'H',
            sr => \N__49454\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_inv_LC_1_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__23897\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23915\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.un7_start_stop_LC_1_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__49478\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35106\,
            lcout => un7_start_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_7_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001100000001"
        )
    port map (
            in0 => \N__23388\,
            in1 => \N__23578\,
            in2 => \N__23241\,
            in3 => \N__19986\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49418\
        );

    \current_shift_inst.PI_CTRL.integrator_1_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001001000"
        )
    port map (
            in0 => \N__21123\,
            in1 => \N__23390\,
            in2 => \N__19980\,
            in3 => \N__23213\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49418\
        );

    \current_shift_inst.PI_CTRL.integrator_3_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__19953\,
            in1 => \N__23389\,
            in2 => \_gnd_net_\,
            in3 => \N__23212\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49935\,
            ce => 'H',
            sr => \N__49418\
        );

    \current_shift_inst.PI_CTRL.integrator_19_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23387\,
            in1 => \N__23586\,
            in2 => \N__23243\,
            in3 => \N__19947\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49924\,
            ce => 'H',
            sr => \N__49422\
        );

    \current_shift_inst.PI_CTRL.integrator_4_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23423\,
            in1 => \N__23585\,
            in2 => \N__23239\,
            in3 => \N__19941\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_23_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__23581\,
            in1 => \N__23426\,
            in2 => \N__23245\,
            in3 => \N__19932\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_17_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23420\,
            in1 => \N__23582\,
            in2 => \N__23237\,
            in3 => \N__19926\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_20_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001010"
        )
    port map (
            in0 => \N__23580\,
            in1 => \N__23425\,
            in2 => \N__23244\,
            in3 => \N__19920\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_24_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101100"
        )
    port map (
            in0 => \N__23422\,
            in1 => \N__23584\,
            in2 => \N__20055\,
            in3 => \N__23223\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_14_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23579\,
            in1 => \N__23424\,
            in2 => \N__20046\,
            in3 => \N__23196\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_22_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23421\,
            in1 => \N__23583\,
            in2 => \N__23238\,
            in3 => \N__20037\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49912\,
            ce => 'H',
            sr => \N__49427\
        );

    \current_shift_inst.PI_CTRL.integrator_25_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100111111001000"
        )
    port map (
            in0 => \N__23371\,
            in1 => \N__20031\,
            in2 => \N__23207\,
            in3 => \N__23529\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_11_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23525\,
            in1 => \N__23373\,
            in2 => \N__20025\,
            in3 => \N__23150\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_18_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23370\,
            in1 => \N__23527\,
            in2 => \N__23206\,
            in3 => \N__20013\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_21_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23526\,
            in1 => \N__23374\,
            in2 => \N__20007\,
            in3 => \N__23149\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_28_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23372\,
            in1 => \N__23528\,
            in2 => \N__23208\,
            in3 => \N__19998\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49902\,
            ce => 'H',
            sr => \N__49430\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIA77M_10_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21906\,
            in1 => \N__23008\,
            in2 => \N__22938\,
            in3 => \N__22973\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_17_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21670\,
            in1 => \N__21717\,
            in2 => \N__22316\,
            in3 => \N__21779\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI288U3_23_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21907\,
            in1 => \N__22240\,
            in2 => \N__20097\,
            in3 => \N__20094\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_2_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__20929\,
            in1 => \N__21136\,
            in2 => \N__21075\,
            in3 => \N__21017\,
            lcout => \current_shift_inst.PI_CTRL.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__21016\,
            in1 => \N__20928\,
            in2 => \N__20826\,
            in3 => \N__22668\,
            lcout => \current_shift_inst.PI_CTRL.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI516M_11_LC_2_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22883\,
            in1 => \N__21868\,
            in2 => \N__21249\,
            in3 => \N__21311\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI555B_21_LC_2_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22068\,
            in2 => \_gnd_net_\,
            in3 => \N__21559\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIRGP71_5_LC_2_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__21432\,
            in1 => \N__22669\,
            in2 => \_gnd_net_\,
            in3 => \N__21469\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI23CN3_6_LC_2_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__21508\,
            in1 => \N__20088\,
            in2 => \N__20082\,
            in3 => \N__21380\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIVPSH7_10_LC_2_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20079\,
            in1 => \N__20070\,
            in2 => \N__20064\,
            in3 => \N__20136\,
            lcout => \current_shift_inst.PI_CTRL.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIOPLC1_20_LC_2_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__21618\,
            in1 => \N__20130\,
            in2 => \N__22190\,
            in3 => \N__20061\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIEE3E2_23_LC_2_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20124\,
            in1 => \N__23530\,
            in2 => \N__20139\,
            in3 => \N__22239\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIHIBM_25_LC_2_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__22594\,
            in1 => \N__22018\,
            in2 => \N__21974\,
            in3 => \N__22135\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIJG7M_0_17_LC_2_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21719\,
            in1 => \N__21674\,
            in2 => \N__22315\,
            in3 => \N__21778\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIGBD4_13_LC_2_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21194\,
            in1 => \N__22155\,
            in2 => \N__22208\,
            in3 => \N__21839\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_2_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22265\,
            in2 => \_gnd_net_\,
            in3 => \N__21530\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIIE52_10_LC_2_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21209\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIHBC4_13_LC_2_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21840\,
            in1 => \N__21639\,
            in2 => \N__21588\,
            in3 => \N__21195\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILIF4_21_LC_2_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21531\,
            in1 => \N__21888\,
            in2 => \N__22209\,
            in3 => \N__22154\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI1PR8_11_LC_2_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21279\,
            in1 => \N__21936\,
            in2 => \N__20112\,
            in3 => \N__20109\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILFC4_10_LC_2_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21800\,
            in1 => \N__21887\,
            in2 => \N__21330\,
            in3 => \N__21821\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI7RN8_11_LC_2_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21278\,
            in1 => \N__21210\,
            in2 => \N__20187\,
            in3 => \N__20154\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINJE4_19_LC_2_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22100\,
            in1 => \N__21584\,
            in2 => \N__22049\,
            in3 => \N__21638\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI0EK5_27_LC_2_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20184\,
            in1 => \N__21935\,
            in2 => \N__22562\,
            in3 => \N__21989\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0_11_LC_2_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__20169\,
            in2 => \N__20163\,
            in3 => \N__20160\,
            lcout => \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIVR52_17_LC_2_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21749\,
            in2 => \_gnd_net_\,
            in3 => \N__21692\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIPLE4_17_LC_2_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21693\,
            in1 => \N__21750\,
            in2 => \N__22563\,
            in3 => \N__21990\,
            lcout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_2_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22480\,
            in2 => \_gnd_net_\,
            in3 => \N__22375\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_2_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__22448\,
            in1 => \N__22511\,
            in2 => \N__20142\,
            in3 => \N__22415\,
            lcout => \current_shift_inst.PI_CTRL.N_31\,
            ltout => \current_shift_inst.PI_CTRL.N_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_2_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__29758\,
            in1 => \N__20890\,
            in2 => \N__20388\,
            in3 => \N__20274\,
            lcout => \current_shift_inst.PI_CTRL.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_2_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20889\,
            in2 => \_gnd_net_\,
            in3 => \N__20974\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_2_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__29764\,
            in1 => \N__22340\,
            in2 => \N__20379\,
            in3 => \N__20370\,
            lcout => \current_shift_inst.PI_CTRL.N_96\,
            ltout => \current_shift_inst.PI_CTRL.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_2_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__20975\,
            in1 => \N__20253\,
            in2 => \N__20337\,
            in3 => \N__20321\,
            lcout => \current_shift_inst.PI_CTRL.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_2_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__29763\,
            in1 => \N__20309\,
            in2 => \N__20894\,
            in3 => \N__20281\,
            lcout => \current_shift_inst.PI_CTRL.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_1_0_LC_2_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__20612\,
            in1 => \N__20584\,
            in2 => \N__20505\,
            in3 => \N__20632\,
            lcout => \pwm_generator_inst.un2_duty_input_0_o3_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_2_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__29762\,
            in1 => \N__20310\,
            in2 => \_gnd_net_\,
            in3 => \N__20280\,
            lcout => \current_shift_inst.PI_CTRL.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o2_1_LC_2_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__20246\,
            in1 => \N__20543\,
            in2 => \N__20231\,
            in3 => \N__20210\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_LC_2_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111101"
        )
    port map (
            in0 => \N__20561\,
            in1 => \N__20196\,
            in2 => \N__20190\,
            in3 => \N__20524\,
            lcout => \pwm_generator_inst.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_3_LC_2_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20633\,
            in1 => \N__20608\,
            in2 => \N__20589\,
            in3 => \N__20560\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un2_duty_input_0_o3_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_duty_input_0_o3_0_LC_2_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__20542\,
            in1 => \N__20525\,
            in2 => \N__20508\,
            in3 => \N__20497\,
            lcout => \pwm_generator_inst.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_0_c_inv_LC_2_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20466\,
            in2 => \_gnd_net_\,
            in3 => \N__20478\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_2_24_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_1_c_inv_LC_2_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20448\,
            in2 => \_gnd_net_\,
            in3 => \N__20460\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_0\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_2_c_inv_LC_2_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20430\,
            in2 => \_gnd_net_\,
            in3 => \N__20442\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_1\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_3_c_inv_LC_2_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20412\,
            in2 => \_gnd_net_\,
            in3 => \N__20424\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_2\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_4_c_inv_LC_2_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20394\,
            in2 => \_gnd_net_\,
            in3 => \N__20406\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_3\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_5_c_inv_LC_2_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20724\,
            in2 => \_gnd_net_\,
            in3 => \N__20736\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_4\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_6_c_inv_LC_2_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20706\,
            in2 => \_gnd_net_\,
            in3 => \N__20718\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_5\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_7_c_inv_LC_2_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20688\,
            in2 => \_gnd_net_\,
            in3 => \N__20700\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_6\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_8_c_inv_LC_2_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20670\,
            in2 => \_gnd_net_\,
            in3 => \N__20682\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_8\,
            ltout => OPEN,
            carryin => \bfn_2_25_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_inv_LC_2_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20652\,
            in2 => \_gnd_net_\,
            in3 => \N__20664\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_8\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_THRU_LUT4_0_LC_2_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23893\,
            in2 => \_gnd_net_\,
            in3 => \N__20646\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_9\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_10_c_RNIN8RS1_LC_2_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100110011"
        )
    port map (
            in0 => \N__24745\,
            in1 => \N__23841\,
            in2 => \_gnd_net_\,
            in3 => \N__20643\,
            lcout => \pwm_generator_inst.un19_threshold_axb_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_10\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_THRU_LUT4_0_LC_2_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23966\,
            in2 => \_gnd_net_\,
            in3 => \N__20640\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_11\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_THRU_LUT4_0_LC_2_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24093\,
            in2 => \_gnd_net_\,
            in3 => \N__20637\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_12\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_THRU_LUT4_0_LC_2_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24122\,
            in2 => \_gnd_net_\,
            in3 => \N__20772\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_13\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_THRU_LUT4_0_LC_2_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22784\,
            in2 => \_gnd_net_\,
            in3 => \N__20769\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_14\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_THRU_LUT4_0_LC_2_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22810\,
            in2 => \_gnd_net_\,
            in3 => \N__20766\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_2_26_0_\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_THRU_LUT4_0_LC_2_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22719\,
            in2 => \_gnd_net_\,
            in3 => \N__20763\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_16_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_16\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_THRU_LUT4_0_LC_2_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22757\,
            in2 => \_gnd_net_\,
            in3 => \N__20760\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_17_THRU_CO\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un15_threshold_1_cry_17\,
            carryout => \pwm_generator_inst.un15_threshold_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_THRU_LUT4_0_LC_2_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20757\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_inv_LC_2_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__22758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23715\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.N_88_i_i_LC_2_30_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__35105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49477\,
            lcout => \N_88_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_2_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__20745\,
            in1 => \N__23418\,
            in2 => \_gnd_net_\,
            in3 => \N__23221\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49414\
        );

    \current_shift_inst.PI_CTRL.integrator_8_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000001010001"
        )
    port map (
            in0 => \N__23598\,
            in1 => \N__23419\,
            in2 => \N__20817\,
            in3 => \N__23222\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49925\,
            ce => 'H',
            sr => \N__49414\
        );

    \current_shift_inst.PI_CTRL.prop_term_5_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29213\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49419\
        );

    \current_shift_inst.PI_CTRL.integrator_10_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23592\,
            in1 => \N__23381\,
            in2 => \N__20805\,
            in3 => \N__23217\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49419\
        );

    \current_shift_inst.PI_CTRL.prop_term_6_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29192\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49419\
        );

    \current_shift_inst.PI_CTRL.integrator_15_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111000001100"
        )
    port map (
            in0 => \N__23380\,
            in1 => \N__23593\,
            in2 => \N__23242\,
            in3 => \N__20793\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49419\
        );

    \current_shift_inst.PI_CTRL.prop_term_2_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__28688\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49913\,
            ce => 'H',
            sr => \N__49419\
        );

    \current_shift_inst.PI_CTRL.integrator_9_LC_3_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010101011"
        )
    port map (
            in0 => \N__20784\,
            in1 => \N__23427\,
            in2 => \N__23240\,
            in3 => \N__23597\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49423\
        );

    \current_shift_inst.PI_CTRL.prop_term_3_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28664\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49423\
        );

    \current_shift_inst.PI_CTRL.prop_term_9_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29102\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49423\
        );

    \current_shift_inst.PI_CTRL.prop_term_0_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30803\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49903\,
            ce => 'H',
            sr => \N__49423\
        );

    \current_shift_inst.PI_CTRL.prop_term_18_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29327\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49428\
        );

    \current_shift_inst.PI_CTRL.prop_term_4_LC_3_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29244\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49428\
        );

    \current_shift_inst.PI_CTRL.integrator_6_LC_3_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001000101"
        )
    port map (
            in0 => \N__23591\,
            in1 => \N__20838\,
            in2 => \N__23417\,
            in3 => \N__23151\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49428\
        );

    \current_shift_inst.PI_CTRL.prop_term_22_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29678\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49428\
        );

    \current_shift_inst.PI_CTRL.prop_term_10_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29072\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49428\
        );

    \current_shift_inst.PI_CTRL.prop_term_12_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29009\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49890\,
            ce => 'H',
            sr => \N__49428\
        );

    \current_shift_inst.PI_CTRL.integrator_RNII42L1_6_LC_3_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__21423\,
            in1 => \N__21495\,
            in2 => \N__21470\,
            in3 => \N__21366\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI34BM_20_LC_3_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23552\,
            in1 => \N__22186\,
            in2 => \N__21566\,
            in3 => \N__21620\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNIMMAM_25_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22076\,
            in1 => \N__22019\,
            in2 => \N__21970\,
            in3 => \N__22128\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI1V2B_11_LC_3_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21872\,
            in2 => \_gnd_net_\,
            in3 => \N__21306\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI71EC1_12_LC_3_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22595\,
            in1 => \N__21257\,
            in2 => \N__21183\,
            in3 => \N__22848\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI24CN6_12_LC_3_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21180\,
            in1 => \N__21174\,
            in2 => \N__21168\,
            in3 => \N__21165\,
            lcout => \current_shift_inst.PI_CTRL.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_3_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21159\,
            in2 => \N__21141\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_3_17_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_2_LC_3_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21087\,
            in2 => \N__21074\,
            in3 => \N__21024\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_3_LC_3_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21021\,
            in2 => \N__20991\,
            in3 => \N__20946\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_4_LC_3_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20943\,
            in2 => \N__20934\,
            in3 => \N__20856\,
            lcout => \current_shift_inst.PI_CTRL.un7_enablelto4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_5_LC_3_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20853\,
            in2 => \N__22671\,
            in3 => \N__20841\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_6_LC_3_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21519\,
            in2 => \N__21510\,
            in3 => \N__21474\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_7_LC_3_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23619\,
            in2 => \N__21471\,
            in3 => \N__21435\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_8_LC_3_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23049\,
            in2 => \N__21431\,
            in3 => \N__21396\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8\,
            clk => \N__49866\,
            ce => 'H',
            sr => \N__49435\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_9_LC_3_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21393\,
            in2 => \N__21384\,
            in3 => \N__21342\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_3_18_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_10_LC_3_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21339\,
            in2 => \N__22934\,
            in3 => \N__21318\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_11_LC_3_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22842\,
            in2 => \N__21315\,
            in3 => \N__21270\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_12_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21267\,
            in2 => \N__21258\,
            in3 => \N__21198\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_13_LC_3_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23040\,
            in2 => \N__22977\,
            in3 => \N__21186\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_14_LC_3_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22836\,
            in2 => \N__21876\,
            in3 => \N__21831\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_15_LC_3_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23028\,
            in2 => \N__23016\,
            in3 => \N__21810\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_16_LC_3_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23679\,
            in2 => \N__22890\,
            in3 => \N__21789\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16\,
            clk => \N__49855\,
            ce => 'H',
            sr => \N__49439\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_17_LC_3_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24045\,
            in2 => \N__21786\,
            in3 => \N__21741\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_3_19_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_18_LC_3_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21738\,
            in2 => \N__21726\,
            in3 => \N__21681\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_19_LC_3_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23640\,
            in2 => \N__21678\,
            in3 => \N__21627\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_20_LC_3_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21624\,
            in2 => \N__23634\,
            in3 => \N__21573\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_21_LC_3_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22542\,
            in2 => \N__21570\,
            in3 => \N__21522\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_22_LC_3_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22329\,
            in2 => \N__22320\,
            in3 => \N__22254\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_23_LC_3_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23652\,
            in2 => \N__22251\,
            in3 => \N__22194\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_24_LC_3_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22191\,
            in2 => \N__23691\,
            in3 => \N__22146\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24\,
            clk => \N__49843\,
            ce => 'H',
            sr => \N__49442\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_25_LC_3_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23673\,
            in2 => \N__22143\,
            in3 => \N__22089\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_3_20_0_\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_26_LC_3_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23625\,
            in2 => \N__22086\,
            in3 => \N__22032\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_27_LC_3_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23646\,
            in2 => \N__22029\,
            in3 => \N__21981\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_28_LC_3_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24033\,
            in2 => \N__21978\,
            in3 => \N__21924\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_29_LC_3_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23664\,
            in2 => \N__21921\,
            in3 => \N__21879\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_30_LC_3_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24018\,
            in2 => \N__22602\,
            in3 => \N__22548\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30\,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_31_LC_3_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__23590\,
            in1 => \N__29796\,
            in2 => \_gnd_net_\,
            in3 => \N__22545\,
            lcout => \current_shift_inst.PI_CTRL.un8_enablelto31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.prop_term_21_LC_3_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29712\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49833\,
            ce => 'H',
            sr => \N__49445\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_0_LC_3_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22536\,
            lcout => \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49826\,
            ce => 'H',
            sr => \N__49450\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIT0LD_6_LC_3_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22504\,
            in2 => \_gnd_net_\,
            in3 => \N__22485\,
            lcout => OPEN,
            ltout => \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_3_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22447\,
            in1 => \N__22414\,
            in2 => \N__22389\,
            in3 => \N__22382\,
            lcout => \current_shift_inst.PI_CTRL.N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_inv_LC_3_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22717\,
            in2 => \_gnd_net_\,
            in3 => \N__23729\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_inv_LC_3_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23765\,
            in2 => \_gnd_net_\,
            in3 => \N__22783\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_inv_LC_3_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23939\,
            in2 => \_gnd_net_\,
            in3 => \N__23965\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_inv_LC_3_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__24146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24121\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBK93_LC_3_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23865\,
            in2 => \N__24771\,
            in3 => \N__24770\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIGBKZ0Z93\,
            ltout => OPEN,
            carryin => \bfn_3_24_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7C2_LC_3_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22629\,
            in2 => \_gnd_net_\,
            in3 => \N__22623\,
            lcout => \pwm_generator_inst.un19_threshold_cry_0_c_RNIJK7CZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_0\,
            carryout => \pwm_generator_inst.un19_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9D2_LC_3_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23928\,
            in2 => \_gnd_net_\,
            in3 => \N__22620\,
            lcout => \pwm_generator_inst.un19_threshold_cry_1_c_RNIQB9DZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_1\,
            carryout => \pwm_generator_inst.un19_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCD2_LC_3_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24051\,
            in2 => \_gnd_net_\,
            in3 => \N__22617\,
            lcout => \pwm_generator_inst.un19_threshold_cry_2_c_RNITHCDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_2\,
            carryout => \pwm_generator_inst.un19_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFD2_LC_3_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24099\,
            in2 => \_gnd_net_\,
            in3 => \N__22614\,
            lcout => \pwm_generator_inst.un19_threshold_cry_3_c_RNI0OFDZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_3\,
            carryout => \pwm_generator_inst.un19_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BR2_LC_3_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22764\,
            in2 => \_gnd_net_\,
            in3 => \N__22611\,
            lcout => \pwm_generator_inst.un19_threshold_cry_4_c_RNIH7BRZ0Z2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_4\,
            carryout => \pwm_generator_inst.un19_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLN23_LC_3_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22797\,
            in2 => \_gnd_net_\,
            in3 => \N__22608\,
            lcout => \pwm_generator_inst.un19_threshold_cry_5_c_RNIGLNZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_5\,
            carryout => \pwm_generator_inst.un19_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTR23_LC_3_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22692\,
            in2 => \_gnd_net_\,
            in3 => \N__22605\,
            lcout => \pwm_generator_inst.un19_threshold_cry_6_c_RNIKTRZ0Z23\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un19_threshold_cry_6\,
            carryout => \pwm_generator_inst.un19_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNIO5033_LC_3_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22731\,
            in2 => \_gnd_net_\,
            in3 => \N__22830\,
            lcout => \pwm_generator_inst.un19_threshold_cry_7_c_RNIOZ0Z5033\,
            ltout => OPEN,
            carryin => \bfn_3_25_0_\,
            carryout => \pwm_generator_inst.un19_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISD433_LC_3_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000011101111000"
        )
    port map (
            in0 => \N__24755\,
            in1 => \N__22827\,
            in2 => \N__23859\,
            in3 => \N__22821\,
            lcout => \pwm_generator_inst.un15_threshold_1_cry_18_c_RNISDZ0Z433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_inv_LC_3_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__22812\,
            in1 => \_gnd_net_\,
            in2 => \N__23751\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_15_c_RNIFV5J2_LC_3_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110001011100"
        )
    port map (
            in0 => \N__22818\,
            in1 => \N__23750\,
            in2 => \N__24765\,
            in3 => \N__22811\,
            lcout => \pwm_generator_inst.un19_threshold_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_14_c_RNIHJQB2_LC_3_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111110010000"
        )
    port map (
            in0 => \N__22791\,
            in1 => \N__22785\,
            in2 => \N__24764\,
            in3 => \N__23772\,
            lcout => \pwm_generator_inst.un19_threshold_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_17_c_RNILBCJ2_LC_3_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__24757\,
            in1 => \N__22756\,
            in2 => \N__22743\,
            in3 => \N__23714\,
            lcout => \pwm_generator_inst.un19_threshold_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_16_c_RNII59J2_LC_3_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000111010"
        )
    port map (
            in0 => \N__23733\,
            in1 => \N__22725\,
            in2 => \N__24766\,
            in3 => \N__22718\,
            lcout => \pwm_generator_inst.un19_threshold_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.integrator_5_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001010100011"
        )
    port map (
            in0 => \N__22686\,
            in1 => \N__23588\,
            in2 => \N__23247\,
            in3 => \N__23430\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49415\
        );

    \current_shift_inst.PI_CTRL.prop_term_7_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29162\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49415\
        );

    \current_shift_inst.PI_CTRL.integrator_13_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110101000"
        )
    port map (
            in0 => \N__23607\,
            in1 => \N__23429\,
            in2 => \N__23246\,
            in3 => \N__23589\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49904\,
            ce => 'H',
            sr => \N__49415\
        );

    \current_shift_inst.PI_CTRL.integrator_16_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011101010"
        )
    port map (
            in0 => \N__23587\,
            in1 => \N__23428\,
            in2 => \N__23262\,
            in3 => \N__23205\,
            lcout => \current_shift_inst.PI_CTRL.integratorZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.prop_term_8_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29135\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.prop_term_13_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29468\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.prop_term_15_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29411\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49891\,
            ce => 'H',
            sr => \N__49420\
        );

    \current_shift_inst.PI_CTRL.integrator_RNI626M_10_LC_4_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23012\,
            in1 => \N__22969\,
            in2 => \N__22933\,
            in3 => \N__22881\,
            lcout => \current_shift_inst.PI_CTRL.un3_enable_0_a3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.prop_term_11_LC_4_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29039\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.prop_term_14_LC_4_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29444\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.prop_term_24_LC_4_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29628\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49856\,
            ce => 'H',
            sr => \N__49431\
        );

    \current_shift_inst.PI_CTRL.prop_term_16_LC_4_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29390\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \N__49436\
        );

    \current_shift_inst.PI_CTRL.prop_term_25_LC_4_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29594\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \N__49436\
        );

    \current_shift_inst.PI_CTRL.prop_term_29_LC_4_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29865\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49844\,
            ce => 'H',
            sr => \N__49436\
        );

    \current_shift_inst.PI_CTRL.prop_term_23_LC_4_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29655\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \N__49440\
        );

    \current_shift_inst.PI_CTRL.prop_term_27_LC_4_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29531\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \N__49440\
        );

    \current_shift_inst.PI_CTRL.prop_term_19_LC_4_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29303\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \N__49440\
        );

    \current_shift_inst.PI_CTRL.prop_term_20_LC_4_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29271\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49834\,
            ce => 'H',
            sr => \N__49440\
        );

    \current_shift_inst.PI_CTRL.prop_term_26_LC_4_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29564\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49827\,
            ce => 'H',
            sr => \N__49443\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_LC_4_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23840\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_22_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5C_LC_4_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23817\,
            in2 => \_gnd_net_\,
            in3 => \N__23805\,
            lcout => \pwm_generator_inst.un3_threshold_cry_0_c_RNI2R5CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_0\,
            carryout => \pwm_generator_inst.un3_threshold_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6C_LC_4_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23802\,
            in2 => \_gnd_net_\,
            in3 => \N__23790\,
            lcout => \pwm_generator_inst.un3_threshold_cry_1_c_RNI3T6CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_1\,
            carryout => \pwm_generator_inst.un3_threshold_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7C_LC_4_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23787\,
            in2 => \_gnd_net_\,
            in3 => \N__23775\,
            lcout => \pwm_generator_inst.un3_threshold_cry_2_c_RNI4V7CZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_2\,
            carryout => \pwm_generator_inst.un3_threshold_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1Q_LC_4_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24399\,
            in2 => \_gnd_net_\,
            in3 => \N__23754\,
            lcout => \pwm_generator_inst.un3_threshold_cry_3_c_RNIJA1QZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_3\,
            carryout => \pwm_generator_inst.un3_threshold_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKB11_LC_4_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24357\,
            in2 => \N__38572\,
            in3 => \N__23736\,
            lcout => \pwm_generator_inst.un3_threshold_cry_4_c_RNIGKBZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_4\,
            carryout => \pwm_generator_inst.un3_threshold_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_5_c_RNIIOD11_LC_4_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38531\,
            in2 => \N__24315\,
            in3 => \N__23718\,
            lcout => \pwm_generator_inst.un3_threshold_cry_5_c_RNIIODZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_5\,
            carryout => \pwm_generator_inst.un3_threshold_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSF11_LC_4_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24273\,
            in2 => \N__38573\,
            in3 => \N__23694\,
            lcout => \pwm_generator_inst.un3_threshold_cry_6_c_RNIKSFZ0Z11\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_6\,
            carryout => \pwm_generator_inst.un3_threshold_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0I11_LC_4_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24237\,
            in2 => \_gnd_net_\,
            in3 => \N__23844\,
            lcout => \pwm_generator_inst.un3_threshold_cry_7_c_RNIM0IZ0Z11\,
            ltout => OPEN,
            carryin => \bfn_4_23_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_LC_4_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24198\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_8\,
            carryout => \pwm_generator_inst.un3_threshold_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_LC_4_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24159\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_9\,
            carryout => \pwm_generator_inst.un3_threshold_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_LC_4_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24660\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_10\,
            carryout => \pwm_generator_inst.un3_threshold_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_LC_4_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24615\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_11\,
            carryout => \pwm_generator_inst.un3_threshold_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_LC_4_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24570\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_12\,
            carryout => \pwm_generator_inst.un3_threshold_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_LC_4_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24540\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_13\,
            carryout => \pwm_generator_inst.un3_threshold_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_LC_4_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24516\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_14\,
            carryout => \pwm_generator_inst.un3_threshold_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_LC_4_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24492\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_24_0_\,
            carryout => \pwm_generator_inst.un3_threshold_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_LC_4_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24471\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_16\,
            carryout => \pwm_generator_inst.un3_threshold_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_LC_4_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24441\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_17\,
            carryout => \pwm_generator_inst.un3_threshold_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_LC_4_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24789\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un3_threshold_cry_18\,
            carryout => \pwm_generator_inst.un3_threshold_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_THRU_LUT4_0_LC_4_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24006\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_4_c_RNI5DBP6_LC_4_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__26984\,
            in1 => \N__24003\,
            in2 => \N__48870\,
            in3 => \N__26918\,
            lcout => \pwm_generator_inst.threshold_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_1_c_RNIEH9B6_LC_4_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__26983\,
            in1 => \N__23997\,
            in2 => \N__48869\,
            in3 => \N__26917\,
            lcout => \pwm_generator_inst.threshold_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_18_c_RNIGJ417_LC_4_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__26989\,
            in1 => \N__48780\,
            in2 => \N__23991\,
            in3 => \N__26919\,
            lcout => \pwm_generator_inst.threshold_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_11_c_RNITTRT1_LC_4_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__24737\,
            in1 => \N__23979\,
            in2 => \N__23970\,
            in3 => \N__23943\,
            lcout => \pwm_generator_inst.un19_threshold_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNIFGO02_LC_4_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001110101010"
        )
    port map (
            in0 => \N__23922\,
            in1 => \N__23904\,
            in2 => \N__23877\,
            in3 => \N__24736\,
            lcout => \pwm_generator_inst.un19_threshold_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_RNI160U1_LC_4_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001001110"
        )
    port map (
            in0 => \N__24738\,
            in1 => \N__24150\,
            in2 => \N__24135\,
            in3 => \N__24123\,
            lcout => \pwm_generator_inst.un19_threshold_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_13_c_inv_LC_4_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__24092\,
            in1 => \_gnd_net_\,
            in2 => \N__24066\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un15_threshold_1_axb_13\,
            ltout => \pwm_generator_inst.un15_threshold_1_axb_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un15_threshold_1_cry_12_c_RNIV1UT1_LC_4_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011110000010"
        )
    port map (
            in0 => \N__24756\,
            in1 => \N__24078\,
            in2 => \N__24069\,
            in3 => \N__24065\,
            lcout => \pwm_generator_inst.un19_threshold_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_30_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010001110"
        )
    port map (
            in0 => \N__25782\,
            in1 => \N__28194\,
            in2 => \N__25763\,
            in3 => \N__28221\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_15_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24852\,
            in1 => \N__26397\,
            in2 => \_gnd_net_\,
            in3 => \N__36681\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49950\,
            ce => \N__33338\,
            sr => \N__49384\
        );

    \current_shift_inst.PI_CTRL.prop_term_17_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29357\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49867\,
            ce => 'H',
            sr => \N__49421\
        );

    \current_shift_inst.PI_CTRL.prop_term_28_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29492\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49857\,
            ce => 'H',
            sr => \N__49424\
        );

    \current_shift_inst.PI_CTRL.prop_term_30_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29834\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49835\,
            ce => 'H',
            sr => \N__49432\
        );

    \CONSTANT_ONE_LUT4_LC_5_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_axb_4_LC_5_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24432\,
            in2 => \N__24417\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.un3_threshold_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \bfn_5_23_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7P701_LC_5_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24393\,
            in2 => \N__24375\,
            in3 => \N__24351\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_0_c_RNI7PZ0Z701\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_0\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8R801_LC_5_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24348\,
            in2 => \N__24333\,
            in3 => \N__24306\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_1_c_RNI8RZ0Z801\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_1\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9T901_LC_5_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24303\,
            in2 => \N__24288\,
            in3 => \N__24267\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_2_c_RNI9TZ0Z901\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_2\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVA01_LC_5_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24264\,
            in2 => \N__24252\,
            in3 => \N__24231\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_3_c_RNIAVAZ0Z01\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_3\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_9_c_RNO_LC_5_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24228\,
            in2 => \N__24216\,
            in3 => \N__24192\,
            lcout => \pwm_generator_inst.un3_threshold_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_4\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_10_c_RNO_LC_5_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24189\,
            in2 => \N__24174\,
            in3 => \N__24153\,
            lcout => \pwm_generator_inst.un3_threshold_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_5\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_11_c_RNO_LC_5_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24690\,
            in2 => \N__24675\,
            in3 => \N__24654\,
            lcout => \pwm_generator_inst.un3_threshold_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_6\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_12_c_RNO_LC_5_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24651\,
            in2 => \N__24636\,
            in3 => \N__24609\,
            lcout => \pwm_generator_inst.un3_threshold_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \bfn_5_24_0_\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_13_c_RNO_LC_5_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24606\,
            in2 => \N__24591\,
            in3 => \N__24564\,
            lcout => \pwm_generator_inst.un3_threshold_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_8\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_14_c_RNO_LC_5_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48936\,
            in2 => \N__24561\,
            in3 => \N__24534\,
            lcout => \pwm_generator_inst.un3_threshold_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_9\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_15_c_RNO_LC_5_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24531\,
            in2 => \N__48951\,
            in3 => \N__24510\,
            lcout => \pwm_generator_inst.un3_threshold_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_10\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_16_c_RNO_LC_5_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48940\,
            in2 => \N__24507\,
            in3 => \N__24486\,
            lcout => \pwm_generator_inst.un3_threshold_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_11\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_17_c_RNO_LC_5_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24483\,
            in2 => \N__48952\,
            in3 => \N__24465\,
            lcout => \pwm_generator_inst.un3_threshold_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_12\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_18_c_RNO_LC_5_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48944\,
            in2 => \N__24462\,
            in3 => \N__24435\,
            lcout => \pwm_generator_inst.un3_threshold_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_13\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un3_threshold_cry_19_c_RNO_LC_5_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48663\,
            in2 => \N__48953\,
            in3 => \N__24783\,
            lcout => \pwm_generator_inst.un3_threshold_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un2_threshold_add_1_cry_14\,
            carryout => \pwm_generator_inst.un2_threshold_add_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RR81_LC_5_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__24780\,
            in1 => \N__30693\,
            in2 => \_gnd_net_\,
            in3 => \N__24774\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_cry_15_c_RNI1RRZ0Z81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_11_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24896\,
            in1 => \N__25994\,
            in2 => \_gnd_net_\,
            in3 => \N__36649\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__31249\,
            sr => \N__49340\
        );

    \phase_controller_inst1.stoper_tr.target_time_15_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36645\,
            in1 => \N__24848\,
            in2 => \_gnd_net_\,
            in3 => \N__26396\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__31249\,
            sr => \N__49340\
        );

    \phase_controller_inst1.stoper_tr.target_time_7_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__26142\,
            in1 => \_gnd_net_\,
            in2 => \N__36703\,
            in3 => \N__24913\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__31249\,
            sr => \N__49340\
        );

    \phase_controller_inst1.stoper_tr.target_time_5_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30228\,
            in1 => \N__30185\,
            in2 => \_gnd_net_\,
            in3 => \N__36650\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49956\,
            ce => \N__31249\,
            sr => \N__49340\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_18_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__24824\,
            in1 => \N__28076\,
            in2 => \N__24809\,
            in3 => \N__28109\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24917\,
            in1 => \N__26141\,
            in2 => \_gnd_net_\,
            in3 => \N__36632\,
            lcout => \elapsed_time_ns_1_RNIJI91B_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_18_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__24825\,
            in1 => \N__28077\,
            in2 => \N__24810\,
            in3 => \N__28110\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30223\,
            in1 => \N__30184\,
            in2 => \_gnd_net_\,
            in3 => \N__36637\,
            lcout => \elapsed_time_ns_1_RNIHG91B_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36636\,
            in1 => \N__24895\,
            in2 => \_gnd_net_\,
            in3 => \N__25998\,
            lcout => \elapsed_time_ns_1_RNIU7OBB_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_20_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__28050\,
            in1 => \N__25889\,
            in2 => \N__28029\,
            in3 => \N__24933\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_20_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__24932\,
            in1 => \N__28024\,
            in2 => \N__25893\,
            in3 => \N__28049\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24847\,
            in1 => \N__26389\,
            in2 => \_gnd_net_\,
            in3 => \N__36651\,
            lcout => \elapsed_time_ns_1_RNI2COBB_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_18_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31307\,
            in1 => \N__31356\,
            in2 => \_gnd_net_\,
            in3 => \N__36602\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49946\,
            ce => \N__31248\,
            sr => \N__49370\
        );

    \phase_controller_inst1.stoper_tr.target_time_2_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28508\,
            in1 => \N__28481\,
            in2 => \_gnd_net_\,
            in3 => \N__36603\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49946\,
            ce => \N__31248\,
            sr => \N__49370\
        );

    \phase_controller_inst1.stoper_tr.target_time_19_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36545\,
            in1 => \N__28799\,
            in2 => \_gnd_net_\,
            in3 => \N__28776\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49936\,
            ce => \N__31200\,
            sr => \N__49374\
        );

    \phase_controller_inst1.stoper_tr.target_time_30_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30893\,
            in1 => \N__30920\,
            in2 => \_gnd_net_\,
            in3 => \N__36546\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49936\,
            ce => \N__31200\,
            sr => \N__49374\
        );

    \phase_controller_inst1.stoper_tr.target_time_31_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36469\,
            in1 => \N__28974\,
            in2 => \_gnd_net_\,
            in3 => \N__28936\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__31255\,
            sr => \N__49380\
        );

    \phase_controller_inst1.stoper_tr.target_time_20_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33159\,
            in1 => \N__33203\,
            in2 => \_gnd_net_\,
            in3 => \N__36470\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__31255\,
            sr => \N__49380\
        );

    \phase_controller_inst1.stoper_tr.target_time_23_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__25874\,
            in1 => \_gnd_net_\,
            in2 => \N__26682\,
            in3 => \N__36471\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49926\,
            ce => \N__31255\,
            sr => \N__49380\
        );

    \phase_controller_inst2.stoper_tr.target_time_7_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36464\,
            in1 => \N__24921\,
            in2 => \_gnd_net_\,
            in3 => \N__26140\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__33339\,
            sr => \N__49385\
        );

    \phase_controller_inst2.stoper_tr.target_time_22_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36462\,
            in1 => \N__26742\,
            in2 => \_gnd_net_\,
            in3 => \N__25713\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__33339\,
            sr => \N__49385\
        );

    \phase_controller_inst2.stoper_tr.target_time_11_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__24897\,
            in1 => \N__25993\,
            in2 => \_gnd_net_\,
            in3 => \N__36465\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__33339\,
            sr => \N__49385\
        );

    \phase_controller_inst2.stoper_tr.target_time_23_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26681\,
            in1 => \N__25873\,
            in2 => \_gnd_net_\,
            in3 => \N__36466\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__33339\,
            sr => \N__49385\
        );

    \phase_controller_inst2.stoper_tr.target_time_25_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36463\,
            in1 => \N__26589\,
            in2 => \_gnd_net_\,
            in3 => \N__25635\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49914\,
            ce => \N__33339\,
            sr => \N__49385\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_22_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011010100"
        )
    port map (
            in0 => \N__31772\,
            in1 => \N__24873\,
            in2 => \N__24864\,
            in3 => \N__31796\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_22_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__24872\,
            in1 => \N__31773\,
            in2 => \N__31797\,
            in3 => \N__24863\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25931\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49892\,
            ce => \N__27061\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26240\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49892\,
            ce => \N__27061\,
            sr => \N__49393\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36477\,
            in1 => \N__28504\,
            in2 => \_gnd_net_\,
            in3 => \N__28470\,
            lcout => \elapsed_time_ns_1_RNIED91B_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36478\,
            in1 => \N__30916\,
            in2 => \_gnd_net_\,
            in3 => \N__30889\,
            lcout => \elapsed_time_ns_1_RNIVAQBB_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25115\,
            in1 => \N__25921\,
            in2 => \_gnd_net_\,
            in3 => \N__24951\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25103\,
            in1 => \N__26230\,
            in2 => \_gnd_net_\,
            in3 => \N__24948\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25116\,
            in1 => \N__26204\,
            in2 => \_gnd_net_\,
            in3 => \N__24945\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25104\,
            in1 => \N__26185\,
            in2 => \_gnd_net_\,
            in3 => \N__24942\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25117\,
            in1 => \N__26158\,
            in2 => \_gnd_net_\,
            in3 => \N__24939\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25105\,
            in1 => \N__26098\,
            in2 => \_gnd_net_\,
            in3 => \N__24936\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25118\,
            in1 => \N__26074\,
            in2 => \_gnd_net_\,
            in3 => \N__24978\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25106\,
            in1 => \N__26041\,
            in2 => \_gnd_net_\,
            in3 => \N__24975\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_7\,
            clk => \N__49868\,
            ce => \N__25160\,
            sr => \N__49401\
        );

    \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25102\,
            in1 => \N__26017\,
            in2 => \_gnd_net_\,
            in3 => \N__24972\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25114\,
            in1 => \N__26491\,
            in2 => \_gnd_net_\,
            in3 => \N__24969\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25099\,
            in1 => \N__26461\,
            in2 => \_gnd_net_\,
            in3 => \N__24966\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25111\,
            in1 => \N__26432\,
            in2 => \_gnd_net_\,
            in3 => \N__24963\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25100\,
            in1 => \N__26413\,
            in2 => \_gnd_net_\,
            in3 => \N__24960\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25112\,
            in1 => \N__26344\,
            in2 => \_gnd_net_\,
            in3 => \N__24957\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__26312\,
            in2 => \_gnd_net_\,
            in3 => \N__24954\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25113\,
            in1 => \N__26290\,
            in2 => \_gnd_net_\,
            in3 => \N__25005\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_15\,
            clk => \N__49858\,
            ce => \N__25161\,
            sr => \N__49407\
        );

    \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25107\,
            in1 => \N__26263\,
            in2 => \_gnd_net_\,
            in3 => \N__25002\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25119\,
            in1 => \N__26803\,
            in2 => \_gnd_net_\,
            in3 => \N__24999\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25108\,
            in1 => \N__26779\,
            in2 => \_gnd_net_\,
            in3 => \N__24996\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25120\,
            in1 => \N__26758\,
            in2 => \_gnd_net_\,
            in3 => \N__24993\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25109\,
            in1 => \N__26698\,
            in2 => \_gnd_net_\,
            in3 => \N__24990\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25121\,
            in1 => \N__26630\,
            in2 => \_gnd_net_\,
            in3 => \N__24987\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25110\,
            in1 => \N__26605\,
            in2 => \_gnd_net_\,
            in3 => \N__24984\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25122\,
            in1 => \N__26545\,
            in2 => \_gnd_net_\,
            in3 => \N__24981\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_23\,
            clk => \N__49845\,
            ce => \N__25159\,
            sr => \N__49410\
        );

    \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25093\,
            in1 => \N__26521\,
            in2 => \_gnd_net_\,
            in3 => \N__25179\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_7_16_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            clk => \N__49836\,
            ce => \N__25149\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25097\,
            in1 => \N__27172\,
            in2 => \_gnd_net_\,
            in3 => \N__25176\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            clk => \N__49836\,
            ce => \N__25149\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25094\,
            in1 => \N__27130\,
            in2 => \_gnd_net_\,
            in3 => \N__25173\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            clk => \N__49836\,
            ce => \N__25149\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25098\,
            in1 => \N__27088\,
            in2 => \_gnd_net_\,
            in3 => \N__25170\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            clk => \N__49836\,
            ce => \N__25149\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__25095\,
            in1 => \N__27149\,
            in2 => \_gnd_net_\,
            in3 => \N__25167\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.counter_cry_28\,
            clk => \N__49836\,
            ce => \N__25149\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__27107\,
            in1 => \N__25096\,
            in2 => \_gnd_net_\,
            in3 => \N__25164\,
            lcout => \delay_measurement_inst.delay_tr_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49836\,
            ce => \N__25149\,
            sr => \N__49416\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__25313\,
            in1 => \_gnd_net_\,
            in2 => \N__25296\,
            in3 => \N__25274\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_166_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25312\,
            in2 => \_gnd_net_\,
            in3 => \N__25292\,
            lcout => \delay_measurement_inst.delay_tr_timer.N_165_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25311\,
            lcout => \delay_measurement_inst.delay_tr_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.running_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__25314\,
            in1 => \N__25291\,
            in2 => \_gnd_net_\,
            in3 => \N__25275\,
            lcout => \delay_measurement_inst.delay_tr_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49821\,
            ce => 'H',
            sr => \N__49425\
        );

    \delay_measurement_inst.stop_timer_tr_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25273\,
            lcout => \delay_measurement_inst.stop_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25248\,
            ce => 'H',
            sr => \N__49429\
        );

    \delay_measurement_inst.start_timer_tr_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25272\,
            lcout => \delay_measurement_inst.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__25247\,
            ce => 'H',
            sr => \N__49433\
        );

    \pwm_generator_inst.un19_threshold_cry_2_c_RNIHNCB6_LC_7_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__27003\,
            in1 => \N__25236\,
            in2 => \N__48852\,
            in3 => \N__26912\,
            lcout => \pwm_generator_inst.threshold_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_3_c_RNIKTFB6_LC_7_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__26913\,
            in1 => \N__25227\,
            in2 => \N__48849\,
            in3 => \N__27004\,
            lcout => \pwm_generator_inst.threshold_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_0_c_RNI7Q7A6_LC_7_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__27002\,
            in1 => \N__25218\,
            in2 => \N__48851\,
            in3 => \N__26911\,
            lcout => \pwm_generator_inst.threshold_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_6_c_RNI83S07_LC_7_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__27006\,
            in1 => \N__26915\,
            in2 => \N__25209\,
            in3 => \N__48796\,
            lcout => \pwm_generator_inst.threshold_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_5_c_RNI4RN07_LC_7_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__26914\,
            in1 => \N__27005\,
            in2 => \N__48850\,
            in3 => \N__25197\,
            lcout => \pwm_generator_inst.threshold_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un19_threshold_cry_7_c_RNICB017_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__26990\,
            in1 => \N__25188\,
            in2 => \N__48781\,
            in3 => \N__26916\,
            lcout => \pwm_generator_inst.threshold_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_0_LC_7_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27402\,
            in1 => \N__27563\,
            in2 => \_gnd_net_\,
            in3 => \N__25341\,
            lcout => \pwm_generator_inst.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_26_0_\,
            carryout => \pwm_generator_inst.counter_cry_0\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_1_LC_7_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27387\,
            in1 => \N__27500\,
            in2 => \_gnd_net_\,
            in3 => \N__25338\,
            lcout => \pwm_generator_inst.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_0\,
            carryout => \pwm_generator_inst.counter_cry_1\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_2_LC_7_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27403\,
            in1 => \N__27542\,
            in2 => \_gnd_net_\,
            in3 => \N__25335\,
            lcout => \pwm_generator_inst.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_1\,
            carryout => \pwm_generator_inst.counter_cry_2\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_3_LC_7_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27388\,
            in1 => \N__27476\,
            in2 => \_gnd_net_\,
            in3 => \N__25332\,
            lcout => \pwm_generator_inst.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_2\,
            carryout => \pwm_generator_inst.counter_cry_3\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_4_LC_7_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27404\,
            in1 => \N__27521\,
            in2 => \_gnd_net_\,
            in3 => \N__25329\,
            lcout => \pwm_generator_inst.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_3\,
            carryout => \pwm_generator_inst.counter_cry_4\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_5_LC_7_26_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27389\,
            in1 => \N__27424\,
            in2 => \_gnd_net_\,
            in3 => \N__25326\,
            lcout => \pwm_generator_inst.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_4\,
            carryout => \pwm_generator_inst.counter_cry_5\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_6_LC_7_26_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27405\,
            in1 => \N__27448\,
            in2 => \_gnd_net_\,
            in3 => \N__25323\,
            lcout => \pwm_generator_inst.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_5\,
            carryout => \pwm_generator_inst.counter_cry_6\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_7_LC_7_26_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27390\,
            in1 => \N__27587\,
            in2 => \_gnd_net_\,
            in3 => \N__25320\,
            lcout => \pwm_generator_inst.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.counter_cry_6\,
            carryout => \pwm_generator_inst.counter_cry_7\,
            clk => \N__49805\,
            ce => 'H',
            sr => \N__49451\
        );

    \pwm_generator_inst.counter_8_LC_7_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27392\,
            in1 => \N__27629\,
            in2 => \_gnd_net_\,
            in3 => \N__25317\,
            lcout => \pwm_generator_inst.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_27_0_\,
            carryout => \pwm_generator_inst.counter_cry_8\,
            clk => \N__49801\,
            ce => 'H',
            sr => \N__49452\
        );

    \pwm_generator_inst.counter_9_LC_7_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__27608\,
            in1 => \N__27391\,
            in2 => \_gnd_net_\,
            in3 => \N__25446\,
            lcout => \pwm_generator_inst.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49801\,
            ce => 'H',
            sr => \N__49452\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_1_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27795\,
            in2 => \N__25443\,
            in3 => \N__27778\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_2_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25434\,
            in2 => \N__25422\,
            in3 => \N__27762\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29730\,
            in2 => \N__25413\,
            in3 => \N__27744\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_4_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27726\,
            in1 => \N__25656\,
            in2 => \N__25401\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_5_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25392\,
            in2 => \N__25386\,
            in3 => \N__27708\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_6_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27333\,
            in2 => \N__25374\,
            in3 => \N__27690\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_7_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25365\,
            in2 => \N__25359\,
            in3 => \N__27672\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_8_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25836\,
            in2 => \N__25350\,
            in3 => \N__27651\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_9_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29973\,
            in2 => \N__25524\,
            in3 => \N__27930\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_10_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25722\,
            in2 => \N__25515\,
            in3 => \N__27912\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_11_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25506\,
            in2 => \N__25500\,
            in3 => \N__27894\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_12_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25905\,
            in2 => \N__25491\,
            in3 => \N__27876\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_13_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27339\,
            in2 => \N__25482\,
            in3 => \N__27858\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_14_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31281\,
            in2 => \N__25470\,
            in3 => \N__27837\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_inv_15_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27816\,
            in1 => \N__25452\,
            in2 => \N__25461\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_16_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29961\,
            in2 => \N__29901\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_18_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25590\,
            in2 => \N__25584\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_20_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25572\,
            in2 => \N__25563\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_22_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25662\,
            in2 => \N__25533\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_24_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25599\,
            in2 => \N__25647\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_26_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25815\,
            in2 => \N__25827\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_28_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28173\,
            in2 => \N__28128\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_30_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25734\,
            in2 => \N__25551\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25536\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_22_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__25692\,
            in1 => \N__27983\,
            in2 => \N__25683\,
            in3 => \N__28001\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__26740\,
            in1 => \N__36633\,
            in2 => \_gnd_net_\,
            in3 => \N__25706\,
            lcout => \elapsed_time_ns_1_RNI0BPBB_0_22\,
            ltout => \elapsed_time_ns_1_RNI0BPBB_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_22_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36634\,
            in1 => \_gnd_net_\,
            in2 => \N__25695\,
            in3 => \N__26741\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49951\,
            ce => \N__31223\,
            sr => \N__49349\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_22_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__25691\,
            in1 => \N__27982\,
            in2 => \N__25682\,
            in3 => \N__28000\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_4_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28344\,
            in1 => \N__28371\,
            in2 => \_gnd_net_\,
            in3 => \N__36635\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49951\,
            ce => \N__31223\,
            sr => \N__49349\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_24_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__25845\,
            in1 => \N__27947\,
            in2 => \N__25614\,
            in3 => \N__27965\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26587\,
            in1 => \N__25628\,
            in2 => \_gnd_net_\,
            in3 => \N__36638\,
            lcout => \elapsed_time_ns_1_RNI3EPBB_0_25\,
            ltout => \elapsed_time_ns_1_RNI3EPBB_0_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_25_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36640\,
            in1 => \_gnd_net_\,
            in2 => \N__25617\,
            in3 => \N__26588\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__31211\,
            sr => \N__49358\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_24_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__25844\,
            in1 => \N__27946\,
            in2 => \N__25613\,
            in3 => \N__27964\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_24_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36639\,
            in1 => \N__28632\,
            in2 => \_gnd_net_\,
            in3 => \N__28611\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__31211\,
            sr => \N__49358\
        );

    \phase_controller_inst1.stoper_tr.target_time_8_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36641\,
            in1 => \N__31004\,
            in2 => \_gnd_net_\,
            in3 => \N__30977\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49947\,
            ce => \N__31211\,
            sr => \N__49358\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_26_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__28244\,
            in1 => \N__28265\,
            in2 => \N__25803\,
            in3 => \N__25791\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_26_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__25790\,
            in1 => \N__28243\,
            in2 => \N__28269\,
            in3 => \N__25799\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28916\,
            in1 => \N__28877\,
            in2 => \_gnd_net_\,
            in3 => \N__36542\,
            lcout => \elapsed_time_ns_1_RNI5GPBB_0_27\,
            ltout => \elapsed_time_ns_1_RNI5GPBB_0_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_27_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36544\,
            in1 => \_gnd_net_\,
            in2 => \N__25806\,
            in3 => \N__28917\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => \N__31265\,
            sr => \N__49365\
        );

    \phase_controller_inst1.stoper_tr.target_time_26_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36543\,
            in1 => \N__30632\,
            in2 => \_gnd_net_\,
            in3 => \N__30606\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49937\,
            ce => \N__31265\,
            sr => \N__49365\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_30_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__25775\,
            in1 => \N__28189\,
            in2 => \N__25764\,
            in3 => \N__28216\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25986\,
            in1 => \N__30075\,
            in2 => \N__28542\,
            in3 => \N__30145\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_10_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30076\,
            in1 => \N__30103\,
            in2 => \_gnd_net_\,
            in3 => \N__36597\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__31201\,
            sr => \N__49371\
        );

    \phase_controller_inst1.stoper_tr.target_time_12_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28563\,
            in1 => \N__28540\,
            in2 => \_gnd_net_\,
            in3 => \N__36598\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49927\,
            ce => \N__31201\,
            sr => \N__49371\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH9BP1_25_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26578\,
            in1 => \N__30744\,
            in2 => \N__30605\,
            in3 => \N__30885\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6T9P1_21_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26676\,
            in1 => \N__26731\,
            in2 => \N__28610\,
            in3 => \N__28841\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_21_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28865\,
            in1 => \N__28842\,
            in2 => \_gnd_net_\,
            in3 => \N__36472\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49915\,
            ce => \N__31254\,
            sr => \N__49375\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36417\,
            in1 => \N__25875\,
            in2 => \_gnd_net_\,
            in3 => \N__26677\,
            lcout => \elapsed_time_ns_1_RNI1CPBB_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIAT5P1_13_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__26379\,
            in1 => \N__31576\,
            in2 => \N__30264\,
            in3 => \N__32470\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__36414\,
            in1 => \N__28798\,
            in2 => \N__28775\,
            in3 => \_gnd_net_\,
            lcout => \elapsed_time_ns_1_RNI6GOBB_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1J1U1_5_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25857\,
            in1 => \N__30213\,
            in2 => \N__25941\,
            in3 => \N__28423\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__28290\,
            in1 => \N__25947\,
            in2 => \N__25848\,
            in3 => \N__28965\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3\,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28631\,
            in2 => \N__25953\,
            in3 => \N__28605\,
            lcout => \elapsed_time_ns_1_RNI2DPBB_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36415\,
            in1 => \N__28562\,
            in2 => \_gnd_net_\,
            in3 => \N__28541\,
            lcout => \elapsed_time_ns_1_RNIV8OBB_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28966\,
            in1 => \N__28937\,
            in2 => \_gnd_net_\,
            in3 => \N__36416\,
            lcout => \elapsed_time_ns_1_RNI0CQBB_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30631\,
            in1 => \N__30597\,
            in2 => \_gnd_net_\,
            in3 => \N__36406\,
            lcout => \elapsed_time_ns_1_RNI4FPBB_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31391\,
            in1 => \N__32662\,
            in2 => \N__28477\,
            in3 => \N__28362\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIRFVB1_27_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33057\,
            in2 => \N__25950\,
            in3 => \N__28910\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36407\,
            in1 => \N__28343\,
            in2 => \_gnd_net_\,
            in3 => \N__28363\,
            lcout => \elapsed_time_ns_1_RNIGF91B_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28864\,
            in1 => \N__28840\,
            in2 => \_gnd_net_\,
            in3 => \N__36408\,
            lcout => \elapsed_time_ns_1_RNIV9PBB_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIPDL7_7_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__26125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30960\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26210\,
            in2 => \N__25932\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3\,
            ltout => OPEN,
            carryin => \bfn_8_11_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26186\,
            in2 => \N__26241\,
            in3 => \N__26214\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26211\,
            in2 => \N__26165\,
            in3 => \N__26190\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26187\,
            in2 => \N__26105\,
            in3 => \N__26169\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26075\,
            in2 => \N__26166\,
            in3 => \N__26109\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26048\,
            in2 => \N__26106\,
            in3 => \N__26082\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26018\,
            in2 => \N__26079\,
            in3 => \N__26055\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26492\,
            in2 => \N__26052\,
            in3 => \N__26025\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49879\,
            ce => \N__27063\,
            sr => \N__49389\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26462\,
            in2 => \N__26022\,
            in3 => \N__25956\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11\,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26438\,
            in2 => \N__26499\,
            in3 => \N__26469\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26414\,
            in2 => \N__26466\,
            in3 => \N__26442\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26439\,
            in2 => \N__26351\,
            in3 => \N__26418\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26415\,
            in2 => \N__26324\,
            in3 => \N__26355\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26291\,
            in2 => \N__26352\,
            in3 => \N__26328\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26264\,
            in2 => \N__26325\,
            in3 => \N__26298\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26804\,
            in2 => \N__26295\,
            in3 => \N__26271\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49869\,
            ce => \N__27062\,
            sr => \N__49394\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26780\,
            in2 => \N__26268\,
            in3 => \N__26244\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26759\,
            in2 => \N__26808\,
            in3 => \N__26784\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26781\,
            in2 => \N__26709\,
            in3 => \N__26763\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26760\,
            in2 => \N__26642\,
            in3 => \N__26712\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26708\,
            in2 => \N__26612\,
            in3 => \N__26646\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26552\,
            in2 => \N__26643\,
            in3 => \N__26616\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26522\,
            in2 => \N__26613\,
            in3 => \N__26559\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27173\,
            in2 => \N__26556\,
            in3 => \N__26529\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49859\,
            ce => \N__27060\,
            sr => \N__49397\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27131\,
            in2 => \N__26526\,
            in3 => \N__26502\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49846\,
            ce => \N__27059\,
            sr => \N__49402\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27089\,
            in2 => \N__27177\,
            in3 => \N__27153\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49846\,
            ce => \N__27059\,
            sr => \N__49402\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27150\,
            in2 => \N__27135\,
            in3 => \N__27111\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49846\,
            ce => \N__27059\,
            sr => \N__49402\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27108\,
            in2 => \N__27093\,
            in3 => \N__27069\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49846\,
            ce => \N__27059\,
            sr => \N__49402\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27066\,
            lcout => \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49846\,
            ce => \N__27059\,
            sr => \N__49402\
        );

    \pwm_generator_inst.un15_threshold_1_cry_9_c_RNI4HK77_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__26988\,
            in1 => \N__26934\,
            in2 => \N__48730\,
            in3 => \N__26878\,
            lcout => \pwm_generator_inst.threshold_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_8_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26850\,
            in2 => \N__26859\,
            in3 => \N__27567\,
            lcout => \pwm_generator_inst.counter_i_0\,
            ltout => OPEN,
            carryin => \bfn_8_24_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_8_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26832\,
            in2 => \N__26844\,
            in3 => \N__27501\,
            lcout => \pwm_generator_inst.counter_i_1\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_0\,
            carryout => \pwm_generator_inst.un14_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_8_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26814\,
            in2 => \N__26826\,
            in3 => \N__27543\,
            lcout => \pwm_generator_inst.counter_i_2\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_1\,
            carryout => \pwm_generator_inst.un14_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_8_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27318\,
            in2 => \N__27327\,
            in3 => \N__27477\,
            lcout => \pwm_generator_inst.counter_i_3\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_2\,
            carryout => \pwm_generator_inst.un14_counter_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_8_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27297\,
            in2 => \N__27312\,
            in3 => \N__27522\,
            lcout => \pwm_generator_inst.counter_i_4\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_3\,
            carryout => \pwm_generator_inst.un14_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_8_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27426\,
            in1 => \N__27276\,
            in2 => \N__27291\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_5\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_4\,
            carryout => \pwm_generator_inst.un14_counter_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_8_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27450\,
            in1 => \N__27261\,
            in2 => \N__27270\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_6\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_5\,
            carryout => \pwm_generator_inst.un14_counter_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_8_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27588\,
            in1 => \N__27246\,
            in2 => \N__27255\,
            in3 => \_gnd_net_\,
            lcout => \pwm_generator_inst.counter_i_7\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_6\,
            carryout => \pwm_generator_inst.un14_counter_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_8_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27228\,
            in2 => \N__27237\,
            in3 => \N__27630\,
            lcout => \pwm_generator_inst.counter_i_8\,
            ltout => OPEN,
            carryin => \bfn_8_25_0_\,
            carryout => \pwm_generator_inst.un14_counter_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_8_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27210\,
            in2 => \N__27222\,
            in3 => \N__27609\,
            lcout => \pwm_generator_inst.counter_i_9\,
            ltout => OPEN,
            carryin => \pwm_generator_inst.un14_counter_cry_8\,
            carryout => \pwm_generator_inst.un14_counter_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.pwm_out_LC_8_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27204\,
            lcout => pwm_output_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49806\,
            ce => 'H',
            sr => \N__49446\
        );

    \pwm_generator_inst.counter_RNIVDL3_9_LC_8_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27625\,
            in1 => \N__27604\,
            in2 => \_gnd_net_\,
            in3 => \N__27586\,
            lcout => \pwm_generator_inst.un1_counterlto9_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNISQD2_0_LC_8_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27562\,
            in2 => \_gnd_net_\,
            in3 => \N__27538\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlto2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIBO26_1_LC_8_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__27520\,
            in1 => \N__27499\,
            in2 => \N__27480\,
            in3 => \N__27475\,
            lcout => OPEN,
            ltout => \pwm_generator_inst.un1_counterlt9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.counter_RNIFA6C_5_LC_8_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__27456\,
            in1 => \N__27449\,
            in2 => \N__27429\,
            in3 => \N__27425\,
            lcout => \pwm_generator_inst.un1_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_8_30_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__27363\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_clk_12mhz_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_1_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__32616\,
            in1 => \N__30000\,
            in2 => \N__27788\,
            in3 => \N__31232\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49955\,
            ce => 'H',
            sr => \N__49316\
        );

    \phase_controller_inst1.stoper_tr.target_time_13_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__30303\,
            in1 => \_gnd_net_\,
            in2 => \N__36721\,
            in3 => \N__30271\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => \N__31250\,
            sr => \N__49324\
        );

    \phase_controller_inst1.stoper_tr.target_time_6_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28437\,
            in1 => \N__36704\,
            in2 => \_gnd_net_\,
            in3 => \N__28395\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => \N__31250\,
            sr => \N__49324\
        );

    \phase_controller_inst1.stoper_tr.target_time_1_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__32639\,
            in1 => \_gnd_net_\,
            in2 => \N__36722\,
            in3 => \N__32691\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49954\,
            ce => \N__31250\,
            sr => \N__49324\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29718\,
            in2 => \N__27789\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_2_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31117\,
            in1 => \N__27761\,
            in2 => \_gnd_net_\,
            in3 => \N__27747\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_3_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31121\,
            in1 => \N__27743\,
            in2 => \N__29985\,
            in3 => \N__27729\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_4_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31118\,
            in1 => \N__27725\,
            in2 => \_gnd_net_\,
            in3 => \N__27711\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_5_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31122\,
            in1 => \N__27707\,
            in2 => \_gnd_net_\,
            in3 => \N__27693\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_6_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31119\,
            in1 => \N__27689\,
            in2 => \_gnd_net_\,
            in3 => \N__27675\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_7_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31123\,
            in1 => \N__27668\,
            in2 => \_gnd_net_\,
            in3 => \N__27654\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_8_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31120\,
            in1 => \N__27650\,
            in2 => \_gnd_net_\,
            in3 => \N__27633\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49952\,
            ce => 'H',
            sr => \N__49332\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_9_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31219\,
            in1 => \N__27929\,
            in2 => \_gnd_net_\,
            in3 => \N__27915\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_10_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31212\,
            in1 => \N__27911\,
            in2 => \_gnd_net_\,
            in3 => \N__27897\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_11_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31216\,
            in1 => \N__27893\,
            in2 => \_gnd_net_\,
            in3 => \N__27879\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_12_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31213\,
            in1 => \N__27875\,
            in2 => \_gnd_net_\,
            in3 => \N__27861\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_13_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31217\,
            in1 => \N__27854\,
            in2 => \_gnd_net_\,
            in3 => \N__27840\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_14_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31214\,
            in1 => \N__27833\,
            in2 => \_gnd_net_\,
            in3 => \N__27819\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_15_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31218\,
            in1 => \N__27815\,
            in2 => \_gnd_net_\,
            in3 => \N__27801\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_16_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31215\,
            in1 => \N__29939\,
            in2 => \_gnd_net_\,
            in3 => \N__27798\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49948\,
            ce => 'H',
            sr => \N__49341\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_17_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31224\,
            in1 => \N__29921\,
            in2 => \_gnd_net_\,
            in3 => \N__28113\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_18_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31228\,
            in1 => \N__28102\,
            in2 => \_gnd_net_\,
            in3 => \N__28080\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_19_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31225\,
            in1 => \N__28075\,
            in2 => \_gnd_net_\,
            in3 => \N__28053\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_20_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31229\,
            in1 => \N__28048\,
            in2 => \_gnd_net_\,
            in3 => \N__28032\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_21_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__31226\,
            in1 => \_gnd_net_\,
            in2 => \N__28028\,
            in3 => \N__28005\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_22_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31230\,
            in1 => \N__28002\,
            in2 => \_gnd_net_\,
            in3 => \N__27987\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_23_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31227\,
            in1 => \N__27984\,
            in2 => \_gnd_net_\,
            in3 => \N__27969\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_24_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31231\,
            in1 => \N__27966\,
            in2 => \_gnd_net_\,
            in3 => \N__27951\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49938\,
            ce => 'H',
            sr => \N__49350\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_25_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31233\,
            in1 => \N__27948\,
            in2 => \_gnd_net_\,
            in3 => \N__27933\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_26_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31237\,
            in1 => \N__28264\,
            in2 => \_gnd_net_\,
            in3 => \N__28248\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_27_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31234\,
            in1 => \N__28245\,
            in2 => \_gnd_net_\,
            in3 => \N__28230\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_28_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31238\,
            in1 => \N__28145\,
            in2 => \_gnd_net_\,
            in3 => \N__28227\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_29_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31235\,
            in1 => \N__28161\,
            in2 => \_gnd_net_\,
            in3 => \N__28224\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_30_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31239\,
            in1 => \N__28220\,
            in2 => \_gnd_net_\,
            in3 => \N__28200\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.accumulated_time_31_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31236\,
            in1 => \N__28193\,
            in2 => \_gnd_net_\,
            in3 => \N__28197\,
            lcout => \phase_controller_inst1.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49928\,
            ce => 'H',
            sr => \N__49359\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_28_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__28160\,
            in1 => \N__28141\,
            in2 => \N__28323\,
            in3 => \N__29874\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_28_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__29873\,
            in1 => \N__28159\,
            in2 => \N__28146\,
            in3 => \N__28319\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_29_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30769\,
            in1 => \N__30753\,
            in2 => \_gnd_net_\,
            in3 => \N__36682\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49916\,
            ce => \N__31264\,
            sr => \N__49366\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36413\,
            in1 => \N__30105\,
            in2 => \_gnd_net_\,
            in3 => \N__30083\,
            lcout => \elapsed_time_ns_1_RNIT6OBB_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30773\,
            in1 => \N__30752\,
            in2 => \_gnd_net_\,
            in3 => \N__36409\,
            lcout => \elapsed_time_ns_1_RNI7IPBB_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIH57P1_17_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__28768\,
            in1 => \N__31348\,
            in2 => \N__33204\,
            in3 => \N__36762\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII9257_13_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__28311\,
            in1 => \N__28305\,
            in2 => \N__28299\,
            in3 => \N__28296\,
            lcout => \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36412\,
            in1 => \N__28430\,
            in2 => \_gnd_net_\,
            in3 => \N__28393\,
            lcout => \elapsed_time_ns_1_RNIIH91B_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31000\,
            in1 => \N__30970\,
            in2 => \_gnd_net_\,
            in3 => \N__36410\,
            lcout => \elapsed_time_ns_1_RNIKJ91B_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33067\,
            in1 => \N__33026\,
            in2 => \_gnd_net_\,
            in3 => \N__36411\,
            lcout => \elapsed_time_ns_1_RNI6HPBB_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_24_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__31751\,
            in1 => \N__28280\,
            in2 => \N__31728\,
            in3 => \N__28572\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_24_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__28571\,
            in1 => \N__31727\,
            in2 => \N__28284\,
            in3 => \N__31752\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_24_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36467\,
            in1 => \N__28627\,
            in2 => \_gnd_net_\,
            in3 => \N__28609\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49893\,
            ce => \N__33335\,
            sr => \N__49376\
        );

    \phase_controller_inst2.stoper_tr.target_time_12_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28558\,
            in1 => \N__28536\,
            in2 => \_gnd_net_\,
            in3 => \N__36468\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49893\,
            ce => \N__33335\,
            sr => \N__49376\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_20_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001100"
        )
    port map (
            in0 => \N__31841\,
            in1 => \N__28811\,
            in2 => \N__31821\,
            in3 => \N__28446\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_20_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__28445\,
            in1 => \N__31820\,
            in2 => \N__28815\,
            in3 => \N__31842\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_2_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28509\,
            in1 => \N__28482\,
            in2 => \_gnd_net_\,
            in3 => \N__36473\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49880\,
            ce => \N__33337\,
            sr => \N__49381\
        );

    \phase_controller_inst2.stoper_tr.target_time_20_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33155\,
            in1 => \N__33201\,
            in2 => \_gnd_net_\,
            in3 => \N__36560\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => \N__33340\,
            sr => \N__49386\
        );

    \phase_controller_inst2.stoper_tr.target_time_6_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36672\,
            in1 => \N__28422\,
            in2 => \_gnd_net_\,
            in3 => \N__28394\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => \N__33340\,
            sr => \N__49386\
        );

    \phase_controller_inst2.stoper_tr.target_time_4_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28364\,
            in1 => \N__28339\,
            in2 => \_gnd_net_\,
            in3 => \N__36561\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => \N__33340\,
            sr => \N__49386\
        );

    \phase_controller_inst2.stoper_tr.target_time_18_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31314\,
            in1 => \N__31338\,
            in2 => \_gnd_net_\,
            in3 => \N__36559\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49870\,
            ce => \N__33340\,
            sr => \N__49386\
        );

    \phase_controller_inst2.stoper_tr.target_time_31_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__28973\,
            in1 => \N__28938\,
            in2 => \_gnd_net_\,
            in3 => \N__36558\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => \N__33341\,
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.target_time_27_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36555\,
            in1 => \N__28909\,
            in2 => \_gnd_net_\,
            in3 => \N__28884\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => \N__33341\,
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.target_time_21_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28866\,
            in1 => \N__28834\,
            in2 => \_gnd_net_\,
            in3 => \N__36557\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => \N__33341\,
            sr => \N__49390\
        );

    \phase_controller_inst2.stoper_tr.target_time_19_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__28800\,
            in1 => \N__28758\,
            in2 => \_gnd_net_\,
            in3 => \N__36556\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49860\,
            ce => \N__33341\,
            sr => \N__49390\
        );

    \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31899\,
            in1 => \N__28740\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axb_0\,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32127\,
            in2 => \_gnd_net_\,
            in3 => \N__28698\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_0\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32115\,
            in3 => \N__28668\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_1\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_3_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32100\,
            in2 => \_gnd_net_\,
            in3 => \N__28635\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_2\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_4_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32088\,
            in2 => \_gnd_net_\,
            in3 => \N__29217\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_3\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_5_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32076\,
            in3 => \N__29196\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_4\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_6_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32061\,
            in2 => \_gnd_net_\,
            in3 => \N__29172\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_5\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32049\,
            in3 => \N__29142\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_6\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_7\,
            clk => \N__49847\,
            ce => 'H',
            sr => \N__49395\
        );

    \current_shift_inst.PI_CTRL.error_control_8_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32034\,
            in3 => \N__29109\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_8\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_9_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32019\,
            in2 => \_gnd_net_\,
            in3 => \N__29079\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_8\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_10_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32235\,
            in3 => \N__29046\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_9\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_11_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32220\,
            in2 => \_gnd_net_\,
            in3 => \N__29013\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_10\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_12_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32208\,
            in2 => \_gnd_net_\,
            in3 => \N__28977\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_11\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_13_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32196\,
            in3 => \N__29448\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_12\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_14_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32181\,
            in2 => \_gnd_net_\,
            in3 => \N__29418\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_13\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_15_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32169\,
            in3 => \N__29394\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_14\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_15\,
            clk => \N__49837\,
            ce => 'H',
            sr => \N__49398\
        );

    \current_shift_inst.PI_CTRL.error_control_16_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32154\,
            in2 => \_gnd_net_\,
            in3 => \N__29361\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_16\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_17_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32142\,
            in3 => \N__29337\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_16\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_18_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32340\,
            in2 => \_gnd_net_\,
            in3 => \N__29307\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_17\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_19_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32328\,
            in2 => \_gnd_net_\,
            in3 => \N__29274\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_18\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_20_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32316\,
            in3 => \N__29247\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_19\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_21_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32301\,
            in2 => \_gnd_net_\,
            in3 => \N__29688\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_20\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_22_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32289\,
            in3 => \N__29658\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_21\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_23_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32274\,
            in3 => \N__29631\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_22\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_23\,
            clk => \N__49828\,
            ce => 'H',
            sr => \N__49403\
        );

    \current_shift_inst.PI_CTRL.error_control_24_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32259\,
            in2 => \_gnd_net_\,
            in3 => \N__29601\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_24\,
            ltout => OPEN,
            carryin => \bfn_9_16_0_\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_25_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32247\,
            in2 => \_gnd_net_\,
            in3 => \N__29568\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_24\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_26_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32448\,
            in2 => \_gnd_net_\,
            in3 => \N__29535\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_25\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_27_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32436\,
            in2 => \_gnd_net_\,
            in3 => \N__29502\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_26\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_28_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32424\,
            in3 => \N__29472\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_27\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_29_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32409\,
            in3 => \N__29841\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_28\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_30_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30717\,
            in2 => \_gnd_net_\,
            in3 => \N__29811\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.PI_CTRL.error_control_2_cry_29\,
            carryout => \current_shift_inst.PI_CTRL.error_control_2_cry_30\,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.error_control_31_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32391\,
            in2 => \_gnd_net_\,
            in3 => \N__29808\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49822\,
            ce => 'H',
            sr => \N__49408\
        );

    \current_shift_inst.PI_CTRL.prop_term_31_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29805\,
            lcout => \current_shift_inst.PI_CTRL.prop_termZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49814\,
            ce => 'H',
            sr => \N__49426\
        );

    \current_shift_inst.PI_CTRL.control_out_10_LC_9_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29787\,
            lcout => \N_19_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49808\,
            ce => 'H',
            sr => \N__49437\
        );

    \phase_controller_inst1.stoper_tr.target_time_3_LC_10_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31376\,
            in1 => \N__31419\,
            in2 => \_gnd_net_\,
            in3 => \N__36702\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49953\,
            ce => \N__31256\,
            sr => \N__49302\
        );

    \phase_controller_inst1.stoper_tr.running_LC_10_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010011101110"
        )
    port map (
            in0 => \N__32605\,
            in1 => \N__31431\,
            in2 => \N__32583\,
            in3 => \N__32535\,
            lcout => \phase_controller_inst1.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49939\,
            ce => 'H',
            sr => \N__49317\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI3C8N_30_LC_10_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32534\,
            in2 => \_gnd_net_\,
            in3 => \N__32575\,
            lcout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29721\,
            in3 => \N__32603\,
            lcout => \phase_controller_inst1.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1_30_LC_10_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29996\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNI9P8V1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_9_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30121\,
            in1 => \N__30162\,
            in2 => \_gnd_net_\,
            in3 => \N__36712\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49929\,
            ce => \N__31199\,
            sr => \N__49325\
        );

    \phase_controller_inst1.stoper_tr.target_time_16_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32506\,
            in1 => \N__32486\,
            in2 => \_gnd_net_\,
            in3 => \N__36711\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49929\,
            ce => \N__31199\,
            sr => \N__49325\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0_16_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__29917\,
            in1 => \N__29886\,
            in2 => \N__29940\,
            in3 => \N__29949\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_16_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__29948\,
            in1 => \N__29938\,
            in2 => \N__29922\,
            in3 => \N__29885\,
            lcout => \phase_controller_inst1.stoper_tr.un4_running_cry_c_RNO_0Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36631\,
            in1 => \N__30125\,
            in2 => \_gnd_net_\,
            in3 => \N__30154\,
            lcout => \elapsed_time_ns_1_RNILK91B_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30298\,
            in1 => \N__36630\,
            in2 => \_gnd_net_\,
            in3 => \N__30278\,
            lcout => \elapsed_time_ns_1_RNI0AOBB_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_17_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36237\,
            in1 => \N__36773\,
            in2 => \_gnd_net_\,
            in3 => \N__36679\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49906\,
            ce => \N__31266\,
            sr => \N__49342\
        );

    \phase_controller_inst1.stoper_tr.target_time_28_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33072\,
            in1 => \N__33022\,
            in2 => \_gnd_net_\,
            in3 => \N__36680\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49906\,
            ce => \N__31266\,
            sr => \N__49342\
        );

    \phase_controller_inst2.stoper_tr.target_time_13_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36673\,
            in1 => \N__30299\,
            in2 => \_gnd_net_\,
            in3 => \N__30279\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => \N__33333\,
            sr => \N__49351\
        );

    \phase_controller_inst2.stoper_tr.target_time_5_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30227\,
            in1 => \N__30189\,
            in2 => \_gnd_net_\,
            in3 => \N__36677\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => \N__33333\,
            sr => \N__49351\
        );

    \phase_controller_inst2.stoper_tr.target_time_1_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36674\,
            in1 => \N__32646\,
            in2 => \_gnd_net_\,
            in3 => \N__32683\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => \N__33333\,
            sr => \N__49351\
        );

    \phase_controller_inst2.stoper_tr.target_time_9_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30161\,
            in1 => \N__30126\,
            in2 => \_gnd_net_\,
            in3 => \N__36678\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => \N__33333\,
            sr => \N__49351\
        );

    \phase_controller_inst2.stoper_tr.target_time_3_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36675\,
            in1 => \N__31380\,
            in2 => \_gnd_net_\,
            in3 => \N__31418\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => \N__33333\,
            sr => \N__49351\
        );

    \phase_controller_inst2.stoper_tr.target_time_10_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30104\,
            in1 => \N__30087\,
            in2 => \_gnd_net_\,
            in3 => \N__36676\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49895\,
            ce => \N__33333\,
            sr => \N__49351\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_1_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30039\,
            in2 => \N__30048\,
            in3 => \N__32770\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_10_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_2_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30021\,
            in2 => \N__30033\,
            in3 => \N__31535\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30006\,
            in2 => \N__30015\,
            in3 => \N__31520\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_4_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30441\,
            in2 => \N__30432\,
            in3 => \N__31505\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_5_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30423\,
            in2 => \N__30417\,
            in3 => \N__31490\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_6_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30405\,
            in2 => \N__30396\,
            in3 => \N__31475\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_7_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30387\,
            in2 => \N__30375\,
            in3 => \N__31460\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_8_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31445\,
            in1 => \N__30945\,
            in2 => \N__30366\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_9_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30357\,
            in2 => \N__30348\,
            in3 => \N__31700\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_10_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30339\,
            in2 => \N__30330\,
            in3 => \N__31685\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_11_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30321\,
            in2 => \N__30312\,
            in3 => \N__31670\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_12_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30534\,
            in2 => \N__30543\,
            in3 => \N__31655\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_13_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31640\,
            in1 => \N__30528\,
            in2 => \N__30519\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_14_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30510\,
            in2 => \N__31548\,
            in3 => \N__31625\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_inv_15_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30504\,
            in2 => \N__30489\,
            in3 => \N__31610\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_16_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33099\,
            in2 => \N__32940\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_18_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30816\,
            in2 => \N__30849\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_20_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30480\,
            in2 => \N__30474\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_22_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30462\,
            in2 => \N__30453\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_24_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30678\,
            in2 => \N__30672\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_26_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30639\,
            in2 => \N__30660\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_28_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33222\,
            in2 => \N__33087\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_30_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30927\,
            in2 => \N__30552\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_LUT4_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30663\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_26_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__32005\,
            in1 => \N__31988\,
            in2 => \N__30651\,
            in3 => \N__30561\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_26_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__30560\,
            in1 => \N__32006\,
            in2 => \N__31989\,
            in3 => \N__30650\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_26_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30633\,
            in1 => \N__30604\,
            in2 => \_gnd_net_\,
            in3 => \N__36671\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49849\,
            ce => \N__33336\,
            sr => \N__49377\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_30_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__30857\,
            in1 => \N__31934\,
            in2 => \N__30939\,
            in3 => \N__31957\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_30_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101100100010"
        )
    port map (
            in0 => \N__31933\,
            in1 => \N__30938\,
            in2 => \N__31959\,
            in3 => \N__30858\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_30_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__36670\,
            in1 => \N__30921\,
            in2 => \_gnd_net_\,
            in3 => \N__30894\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49849\,
            ce => \N__33336\,
            sr => \N__49377\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_18_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110101000100"
        )
    port map (
            in0 => \N__31862\,
            in1 => \N__30824\,
            in2 => \N__31887\,
            in3 => \N__30837\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_18_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__30836\,
            in1 => \N__31886\,
            in2 => \N__30828\,
            in3 => \N__31863\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_0_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31919\,
            in2 => \_gnd_net_\,
            in3 => \N__37830\,
            lcout => \current_shift_inst.PI_CTRL.prop_term_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49830\,
            ce => 'H',
            sr => \N__49387\
        );

    \phase_controller_inst2.stoper_tr.target_time_29_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30777\,
            in1 => \N__30751\,
            in2 => \_gnd_net_\,
            in3 => \N__36714\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49823\,
            ce => \N__33342\,
            sr => \N__49391\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32387\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_16_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__48891\,
            in1 => \N__30711\,
            in2 => \N__48729\,
            in3 => \N__48932\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__32526\,
            in1 => \N__31430\,
            in2 => \_gnd_net_\,
            in3 => \N__32550\,
            lcout => \phase_controller_inst1.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.start_latched_RNI59OS_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__32551\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32527\,
            lcout => \phase_controller_inst1.stoper_tr.start_latched_RNI59OSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31375\,
            in1 => \N__31414\,
            in2 => \_gnd_net_\,
            in3 => \N__36687\,
            lcout => \elapsed_time_ns_1_RNIFE91B_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32508\,
            in1 => \N__32485\,
            in2 => \_gnd_net_\,
            in3 => \N__36688\,
            lcout => \elapsed_time_ns_1_RNI3DOBB_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.start_timer_tr_RNO_0_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__32887\,
            in1 => \N__33724\,
            in2 => \N__38322\,
            in3 => \N__32847\,
            lcout => \phase_controller_inst2.N_54_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31306\,
            in1 => \N__31355\,
            in2 => \_gnd_net_\,
            in3 => \N__36689\,
            lcout => \elapsed_time_ns_1_RNI5FOBB_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31591\,
            in1 => \N__31559\,
            in2 => \_gnd_net_\,
            in3 => \N__36690\,
            lcout => \elapsed_time_ns_1_RNI1BOBB_0_14\,
            ltout => \elapsed_time_ns_1_RNI1BOBB_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.target_time_14_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__36691\,
            in1 => \_gnd_net_\,
            in2 => \N__31284\,
            in3 => \N__31592\,
            lcout => \phase_controller_inst1.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49896\,
            ce => \N__31263\,
            sr => \N__49333\
        );

    \phase_controller_inst2.stoper_tr.target_time_8_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__31005\,
            in1 => \N__30978\,
            in2 => \_gnd_net_\,
            in3 => \N__36701\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => \N__33332\,
            sr => \N__49343\
        );

    \phase_controller_inst2.stoper_tr.target_time_14_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31593\,
            in1 => \N__31560\,
            in2 => \_gnd_net_\,
            in3 => \N__36700\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49881\,
            ce => \N__33332\,
            sr => \N__49343\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32709\,
            in2 => \N__32771\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33668\,
            in1 => \N__31536\,
            in2 => \_gnd_net_\,
            in3 => \N__31524\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_3_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__33676\,
            in1 => \N__31521\,
            in2 => \N__33132\,
            in3 => \N__31509\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_4_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33669\,
            in1 => \N__31506\,
            in2 => \_gnd_net_\,
            in3 => \N__31494\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_5_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33677\,
            in1 => \N__31491\,
            in2 => \_gnd_net_\,
            in3 => \N__31479\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_6_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33670\,
            in1 => \N__31476\,
            in2 => \_gnd_net_\,
            in3 => \N__31464\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_7_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33678\,
            in1 => \N__31461\,
            in2 => \_gnd_net_\,
            in3 => \N__31449\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_8_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33671\,
            in1 => \N__31446\,
            in2 => \_gnd_net_\,
            in3 => \N__31434\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_7\,
            clk => \N__49872\,
            ce => 'H',
            sr => \N__49352\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_9_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33675\,
            in1 => \N__31701\,
            in2 => \_gnd_net_\,
            in3 => \N__31689\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_10_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33679\,
            in1 => \N__31686\,
            in2 => \_gnd_net_\,
            in3 => \N__31674\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_11_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33672\,
            in1 => \N__31671\,
            in2 => \_gnd_net_\,
            in3 => \N__31659\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_12_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33680\,
            in1 => \N__31656\,
            in2 => \_gnd_net_\,
            in3 => \N__31644\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_13_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33673\,
            in1 => \N__31641\,
            in2 => \_gnd_net_\,
            in3 => \N__31629\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_14_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33681\,
            in1 => \N__31626\,
            in2 => \_gnd_net_\,
            in3 => \N__31614\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_15_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33674\,
            in1 => \N__31611\,
            in2 => \_gnd_net_\,
            in3 => \N__31599\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_16_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33682\,
            in1 => \N__32962\,
            in2 => \_gnd_net_\,
            in3 => \N__31596\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_15\,
            clk => \N__49862\,
            ce => 'H',
            sr => \N__49360\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_17_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33692\,
            in1 => \N__33000\,
            in2 => \_gnd_net_\,
            in3 => \N__31890\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_18_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33696\,
            in1 => \N__31882\,
            in2 => \_gnd_net_\,
            in3 => \N__31866\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_19_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33693\,
            in1 => \N__31861\,
            in2 => \_gnd_net_\,
            in3 => \N__31845\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_20_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33697\,
            in1 => \N__31840\,
            in2 => \_gnd_net_\,
            in3 => \N__31824\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_21_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33694\,
            in1 => \N__31816\,
            in2 => \_gnd_net_\,
            in3 => \N__31800\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_22_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33698\,
            in1 => \N__31792\,
            in2 => \_gnd_net_\,
            in3 => \N__31776\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_23_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33695\,
            in1 => \N__31771\,
            in2 => \_gnd_net_\,
            in3 => \N__31755\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_24_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33699\,
            in1 => \N__31745\,
            in2 => \_gnd_net_\,
            in3 => \N__31731\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_23\,
            clk => \N__49850\,
            ce => 'H',
            sr => \N__49367\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_25_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33689\,
            in1 => \N__31718\,
            in2 => \_gnd_net_\,
            in3 => \N__31704\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_26_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33685\,
            in1 => \N__32007\,
            in2 => \_gnd_net_\,
            in3 => \N__31992\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_27_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33690\,
            in1 => \N__31984\,
            in2 => \_gnd_net_\,
            in3 => \N__31968\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_28_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33686\,
            in1 => \N__33240\,
            in2 => \_gnd_net_\,
            in3 => \N__31965\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_29_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33691\,
            in1 => \N__33282\,
            in2 => \_gnd_net_\,
            in3 => \N__31962\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_30_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__33687\,
            in1 => \N__31958\,
            in2 => \_gnd_net_\,
            in3 => \N__31941\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_29\,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_31_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__31935\,
            in1 => \N__33688\,
            in2 => \_gnd_net_\,
            in3 => \N__31938\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49839\,
            ce => 'H',
            sr => \N__49372\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38489\,
            lcout => \current_shift_inst.N_1263_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37829\,
            in2 => \N__31920\,
            in3 => \N__31918\,
            lcout => \current_shift_inst.control_input_1\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \current_shift_inst.control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37353\,
            in2 => \_gnd_net_\,
            in3 => \N__32118\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_0\,
            carryout => \current_shift_inst.control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33300\,
            in2 => \_gnd_net_\,
            in3 => \N__32103\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_1\,
            carryout => \current_shift_inst.control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38022\,
            in2 => \_gnd_net_\,
            in3 => \N__32091\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_2\,
            carryout => \current_shift_inst.control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38145\,
            in2 => \_gnd_net_\,
            in3 => \N__32079\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_3\,
            carryout => \current_shift_inst.control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37860\,
            in2 => \_gnd_net_\,
            in3 => \N__32064\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_4\,
            carryout => \current_shift_inst.control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33210\,
            in2 => \_gnd_net_\,
            in3 => \N__32052\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_5\,
            carryout => \current_shift_inst.control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38100\,
            in2 => \_gnd_net_\,
            in3 => \N__32037\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_6\,
            carryout => \current_shift_inst.control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38052\,
            in2 => \_gnd_net_\,
            in3 => \N__32022\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \current_shift_inst.control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33384\,
            in2 => \_gnd_net_\,
            in3 => \N__32010\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_8\,
            carryout => \current_shift_inst.control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33411\,
            in2 => \_gnd_net_\,
            in3 => \N__32223\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_9\,
            carryout => \current_shift_inst.control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33366\,
            in2 => \_gnd_net_\,
            in3 => \N__32211\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_10\,
            carryout => \current_shift_inst.control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33378\,
            in2 => \_gnd_net_\,
            in3 => \N__32199\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_11\,
            carryout => \current_shift_inst.control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33372\,
            in2 => \_gnd_net_\,
            in3 => \N__32184\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_12\,
            carryout => \current_shift_inst.control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33441\,
            in2 => \_gnd_net_\,
            in3 => \N__32172\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_13\,
            carryout => \current_shift_inst.control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33360\,
            in2 => \_gnd_net_\,
            in3 => \N__32157\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_14\,
            carryout => \current_shift_inst.control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33435\,
            in2 => \_gnd_net_\,
            in3 => \N__32145\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \current_shift_inst.control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32364\,
            in2 => \_gnd_net_\,
            in3 => \N__32130\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_16\,
            carryout => \current_shift_inst.control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33429\,
            in2 => \_gnd_net_\,
            in3 => \N__32331\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_17\,
            carryout => \current_shift_inst.control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33423\,
            in2 => \_gnd_net_\,
            in3 => \N__32319\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_18\,
            carryout => \current_shift_inst.control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33417\,
            in2 => \_gnd_net_\,
            in3 => \N__32304\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_19\,
            carryout => \current_shift_inst.control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36807\,
            in2 => \_gnd_net_\,
            in3 => \N__32292\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_20\,
            carryout => \current_shift_inst.control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36105\,
            in2 => \_gnd_net_\,
            in3 => \N__32277\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_21\,
            carryout => \current_shift_inst.control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33402\,
            in2 => \_gnd_net_\,
            in3 => \N__32262\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_22\,
            carryout => \current_shift_inst.control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33396\,
            in2 => \_gnd_net_\,
            in3 => \N__32250\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_11_16_0_\,
            carryout => \current_shift_inst.control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33390\,
            in2 => \_gnd_net_\,
            in3 => \N__32238\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_24\,
            carryout => \current_shift_inst.control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32376\,
            in2 => \_gnd_net_\,
            in3 => \N__32439\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_25\,
            carryout => \current_shift_inst.control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33549\,
            in2 => \_gnd_net_\,
            in3 => \N__32427\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_26\,
            carryout => \current_shift_inst.control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36048\,
            in2 => \_gnd_net_\,
            in3 => \N__32412\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_27\,
            carryout => \current_shift_inst.control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32370\,
            in2 => \_gnd_net_\,
            in3 => \N__32397\,
            lcout => \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.control_input_cry_28\,
            carryout => \current_shift_inst.control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38496\,
            in2 => \_gnd_net_\,
            in3 => \N__32394\,
            lcout => \current_shift_inst.control_input_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34659\,
            in1 => \N__36093\,
            in2 => \_gnd_net_\,
            in3 => \N__38497\,
            lcout => \current_shift_inst.control_input_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38498\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34566\,
            in1 => \N__35799\,
            in2 => \_gnd_net_\,
            in3 => \N__38479\,
            lcout => \current_shift_inst.control_input_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.S2_LC_11_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32865\,
            lcout => s4_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49799\,
            ce => 'H',
            sr => \N__49434\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32638\,
            in1 => \N__32684\,
            in2 => \_gnd_net_\,
            in3 => \N__36686\,
            lcout => \elapsed_time_ns_1_RNIDC91B_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_RNO_0_3_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__33469\,
            in1 => \N__33802\,
            in2 => \N__33498\,
            in3 => \N__34887\,
            lcout => \phase_controller_inst1.state_ns_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_tr.time_passed_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000110010101100"
        )
    port map (
            in0 => \N__32533\,
            in1 => \N__33496\,
            in2 => \N__32615\,
            in3 => \N__32582\,
            lcout => \phase_controller_inst1.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49303\
        );

    \phase_controller_inst1.start_timer_tr_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001111110011"
        )
    port map (
            in0 => \N__33495\,
            in1 => \N__33840\,
            in2 => \N__32556\,
            in3 => \N__33473\,
            lcout => \phase_controller_inst1.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49303\
        );

    \phase_controller_inst1.stoper_tr.start_latched_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32555\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49917\,
            ce => 'H',
            sr => \N__49303\
        );

    \phase_controller_inst2.stoper_tr.target_time_16_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32507\,
            in1 => \N__32490\,
            in2 => \_gnd_net_\,
            in3 => \N__36713\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49905\,
            ce => \N__33331\,
            sr => \N__49310\
        );

    \phase_controller_inst2.start_timer_hc_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__33748\,
            in1 => \N__33707\,
            in2 => \N__38979\,
            in3 => \N__32914\,
            lcout => \phase_controller_inst2.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49894\,
            ce => 'H',
            sr => \N__49318\
        );

    \phase_controller_inst2.state_2_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101000110000"
        )
    port map (
            in0 => \N__32915\,
            in1 => \N__38321\,
            in2 => \N__33729\,
            in3 => \N__33749\,
            lcout => \phase_controller_inst2.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49894\,
            ce => 'H',
            sr => \N__49318\
        );

    \phase_controller_inst2.state_1_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__32854\,
            in1 => \N__33708\,
            in2 => \_gnd_net_\,
            in3 => \N__32888\,
            lcout => \phase_controller_inst2.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49894\,
            ce => 'H',
            sr => \N__49318\
        );

    \phase_controller_inst2.state_RNO_0_3_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__32922\,
            in1 => \N__33747\,
            in2 => \N__32802\,
            in3 => \N__32827\,
            lcout => \phase_controller_inst2.state_ns_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.state_0_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__32895\,
            in1 => \N__32828\,
            in2 => \N__32801\,
            in3 => \N__32858\,
            lcout => \phase_controller_inst2.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49871\,
            ce => 'H',
            sr => \N__49334\
        );

    \phase_controller_inst2.stoper_tr.time_passed_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000101011001100"
        )
    port map (
            in0 => \N__35710\,
            in1 => \N__32796\,
            in2 => \N__32745\,
            in3 => \N__35622\,
            lcout => \phase_controller_inst2.tr_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \N__49344\
        );

    \phase_controller_inst2.start_timer_tr_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111001111110011"
        )
    port map (
            in0 => \N__32829\,
            in1 => \N__32811\,
            in2 => \N__35656\,
            in3 => \N__32797\,
            lcout => \phase_controller_inst2.start_timer_trZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \N__49344\
        );

    \phase_controller_inst2.stoper_tr.accumulated_time_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__32703\,
            in1 => \N__35621\,
            in2 => \N__32772\,
            in3 => \N__33683\,
            lcout => \phase_controller_inst2.stoper_tr.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49861\,
            ce => 'H',
            sr => \N__49344\
        );

    \phase_controller_inst2.stoper_tr.running_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010111001100"
        )
    port map (
            in0 => \N__35706\,
            in1 => \N__35678\,
            in2 => \N__32744\,
            in3 => \N__35620\,
            lcout => \phase_controller_inst2.stoper_tr.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \N__49353\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNI54EN_30_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35705\,
            in2 => \_gnd_net_\,
            in3 => \N__32737\,
            lcout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_tr.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32712\,
            in3 => \N__35618\,
            lcout => \phase_controller_inst2.stoper_tr.un1_accumulated_time_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35660\,
            lcout => \phase_controller_inst2.stoper_tr.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49848\,
            ce => 'H',
            sr => \N__49353\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1_30_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35619\,
            in2 => \_gnd_net_\,
            in3 => \N__32702\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNIEA6F1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_28_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000100110000"
        )
    port map (
            in0 => \N__40847\,
            in1 => \N__40823\,
            in2 => \N__33111\,
            in3 => \N__33120\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_28_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__33119\,
            in1 => \N__40848\,
            in2 => \N__40827\,
            in3 => \N__33107\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_28_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39696\,
            in1 => \N__34269\,
            in2 => \_gnd_net_\,
            in3 => \N__47075\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49838\,
            ce => \N__47153\,
            sr => \N__49361\
        );

    \phase_controller_inst2.stoper_hc.target_time_29_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47074\,
            in1 => \N__39654\,
            in2 => \_gnd_net_\,
            in3 => \N__34250\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49838\,
            ce => \N__47153\,
            sr => \N__49361\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__37241\,
            in1 => \N__41120\,
            in2 => \N__41319\,
            in3 => \N__37220\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_16_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000100"
        )
    port map (
            in0 => \N__32999\,
            in1 => \N__32982\,
            in2 => \N__32966\,
            in3 => \N__33354\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_28_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__33293\,
            in1 => \N__33280\,
            in2 => \N__33263\,
            in3 => \N__33238\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_28_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__33068\,
            in1 => \N__33027\,
            in2 => \_gnd_net_\,
            in3 => \N__36720\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49829\,
            ce => \N__33334\,
            sr => \N__49368\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_16_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101000101"
        )
    port map (
            in0 => \N__32998\,
            in1 => \N__32981\,
            in2 => \N__32967\,
            in3 => \N__33353\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.target_time_17_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36230\,
            in1 => \N__36763\,
            in2 => \_gnd_net_\,
            in3 => \N__36719\,
            lcout => \phase_controller_inst2.stoper_tr.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49829\,
            ce => \N__33334\,
            sr => \N__49368\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34383\,
            in1 => \N__35778\,
            in2 => \_gnd_net_\,
            in3 => \N__38490\,
            lcout => \current_shift_inst.control_input_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.un4_running_cry_c_RNO_0_28_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__33294\,
            in1 => \N__33281\,
            in2 => \N__33264\,
            in3 => \N__33239\,
            lcout => \phase_controller_inst2.stoper_tr.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34512\,
            in1 => \N__35754\,
            in2 => \_gnd_net_\,
            in3 => \N__38491\,
            lcout => \current_shift_inst.control_input_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33148\,
            in1 => \N__33202\,
            in2 => \_gnd_net_\,
            in3 => \N__36718\,
            lcout => \elapsed_time_ns_1_RNIU8PBB_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_8_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46913\,
            in1 => \N__37901\,
            in2 => \_gnd_net_\,
            in3 => \N__39273\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49819\,
            ce => \N__47152\,
            sr => \N__49378\
        );

    \phase_controller_inst2.stoper_hc.target_time_30_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39612\,
            in1 => \N__34345\,
            in2 => \_gnd_net_\,
            in3 => \N__46914\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49819\,
            ce => \N__47152\,
            sr => \N__49378\
        );

    \phase_controller_inst2.stoper_hc.target_time_31_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39567\,
            in1 => \N__34453\,
            in2 => \_gnd_net_\,
            in3 => \N__46915\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49819\,
            ce => \N__47152\,
            sr => \N__49378\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34347\,
            in1 => \N__39611\,
            in2 => \_gnd_net_\,
            in3 => \N__46722\,
            lcout => \elapsed_time_ns_1_RNIV2EN9_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_30_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001110"
        )
    port map (
            in0 => \N__34430\,
            in1 => \N__35478\,
            in2 => \N__35520\,
            in3 => \N__34416\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_8_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46723\,
            in1 => \N__37905\,
            in2 => \_gnd_net_\,
            in3 => \N__39272\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49817\,
            ce => \N__37638\,
            sr => \N__49382\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35910\,
            in1 => \N__34491\,
            in2 => \_gnd_net_\,
            in3 => \N__38460\,
            lcout => \current_shift_inst.control_input_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46830\,
            in1 => \N__34246\,
            in2 => \_gnd_net_\,
            in3 => \N__39653\,
            lcout => \elapsed_time_ns_1_RNI7ADN9_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__34455\,
            in1 => \N__39563\,
            in2 => \_gnd_net_\,
            in3 => \N__46831\,
            lcout => \elapsed_time_ns_1_RNI04EN9_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38462\,
            in1 => \N__35865\,
            in2 => \_gnd_net_\,
            in3 => \N__34626\,
            lcout => \current_shift_inst.control_input_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35850\,
            in1 => \N__34614\,
            in2 => \_gnd_net_\,
            in3 => \N__38463\,
            lcout => \current_shift_inst.control_input_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38461\,
            in1 => \N__34470\,
            in2 => \_gnd_net_\,
            in3 => \N__35880\,
            lcout => \current_shift_inst.control_input_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34590\,
            in1 => \N__35826\,
            in2 => \_gnd_net_\,
            in3 => \N__38467\,
            lcout => \current_shift_inst.control_input_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110101"
        )
    port map (
            in0 => \N__34602\,
            in1 => \_gnd_net_\,
            in2 => \N__38492\,
            in3 => \N__35838\,
            lcout => \current_shift_inst.control_input_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38493\,
            in1 => \N__35814\,
            in2 => \_gnd_net_\,
            in3 => \N__34578\,
            lcout => \current_shift_inst.control_input_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38455\,
            in1 => \N__36000\,
            in2 => \_gnd_net_\,
            in3 => \N__34554\,
            lcout => \current_shift_inst.control_input_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34542\,
            in1 => \N__35985\,
            in2 => \_gnd_net_\,
            in3 => \N__38456\,
            lcout => \current_shift_inst.control_input_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38457\,
            in1 => \N__34530\,
            in2 => \_gnd_net_\,
            in3 => \N__35970\,
            lcout => \current_shift_inst.control_input_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__35895\,
            in1 => \N__34479\,
            in2 => \_gnd_net_\,
            in3 => \N__38454\,
            lcout => \current_shift_inst.control_input_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34695\,
            in1 => \N__35949\,
            in2 => \_gnd_net_\,
            in3 => \N__38458\,
            lcout => \current_shift_inst.control_input_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38459\,
            in1 => \N__34683\,
            in2 => \_gnd_net_\,
            in3 => \N__35937\,
            lcout => \current_shift_inst.control_input_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__34671\,
            in1 => \N__35925\,
            in2 => \_gnd_net_\,
            in3 => \N__38494\,
            lcout => \current_shift_inst.control_input_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38495\,
            in1 => \N__34644\,
            in2 => \_gnd_net_\,
            in3 => \N__36078\,
            lcout => \current_shift_inst.control_input_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.stop_timer_hc_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49991\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.stop_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33543\,
            ce => 'H',
            sr => \N__49404\
        );

    \delay_measurement_inst.start_timer_hc_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49990\,
            lcout => \delay_measurement_inst.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33543\,
            ce => 'H',
            sr => \N__49404\
        );

    \phase_controller_inst2.S1_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33759\,
            lcout => s3_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49802\,
            ce => 'H',
            sr => \N__49411\
        );

    \GB_BUFFER_red_c_g_THRU_LUT4_0_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__49476\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_red_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_3_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100011111111"
        )
    port map (
            in0 => \N__35083\,
            in1 => \N__33452\,
            in2 => \N__33875\,
            in3 => \N__33504\,
            lcout => state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => 'H',
            sr => \N__49291\
        );

    \phase_controller_inst1.state_2_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__33809\,
            in1 => \N__33834\,
            in2 => \N__34910\,
            in3 => \N__33857\,
            lcout => \phase_controller_inst1.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => 'H',
            sr => \N__49291\
        );

    \phase_controller_inst1.state_0_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__34777\,
            in1 => \N__34727\,
            in2 => \N__33474\,
            in3 => \N__33497\,
            lcout => \phase_controller_inst1.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => 'H',
            sr => \N__49291\
        );

    \phase_controller_inst1.state_4_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__33453\,
            in1 => \N__33868\,
            in2 => \_gnd_net_\,
            in3 => \N__35084\,
            lcout => \phase_controller_inst1.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => 'H',
            sr => \N__49291\
        );

    \phase_controller_inst1.start_flag_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__35082\,
            in1 => \N__33451\,
            in2 => \N__33876\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49940\,
            ce => 'H',
            sr => \N__49291\
        );

    \phase_controller_inst1.state_RNIE87F_2_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__33856\,
            in1 => \N__33828\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__34778\,
            in1 => \N__33829\,
            in2 => \N__33858\,
            in3 => \N__34722\,
            lcout => \phase_controller_inst1.N_54_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36979\,
            lcout => \phase_controller_inst1.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49304\
        );

    \phase_controller_inst1.stoper_hc.time_passed_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__33833\,
            in1 => \N__33948\,
            in2 => \N__37014\,
            in3 => \N__34142\,
            lcout => \phase_controller_inst1.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49304\
        );

    \phase_controller_inst1.start_timer_hc_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__33810\,
            in1 => \N__34745\,
            in2 => \N__34916\,
            in3 => \N__36978\,
            lcout => \phase_controller_inst1.start_timer_hcZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49918\,
            ce => 'H',
            sr => \N__49304\
        );

    \phase_controller_inst2.state_3_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__35087\,
            in1 => \N__35021\,
            in2 => \N__33768\,
            in3 => \N__35037\,
            lcout => \phase_controller_inst2.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49907\,
            ce => 'H',
            sr => \N__49311\
        );

    \phase_controller_inst2.state_RNIG7JF_2_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38320\,
            in2 => \_gnd_net_\,
            in3 => \N__33725\,
            lcout => \phase_controller_inst2.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.start_latched_RNI7GMN_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35718\,
            in2 => \_gnd_net_\,
            in3 => \N__35655\,
            lcout => \phase_controller_inst2.stoper_tr.start_latched_RNI7GMNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110101010"
        )
    port map (
            in0 => \N__33960\,
            in1 => \N__37012\,
            in2 => \N__34143\,
            in3 => \N__33944\,
            lcout => \phase_controller_inst1.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49882\,
            ce => 'H',
            sr => \N__49326\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNID63H_30_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__37011\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34138\,
            lcout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst1.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33963\,
            in3 => \N__33942\,
            lcout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__37010\,
            in1 => \N__33959\,
            in2 => \_gnd_net_\,
            in3 => \N__36980\,
            lcout => \phase_controller_inst1.stoper_hc.un2_start_0\,
            ltout => \phase_controller_inst1.stoper_hc.un2_start_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1_30_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__33951\,
            in3 => \N__33923\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNI2RQB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_1_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__33943\,
            in1 => \N__37590\,
            in2 => \N__33927\,
            in3 => \N__34946\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49882\,
            ce => 'H',
            sr => \N__49326\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37107\,
            in2 => \N__33915\,
            in3 => \N__34942\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_2_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37095\,
            in2 => \N__33906\,
            in3 => \N__35234\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_3_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35210\,
            in1 => \N__34365\,
            in2 => \N__33897\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_4_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37659\,
            in2 => \N__33885\,
            in3 => \N__35195\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_5_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34974\,
            in2 => \N__34050\,
            in3 => \N__35180\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_6_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34038\,
            in2 => \N__34098\,
            in3 => \N__35165\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_7_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34191\,
            in2 => \N__34032\,
            in3 => \N__35150\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_8_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34023\,
            in2 => \N__34011\,
            in3 => \N__35135\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_9_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34170\,
            in2 => \N__33999\,
            in3 => \N__35120\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_10_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33990\,
            in2 => \N__34311\,
            in3 => \N__35333\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_11_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35318\,
            in1 => \N__34329\,
            in2 => \N__33984\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_12_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__35303\,
            in1 => \N__34356\,
            in2 => \N__33972\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_13_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34074\,
            in2 => \N__35424\,
            in3 => \N__35288\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_14_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36939\,
            in2 => \N__34068\,
            in3 => \N__35273\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_inv_15_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34182\,
            in2 => \N__34059\,
            in3 => \N__35258\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_16_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36864\,
            in2 => \N__36927\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_18_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37284\,
            in2 => \N__37083\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_20_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37146\,
            in2 => \N__37029\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_22_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37716\,
            in2 => \N__37776\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_24_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34989\,
            in2 => \N__35004\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_26_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34107\,
            in2 => \N__34116\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_28_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34200\,
            in2 => \N__34281\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_30_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34158\,
            in2 => \N__34404\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34146\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_26_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__35351\,
            in1 => \N__34290\,
            in2 => \N__34086\,
            in3 => \N__35581\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_26_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__34289\,
            in1 => \N__34085\,
            in2 => \N__35583\,
            in3 => \N__35350\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46849\,
            in1 => \N__45443\,
            in2 => \_gnd_net_\,
            in3 => \N__45407\,
            lcout => \elapsed_time_ns_1_RNII43T9_0_6\,
            ltout => \elapsed_time_ns_1_RNII43T9_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_6_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__45444\,
            in1 => \_gnd_net_\,
            in2 => \N__34101\,
            in3 => \N__46853\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => \N__37607\,
            sr => \N__49362\
        );

    \phase_controller_inst1.stoper_hc.target_time_27_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46852\,
            in1 => \N__47121\,
            in2 => \_gnd_net_\,
            in3 => \N__50382\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => \N__37607\,
            sr => \N__49362\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41630\,
            in1 => \N__41597\,
            in2 => \_gnd_net_\,
            in3 => \N__46850\,
            lcout => \elapsed_time_ns_1_RNI47DN9_0_26\,
            ltout => \elapsed_time_ns_1_RNI47DN9_0_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_26_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46851\,
            in1 => \_gnd_net_\,
            in2 => \N__34293\,
            in3 => \N__41631\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49840\,
            ce => \N__37607\,
            sr => \N__49362\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_28_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100010000"
        )
    port map (
            in0 => \N__35562\,
            in1 => \N__35541\,
            in2 => \N__34224\,
            in3 => \N__34209\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46814\,
            in1 => \N__39694\,
            in2 => \_gnd_net_\,
            in3 => \N__34265\,
            lcout => \elapsed_time_ns_1_RNI69DN9_0_28\,
            ltout => \elapsed_time_ns_1_RNI69DN9_0_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_28_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39695\,
            in1 => \_gnd_net_\,
            in2 => \N__34254\,
            in3 => \N__46816\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49831\,
            ce => \N__37608\,
            sr => \N__49369\
        );

    \phase_controller_inst1.stoper_hc.target_time_29_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46815\,
            in1 => \N__34251\,
            in2 => \_gnd_net_\,
            in3 => \N__39649\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49831\,
            ce => \N__37608\,
            sr => \N__49369\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_28_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100110001"
        )
    port map (
            in0 => \N__35561\,
            in1 => \N__35540\,
            in2 => \N__34223\,
            in3 => \N__34208\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_7_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45383\,
            in1 => \N__45354\,
            in2 => \_gnd_net_\,
            in3 => \N__46817\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49831\,
            ce => \N__37608\,
            sr => \N__49369\
        );

    \phase_controller_inst1.stoper_hc.target_time_15_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46916\,
            in1 => \N__45208\,
            in2 => \_gnd_net_\,
            in3 => \N__45191\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => \N__37641\,
            sr => \N__49373\
        );

    \phase_controller_inst1.stoper_hc.target_time_9_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41400\,
            in1 => \N__46921\,
            in2 => \_gnd_net_\,
            in3 => \N__41433\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => \N__37641\,
            sr => \N__49373\
        );

    \phase_controller_inst1.stoper_hc.target_time_3_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46918\,
            in1 => \N__41475\,
            in2 => \_gnd_net_\,
            in3 => \N__41514\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => \N__37641\,
            sr => \N__49373\
        );

    \phase_controller_inst1.stoper_hc.target_time_12_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41343\,
            in1 => \N__46920\,
            in2 => \_gnd_net_\,
            in3 => \N__41376\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => \N__37641\,
            sr => \N__49373\
        );

    \phase_controller_inst1.stoper_hc.target_time_30_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46917\,
            in1 => \N__39600\,
            in2 => \_gnd_net_\,
            in3 => \N__34346\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => \N__37641\,
            sr => \N__49373\
        );

    \phase_controller_inst1.stoper_hc.target_time_11_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40921\,
            in1 => \N__46919\,
            in2 => \_gnd_net_\,
            in3 => \N__40961\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49824\,
            ce => \N__37641\,
            sr => \N__49373\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41375\,
            in1 => \N__40996\,
            in2 => \N__40962\,
            in3 => \N__41432\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI9JET2_5_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__45442\,
            in1 => \N__39316\,
            in2 => \N__34320\,
            in3 => \N__34317\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI32LR_7_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39268\,
            in2 => \_gnd_net_\,
            in3 => \N__45353\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_10_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40997\,
            in1 => \N__41024\,
            in2 => \_gnd_net_\,
            in3 => \N__46724\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49820\,
            ce => \N__37639\,
            sr => \N__49379\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__35439\,
            in1 => \N__34299\,
            in2 => \N__35733\,
            in3 => \N__39561\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3\,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_31_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__39562\,
            in1 => \_gnd_net_\,
            in2 => \N__34458\,
            in3 => \N__34454\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49818\,
            ce => \N__37642\,
            sr => \N__49383\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_30_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110011101111"
        )
    port map (
            in0 => \N__34431\,
            in1 => \N__35477\,
            in2 => \N__35519\,
            in3 => \N__34415\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36795\,
            in2 => \N__41883\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46369\,
            in2 => \N__46338\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47641\,
            in2 => \N__37959\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39504\,
            in2 => \N__47807\,
            in3 => \N__34389\,
            lcout => \current_shift_inst.un38_control_input_0_s1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47645\,
            in2 => \N__39777\,
            in3 => \N__34386\,
            lcout => \current_shift_inst.un38_control_input_0_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39897\,
            in2 => \N__47808\,
            in3 => \N__34371\,
            lcout => \current_shift_inst.un38_control_input_0_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47649\,
            in2 => \N__38133\,
            in3 => \N__34368\,
            lcout => \current_shift_inst.un38_control_input_0_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36039\,
            in2 => \N__47809\,
            in3 => \N__34518\,
            lcout => \current_shift_inst.un38_control_input_0_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47653\,
            in2 => \N__36171\,
            in3 => \N__34515\,
            lcout => \current_shift_inst.un38_control_input_0_s1_8\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39738\,
            in2 => \N__47810\,
            in3 => \N__34500\,
            lcout => \current_shift_inst.un38_control_input_0_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47657\,
            in2 => \N__48336\,
            in3 => \N__34497\,
            lcout => \current_shift_inst.un38_control_input_0_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36162\,
            in2 => \N__47811\,
            in3 => \N__34494\,
            lcout => \current_shift_inst.un38_control_input_0_s1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47661\,
            in2 => \N__48405\,
            in3 => \N__34482\,
            lcout => \current_shift_inst.un38_control_input_0_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47253\,
            in2 => \N__47812\,
            in3 => \N__34473\,
            lcout => \current_shift_inst.un38_control_input_0_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47665\,
            in2 => \N__38217\,
            in3 => \N__34461\,
            lcout => \current_shift_inst.un38_control_input_0_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39789\,
            in2 => \N__47813\,
            in3 => \N__34617\,
            lcout => \current_shift_inst.un38_control_input_0_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47685\,
            in2 => \N__36834\,
            in3 => \N__34605\,
            lcout => \current_shift_inst.un38_control_input_0_s1_16\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36024\,
            in2 => \N__47818\,
            in3 => \N__34593\,
            lcout => \current_shift_inst.un38_control_input_0_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47689\,
            in2 => \N__36033\,
            in3 => \N__34581\,
            lcout => \current_shift_inst.un38_control_input_0_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36012\,
            in2 => \N__47819\,
            in3 => \N__34569\,
            lcout => \current_shift_inst.un38_control_input_0_s1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47693\,
            in2 => \N__39939\,
            in3 => \N__34557\,
            lcout => \current_shift_inst.un38_control_input_0_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36018\,
            in2 => \N__47820\,
            in3 => \N__34545\,
            lcout => \current_shift_inst.un38_control_input_0_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47697\,
            in2 => \N__39966\,
            in3 => \N__34533\,
            lcout => \current_shift_inst.un38_control_input_0_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36147\,
            in2 => \N__47821\,
            in3 => \N__34521\,
            lcout => \current_shift_inst.un38_control_input_0_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47822\,
            in2 => \N__36843\,
            in3 => \N__34701\,
            lcout => \current_shift_inst.un38_control_input_0_s1_24\,
            ltout => OPEN,
            carryin => \bfn_13_19_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42621\,
            in2 => \N__47872\,
            in3 => \N__34698\,
            lcout => \current_shift_inst.un38_control_input_0_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47826\,
            in2 => \N__36852\,
            in3 => \N__34686\,
            lcout => \current_shift_inst.un38_control_input_0_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36132\,
            in2 => \N__47873\,
            in3 => \N__34674\,
            lcout => \current_shift_inst.un38_control_input_0_s1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47830\,
            in2 => \N__36156\,
            in3 => \N__34662\,
            lcout => \current_shift_inst.un38_control_input_0_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36126\,
            in2 => \N__47874\,
            in3 => \N__34647\,
            lcout => \current_shift_inst.un38_control_input_0_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47834\,
            in2 => \N__36141\,
            in3 => \N__34632\,
            lcout => \current_shift_inst.un38_control_input_0_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s1\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__47835\,
            in1 => \N__48255\,
            in2 => \_gnd_net_\,
            in3 => \N__34629\,
            lcout => \current_shift_inst.un38_control_input_0_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.S2_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34734\,
            lcout => s2_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \N__49412\
        );

    \current_shift_inst.start_timer_s1_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__34855\,
            in1 => \N__34836\,
            in2 => \_gnd_net_\,
            in3 => \N__34914\,
            lcout => \current_shift_inst.start_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \N__49412\
        );

    \phase_controller_inst1.S1_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34915\,
            lcout => s1_phy_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49803\,
            ce => 'H',
            sr => \N__49412\
        );

    \current_shift_inst.stop_timer_s1_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__34837\,
            in1 => \N__34815\,
            in2 => \N__34917\,
            in3 => \N__34856\,
            lcout => \current_shift_inst.stop_timer_sZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49800\,
            ce => 'H',
            sr => \N__49417\
        );

    \current_shift_inst.timer_s1.running_LC_13_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__34814\,
            in1 => \N__34838\,
            in2 => \_gnd_net_\,
            in3 => \N__36198\,
            lcout => \current_shift_inst.timer_s1.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49800\,
            ce => 'H',
            sr => \N__49417\
        );

    \current_shift_inst.timer_s1.running_RNIEOIK_LC_13_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__36196\,
            in1 => \N__34813\,
            in2 => \_gnd_net_\,
            in3 => \N__34839\,
            lcout => \current_shift_inst.timer_s1.N_162_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.running_RNII51H_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36195\,
            in2 => \_gnd_net_\,
            in3 => \N__34812\,
            lcout => \current_shift_inst.timer_s1.N_161_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.state_1_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__34782\,
            in1 => \N__34746\,
            in2 => \_gnd_net_\,
            in3 => \N__34726\,
            lcout => \phase_controller_inst1.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49941\,
            ce => 'H',
            sr => \N__49292\
        );

    \phase_controller_inst2.stoper_hc.start_latched_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38984\,
            lcout => \phase_controller_inst2.stoper_hc.start_latchedZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49930\,
            ce => 'H',
            sr => \N__49296\
        );

    \phase_controller_inst2.state_4_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__35035\,
            in1 => \N__35017\,
            in2 => \_gnd_net_\,
            in3 => \N__35086\,
            lcout => \phase_controller_inst2.stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49305\
        );

    \phase_controller_inst2.start_flag_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111000"
        )
    port map (
            in0 => \N__35085\,
            in1 => \N__35036\,
            in2 => \N__35022\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.start_flagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49919\,
            ce => 'H',
            sr => \N__49305\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_24_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__35396\,
            in1 => \N__34962\,
            in2 => \N__36954\,
            in3 => \N__35375\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_24_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__34961\,
            in1 => \N__35397\,
            in2 => \N__35376\,
            in3 => \N__36953\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45038\,
            in1 => \N__45014\,
            in2 => \_gnd_net_\,
            in3 => \N__46956\,
            lcout => \elapsed_time_ns_1_RNI36DN9_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46957\,
            in1 => \N__39317\,
            in2 => \_gnd_net_\,
            in3 => \N__37040\,
            lcout => \elapsed_time_ns_1_RNIH33T9_0_5\,
            ltout => \elapsed_time_ns_1_RNIH33T9_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_5_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__39318\,
            in1 => \_gnd_net_\,
            in2 => \N__34977\,
            in3 => \N__46960\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49908\,
            ce => \N__37643\,
            sr => \N__49312\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40477\,
            in1 => \N__46958\,
            in2 => \_gnd_net_\,
            in3 => \N__40436\,
            lcout => \elapsed_time_ns_1_RNI25DN9_0_24\,
            ltout => \elapsed_time_ns_1_RNI25DN9_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_24_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46959\,
            in1 => \_gnd_net_\,
            in2 => \N__34965\,
            in3 => \N__40478\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49908\,
            ce => \N__37643\,
            sr => \N__49312\
        );

    \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34953\,
            in2 => \N__34947\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_2_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37506\,
            in1 => \N__35235\,
            in2 => \_gnd_net_\,
            in3 => \N__35223\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_3_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__37587\,
            in1 => \N__35211\,
            in2 => \N__35220\,
            in3 => \N__35199\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37507\,
            in1 => \N__35196\,
            in2 => \_gnd_net_\,
            in3 => \N__35184\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37588\,
            in1 => \N__35181\,
            in2 => \_gnd_net_\,
            in3 => \N__35169\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37508\,
            in1 => \N__35166\,
            in2 => \_gnd_net_\,
            in3 => \N__35154\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_7_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37589\,
            in1 => \N__35151\,
            in2 => \_gnd_net_\,
            in3 => \N__35139\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_8_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37509\,
            in1 => \N__35136\,
            in2 => \_gnd_net_\,
            in3 => \N__35124\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49897\,
            ce => 'H',
            sr => \N__49319\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_9_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37586\,
            in1 => \N__35121\,
            in2 => \_gnd_net_\,
            in3 => \N__35109\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_10_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37555\,
            in1 => \N__35334\,
            in2 => \_gnd_net_\,
            in3 => \N__35322\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_11_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37583\,
            in1 => \N__35319\,
            in2 => \_gnd_net_\,
            in3 => \N__35307\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_12_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37556\,
            in1 => \N__35304\,
            in2 => \_gnd_net_\,
            in3 => \N__35292\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_13_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37584\,
            in1 => \N__35289\,
            in2 => \_gnd_net_\,
            in3 => \N__35277\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_14_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37557\,
            in1 => \N__35274\,
            in2 => \_gnd_net_\,
            in3 => \N__35262\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_15_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37585\,
            in1 => \N__35259\,
            in2 => \_gnd_net_\,
            in3 => \N__35247\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_16_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37558\,
            in1 => \N__36912\,
            in2 => \_gnd_net_\,
            in3 => \N__35244\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49883\,
            ce => 'H',
            sr => \N__49327\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_17_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37622\,
            in1 => \N__36880\,
            in2 => \_gnd_net_\,
            in3 => \N__35241\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_18_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37609\,
            in1 => \N__37299\,
            in2 => \_gnd_net_\,
            in3 => \N__35238\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_19_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37623\,
            in1 => \N__37329\,
            in2 => \_gnd_net_\,
            in3 => \N__35412\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_20_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37610\,
            in1 => \N__37163\,
            in2 => \_gnd_net_\,
            in3 => \N__35409\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_21_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37624\,
            in1 => \N__37179\,
            in2 => \_gnd_net_\,
            in3 => \N__35406\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_22_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37611\,
            in1 => \N__37753\,
            in2 => \_gnd_net_\,
            in3 => \N__35403\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_23_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37625\,
            in1 => \N__37732\,
            in2 => \_gnd_net_\,
            in3 => \N__35400\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_24_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37612\,
            in1 => \N__35395\,
            in2 => \_gnd_net_\,
            in3 => \N__35379\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49873\,
            ce => 'H',
            sr => \N__49335\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_25_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37619\,
            in1 => \N__35371\,
            in2 => \_gnd_net_\,
            in3 => \N__35355\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_26_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37626\,
            in1 => \N__35352\,
            in2 => \_gnd_net_\,
            in3 => \N__35337\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_27_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37620\,
            in1 => \N__35582\,
            in2 => \_gnd_net_\,
            in3 => \N__35565\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_28_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37627\,
            in1 => \N__35560\,
            in2 => \_gnd_net_\,
            in3 => \N__35544\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_29_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37621\,
            in1 => \N__35539\,
            in2 => \_gnd_net_\,
            in3 => \N__35523\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_30_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__37628\,
            in1 => \N__35506\,
            in2 => \_gnd_net_\,
            in3 => \N__35484\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst1.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \phase_controller_inst1.stoper_hc.accumulated_time_31_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__35470\,
            in1 => \N__37629\,
            in2 => \_gnd_net_\,
            in3 => \N__35481\,
            lcout => \phase_controller_inst1.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49863\,
            ce => 'H',
            sr => \N__49345\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI52F01_17_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39464\,
            in1 => \N__44663\,
            in2 => \N__47243\,
            in3 => \N__44574\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIQPH01_21_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41558\,
            in1 => \N__41682\,
            in2 => \N__45516\,
            in3 => \N__40468\,
            lcout => OPEN,
            ltout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2S124_13_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__35589\,
            in1 => \N__35448\,
            in2 => \N__35442\,
            in3 => \N__37269\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_13_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44354\,
            in1 => \N__44321\,
            in2 => \_gnd_net_\,
            in3 => \N__46936\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49851\,
            ce => \N__37630\,
            sr => \N__49354\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46812\,
            in1 => \N__37679\,
            in2 => \_gnd_net_\,
            in3 => \N__39353\,
            lcout => \elapsed_time_ns_1_RNIG23T9_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIPMI72_27_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__39693\,
            in1 => \N__37275\,
            in2 => \_gnd_net_\,
            in3 => \N__47112\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46813\,
            in1 => \N__40925\,
            in2 => \_gnd_net_\,
            in3 => \N__40960\,
            lcout => \elapsed_time_ns_1_RNIUVBN9_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45212\,
            in1 => \N__45190\,
            in2 => \_gnd_net_\,
            in3 => \N__46811\,
            lcout => \elapsed_time_ns_1_RNI24CN9_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__35717\,
            in1 => \N__35679\,
            in2 => \_gnd_net_\,
            in3 => \N__35661\,
            lcout => \phase_controller_inst2.stoper_tr.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI56J01_25_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39648\,
            in1 => \N__41624\,
            in2 => \N__39610\,
            in3 => \N__45003\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36794\,
            in2 => \N__41445\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_13_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_0_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46359\,
            in2 => \N__41853\,
            in3 => \N__38271\,
            lcout => \current_shift_inst.un38_control_input_5_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_0_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_1_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__38272\,
            in1 => \N__47379\,
            in2 => \N__37380\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un38_control_input_5_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_1_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_2_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37815\,
            in2 => \N__47584\,
            in3 => \N__35784\,
            lcout => \current_shift_inst.un38_control_input_0_s0_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_2_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_3_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47383\,
            in2 => \N__41802\,
            in3 => \N__35781\,
            lcout => \current_shift_inst.un38_control_input_0_s0_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_3_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_4_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39750\,
            in2 => \N__47585\,
            in3 => \N__35766\,
            lcout => \current_shift_inst.un38_control_input_0_s0_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_4_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_5_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47387\,
            in2 => \N__37983\,
            in3 => \N__35763\,
            lcout => \current_shift_inst.un38_control_input_0_s0_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_5_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_6_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37800\,
            in2 => \N__47586\,
            in3 => \N__35760\,
            lcout => \current_shift_inst.un38_control_input_0_s0_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_6_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_7_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47391\,
            in2 => \N__37932\,
            in3 => \N__35757\,
            lcout => \current_shift_inst.un38_control_input_0_s0_8\,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_8_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37923\,
            in2 => \N__47587\,
            in3 => \N__35742\,
            lcout => \current_shift_inst.un38_control_input_0_s0_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_8_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_9_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47395\,
            in2 => \N__37809\,
            in3 => \N__35739\,
            lcout => \current_shift_inst.un38_control_input_0_s0_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_9_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_10_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37785\,
            in2 => \N__47588\,
            in3 => \N__35736\,
            lcout => \current_shift_inst.un38_control_input_0_s0_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_10_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_11_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47399\,
            in2 => \N__37794\,
            in3 => \N__35898\,
            lcout => \current_shift_inst.un38_control_input_0_s0_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_11_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_12_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39909\,
            in2 => \N__47589\,
            in3 => \N__35883\,
            lcout => \current_shift_inst.un38_control_input_0_s0_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_12_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_13_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47403\,
            in2 => \N__37974\,
            in3 => \N__35868\,
            lcout => \current_shift_inst.un38_control_input_0_s0_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_13_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_14_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37965\,
            in2 => \N__47590\,
            in3 => \N__35853\,
            lcout => \current_shift_inst.un38_control_input_0_s0_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_14_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_15_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47669\,
            in2 => \N__38088\,
            in3 => \N__35841\,
            lcout => \current_shift_inst.un38_control_input_0_s0_16\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_16_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37917\,
            in2 => \N__47814\,
            in3 => \N__35829\,
            lcout => \current_shift_inst.un38_control_input_0_s0_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_16_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_17_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47673\,
            in2 => \N__38010\,
            in3 => \N__35817\,
            lcout => \current_shift_inst.un38_control_input_0_s0_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_17_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_18_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37911\,
            in2 => \N__47815\,
            in3 => \N__35802\,
            lcout => \current_shift_inst.un38_control_input_0_s0_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_18_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_19_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47677\,
            in2 => \N__48270\,
            in3 => \N__35787\,
            lcout => \current_shift_inst.un38_control_input_0_s0_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_19_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_20_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38205\,
            in2 => \N__47816\,
            in3 => \N__35988\,
            lcout => \current_shift_inst.un38_control_input_0_s0_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_20_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_21_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47681\,
            in2 => \N__37944\,
            in3 => \N__35973\,
            lcout => \current_shift_inst.un38_control_input_0_s0_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_21_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_22_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38226\,
            in2 => \N__47817\,
            in3 => \N__35958\,
            lcout => \current_shift_inst.un38_control_input_0_s0_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_22_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_23_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36006\,
            in2 => \N__47836\,
            in3 => \N__35955\,
            lcout => \current_shift_inst.un38_control_input_0_s0_24\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \current_shift_inst.un38_control_input_cry_24_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47721\,
            in2 => \N__38196\,
            in3 => \N__35952\,
            lcout => \current_shift_inst.un38_control_input_0_s0_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_24_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_25_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37992\,
            in2 => \N__47837\,
            in3 => \N__35940\,
            lcout => \current_shift_inst.un38_control_input_0_s0_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_25_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_26_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47725\,
            in2 => \N__38187\,
            in3 => \N__35928\,
            lcout => \current_shift_inst.un38_control_input_0_s0_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_26_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_27_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36177\,
            in2 => \N__47838\,
            in3 => \N__35913\,
            lcout => \current_shift_inst.un38_control_input_0_s0_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_27_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_28_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47729\,
            in2 => \N__38175\,
            in3 => \N__36081\,
            lcout => \current_shift_inst.un38_control_input_0_s0_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_28_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_29_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37998\,
            in2 => \N__47839\,
            in3 => \N__36066\,
            lcout => \current_shift_inst.un38_control_input_0_s0_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un38_control_input_cry_29_s0\,
            carryout => \current_shift_inst.un38_control_input_cry_30_s0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__46590\,
            in1 => \N__36063\,
            in2 => \N__38499\,
            in3 => \N__36051\,
            lcout => \current_shift_inst.control_input_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48208\,
            in1 => \N__47741\,
            in2 => \N__40037\,
            in3 => \N__42009\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__47739\,
            in1 => \N__48211\,
            in2 => \N__42180\,
            in3 => \N__43164\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48210\,
            in1 => \N__47746\,
            in2 => \N__40562\,
            in3 => \N__42211\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__47743\,
            in1 => \N__48213\,
            in2 => \N__42093\,
            in3 => \N__40326\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__48212\,
            in1 => \N__42140\,
            in2 => \N__42612\,
            in3 => \N__47744\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47745\,
            in1 => \N__48214\,
            in2 => \N__43061\,
            in3 => \N__42485\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48215\,
            in1 => \N__47740\,
            in2 => \N__43014\,
            in3 => \N__42389\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47742\,
            in1 => \N__48209\,
            in2 => \N__42713\,
            in3 => \N__41976\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48216\,
            in1 => \N__43382\,
            in2 => \N__47847\,
            in3 => \N__43344\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42390\,
            in1 => \N__47750\,
            in2 => \N__43013\,
            in3 => \N__48222\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI5C531_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \N__47754\,
            in1 => \N__42519\,
            in2 => \N__48251\,
            in3 => \N__40221\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__42310\,
            in1 => \N__47757\,
            in2 => \N__38277\,
            in3 => \N__48224\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__48221\,
            in1 => \N__42419\,
            in2 => \N__47846\,
            in3 => \N__42908\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42353\,
            in1 => \N__47755\,
            in2 => \N__43532\,
            in3 => \N__48223\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__36120\,
            in1 => \N__36111\,
            in2 => \_gnd_net_\,
            in3 => \N__38485\,
            lcout => \current_shift_inst.control_input_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__42457\,
            in1 => \N__47756\,
            in2 => \N__42959\,
            in3 => \N__48220\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47870\,
            in1 => \N__48253\,
            in2 => \N__43062\,
            in3 => \N__42489\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPR031_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110001101"
        )
    port map (
            in0 => \N__48252\,
            in1 => \N__42249\,
            in2 => \N__43260\,
            in3 => \N__47871\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38442\,
            in1 => \N__36822\,
            in2 => \_gnd_net_\,
            in3 => \N__36816\,
            lcout => \current_shift_inst.control_input_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__41882\,
            in1 => \N__38754\,
            in2 => \_gnd_net_\,
            in3 => \N__38253\,
            lcout => \current_shift_inst.un38_control_input_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__36223\,
            in1 => \N__36774\,
            in2 => \_gnd_net_\,
            in3 => \N__36723\,
            lcout => \elapsed_time_ns_1_RNI4EOBB_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_inv_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__46553\,
            in1 => \N__38753\,
            in2 => \_gnd_net_\,
            in3 => \N__36204\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46525\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_fast_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49809\,
            ce => \N__46406\,
            sr => \N__49405\
        );

    \current_shift_inst.timer_s1.running_RNIUKI8_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36197\,
            lcout => \current_shift_inst.timer_s1.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__39001\,
            in1 => \N__38291\,
            in2 => \_gnd_net_\,
            in3 => \N__38980\,
            lcout => \phase_controller_inst2.stoper_hc.un2_start_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.start_latched_RNIFLAI_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37013\,
            in2 => \_gnd_net_\,
            in3 => \N__36981\,
            lcout => \phase_controller_inst1.stoper_hc.start_latched_RNIFLAIZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_17_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44589\,
            in1 => \N__44612\,
            in2 => \_gnd_net_\,
            in3 => \N__47038\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49931\,
            ce => \N__37518\,
            sr => \N__49297\
        );

    \phase_controller_inst1.stoper_hc.target_time_25_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45034\,
            in1 => \N__47076\,
            in2 => \_gnd_net_\,
            in3 => \N__45015\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49920\,
            ce => \N__37644\,
            sr => \N__49306\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44545\,
            in1 => \N__44513\,
            in2 => \_gnd_net_\,
            in3 => \N__47029\,
            lcout => \elapsed_time_ns_1_RNI13CN9_0_14\,
            ltout => \elapsed_time_ns_1_RNI13CN9_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_14_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47030\,
            in1 => \_gnd_net_\,
            in2 => \N__36942\,
            in3 => \N__44546\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => \N__37597\,
            sr => \N__49313\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44611\,
            in1 => \N__44584\,
            in2 => \_gnd_net_\,
            in3 => \N__47028\,
            lcout => \elapsed_time_ns_1_RNI46CN9_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_16_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010011110101"
        )
    port map (
            in0 => \N__36881\,
            in1 => \N__37067\,
            in2 => \N__36897\,
            in3 => \N__36910\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_16_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011011100"
        )
    port map (
            in0 => \N__36911\,
            in1 => \N__36893\,
            in2 => \N__37068\,
            in3 => \N__36882\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44416\,
            in1 => \N__47027\,
            in2 => \_gnd_net_\,
            in3 => \N__44375\,
            lcout => \elapsed_time_ns_1_RNI35CN9_0_16\,
            ltout => \elapsed_time_ns_1_RNI35CN9_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_16_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47031\,
            in1 => \_gnd_net_\,
            in2 => \N__37071\,
            in3 => \N__44417\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49909\,
            ce => \N__37597\,
            sr => \N__49313\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__40710\,
            in1 => \N__40733\,
            in2 => \N__37056\,
            in3 => \N__47190\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_18_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__47189\,
            in1 => \N__40709\,
            in2 => \N__40737\,
            in3 => \N__37052\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_19_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37263\,
            in1 => \N__39465\,
            in2 => \_gnd_net_\,
            in3 => \N__47035\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49898\,
            ce => \N__47156\,
            sr => \N__49320\
        );

    \phase_controller_inst2.stoper_hc.target_time_2_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__47033\,
            in1 => \N__37200\,
            in2 => \N__39537\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49898\,
            ce => \N__47156\,
            sr => \N__49320\
        );

    \phase_controller_inst2.stoper_hc.target_time_3_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41474\,
            in1 => \N__41509\,
            in2 => \_gnd_net_\,
            in3 => \N__47036\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49898\,
            ce => \N__47156\,
            sr => \N__49320\
        );

    \phase_controller_inst2.stoper_hc.target_time_4_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47034\,
            in1 => \N__37683\,
            in2 => \_gnd_net_\,
            in3 => \N__39352\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49898\,
            ce => \N__47156\,
            sr => \N__49320\
        );

    \phase_controller_inst2.stoper_hc.target_time_5_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37044\,
            in1 => \N__39315\,
            in2 => \_gnd_net_\,
            in3 => \N__47037\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49898\,
            ce => \N__47156\,
            sr => \N__49320\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_20_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000101010000"
        )
    port map (
            in0 => \N__37178\,
            in1 => \N__37159\,
            in2 => \N__37131\,
            in3 => \N__37116\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_20_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__37115\,
            in1 => \N__37177\,
            in2 => \N__37164\,
            in3 => \N__37130\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__46965\,
            in1 => \_gnd_net_\,
            in2 => \N__45514\,
            in3 => \N__45467\,
            lcout => \elapsed_time_ns_1_RNIV1DN9_0_21\,
            ltout => \elapsed_time_ns_1_RNIV1DN9_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_21_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45507\,
            in2 => \N__37134\,
            in3 => \N__46970\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__37519\,
            sr => \N__49328\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46964\,
            in1 => \N__44661\,
            in2 => \_gnd_net_\,
            in3 => \N__44624\,
            lcout => \elapsed_time_ns_1_RNIU0DN9_0_20\,
            ltout => \elapsed_time_ns_1_RNIU0DN9_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_20_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__44662\,
            in1 => \_gnd_net_\,
            in2 => \N__37119\,
            in3 => \N__46969\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__37519\,
            sr => \N__49328\
        );

    \phase_controller_inst1.stoper_hc.target_time_1_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__50325\,
            in1 => \_gnd_net_\,
            in2 => \N__47039\,
            in3 => \N__45146\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__37519\,
            sr => \N__49328\
        );

    \phase_controller_inst1.stoper_hc.target_time_2_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37199\,
            in1 => \N__39533\,
            in2 => \_gnd_net_\,
            in3 => \N__46971\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49884\,
            ce => \N__37519\,
            sr => \N__49328\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_18_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010110010"
        )
    port map (
            in0 => \N__37338\,
            in1 => \N__37328\,
            in2 => \N__37313\,
            in3 => \N__37298\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47232\,
            in1 => \N__47058\,
            in2 => \_gnd_net_\,
            in3 => \N__47201\,
            lcout => \elapsed_time_ns_1_RNI57CN9_0_18\,
            ltout => \elapsed_time_ns_1_RNI57CN9_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_18_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__47059\,
            in1 => \_gnd_net_\,
            in2 => \N__37341\,
            in3 => \N__47233\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__37634\,
            sr => \N__49336\
        );

    \phase_controller_inst1.stoper_hc.target_time_19_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37258\,
            in1 => \N__39460\,
            in2 => \_gnd_net_\,
            in3 => \N__47060\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49874\,
            ce => \N__37634\,
            sr => \N__49336\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_18_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001011110011"
        )
    port map (
            in0 => \N__37337\,
            in1 => \N__37327\,
            in2 => \N__37314\,
            in3 => \N__37297\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41496\,
            in1 => \N__39337\,
            in2 => \N__39532\,
            in3 => \N__50319\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUPD01_13_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__45172\,
            in1 => \N__44530\,
            in2 => \N__44407\,
            in3 => \N__44310\,
            lcout => \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__37262\,
            in1 => \N__39450\,
            in2 => \_gnd_net_\,
            in3 => \N__46934\,
            lcout => \elapsed_time_ns_1_RNI68CN9_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_30_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011111011"
        )
    port map (
            in0 => \N__37242\,
            in1 => \N__41318\,
            in2 => \N__41127\,
            in3 => \N__37221\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46935\,
            in1 => \N__37198\,
            in2 => \_gnd_net_\,
            in3 => \N__39525\,
            lcout => \elapsed_time_ns_1_RNIE03T9_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46933\,
            in1 => \N__45376\,
            in2 => \_gnd_net_\,
            in3 => \N__45342\,
            lcout => \elapsed_time_ns_1_RNIJ53T9_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_0_22_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__37704\,
            in1 => \N__37692\,
            in2 => \N__37758\,
            in3 => \N__37736\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNO_22_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__37691\,
            in1 => \N__37757\,
            in2 => \N__37737\,
            in3 => \N__37703\,
            lcout => \phase_controller_inst1.stoper_hc.un4_running_cry_c_RNOZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_23_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46942\,
            in1 => \N__41585\,
            in2 => \_gnd_net_\,
            in3 => \N__41550\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49852\,
            ce => \N__37640\,
            sr => \N__49355\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41676\,
            in1 => \N__46940\,
            in2 => \_gnd_net_\,
            in3 => \N__41651\,
            lcout => \elapsed_time_ns_1_RNI03DN9_0_22\,
            ltout => \elapsed_time_ns_1_RNI03DN9_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst1.stoper_hc.target_time_22_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__46941\,
            in1 => \_gnd_net_\,
            in2 => \N__37695\,
            in3 => \N__41677\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49852\,
            ce => \N__37640\,
            sr => \N__49355\
        );

    \phase_controller_inst1.stoper_hc.target_time_4_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46943\,
            in1 => \N__37675\,
            in2 => \_gnd_net_\,
            in3 => \N__39354\,
            lcout => \phase_controller_inst1.stoper_hc.target_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49852\,
            ce => \N__37640\,
            sr => \N__49355\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48093\,
            in1 => \N__47419\,
            in2 => \N__40095\,
            in3 => \N__41778\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITRK61_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__38427\,
            in1 => \N__37371\,
            in2 => \_gnd_net_\,
            in3 => \N__37365\,
            lcout => \current_shift_inst.control_input_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39264\,
            in1 => \N__37900\,
            in2 => \_gnd_net_\,
            in3 => \N__46881\,
            lcout => \elapsed_time_ns_1_RNIK63T9_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__38428\,
            in1 => \N__37881\,
            in2 => \_gnd_net_\,
            in3 => \N__37866\,
            lcout => \current_shift_inst.control_input_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__37848\,
            in1 => \N__37842\,
            in2 => \_gnd_net_\,
            in3 => \N__38426\,
            lcout => \current_shift_inst.control_input_axb_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47418\,
            in1 => \N__48094\,
            in2 => \N__42870\,
            in3 => \N__41751\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48393\,
            in1 => \N__48166\,
            in2 => \N__47610\,
            in3 => \N__48360\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48165\,
            in1 => \N__47426\,
            in2 => \N__40041\,
            in3 => \N__42008\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__47428\,
            in1 => \N__48168\,
            in2 => \N__48432\,
            in3 => \N__48467\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41023\,
            in1 => \N__41001\,
            in2 => \_gnd_net_\,
            in3 => \N__46912\,
            lcout => \elapsed_time_ns_1_RNITUBN9_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47427\,
            in1 => \N__48167\,
            in2 => \N__43383\,
            in3 => \N__43343\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42759\,
            in1 => \N__48164\,
            in2 => \N__47611\,
            in3 => \N__42053\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__48169\,
            in1 => \N__47429\,
            in2 => \N__43448\,
            in3 => \N__43485\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47616\,
            in1 => \N__48082\,
            in2 => \N__43110\,
            in3 => \N__42279\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48079\,
            in1 => \N__47618\,
            in2 => \N__40094\,
            in3 => \N__41774\,
            lcout => \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47614\,
            in1 => \N__48085\,
            in2 => \N__40263\,
            in3 => \N__42558\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48080\,
            in1 => \N__47613\,
            in2 => \N__42714\,
            in3 => \N__41972\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47612\,
            in1 => \N__48081\,
            in2 => \N__40170\,
            in3 => \N__41943\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48083\,
            in1 => \N__47617\,
            in2 => \N__40563\,
            in3 => \N__42213\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__47615\,
            in1 => \N__48084\,
            in2 => \N__42141\,
            in3 => \N__42605\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__38163\,
            in1 => \N__38154\,
            in2 => \_gnd_net_\,
            in3 => \N__38430\,
            lcout => \current_shift_inst.control_input_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48207\,
            in1 => \N__42758\,
            in2 => \N__47795\,
            in3 => \N__42054\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__38121\,
            in1 => \N__38112\,
            in2 => \_gnd_net_\,
            in3 => \N__38431\,
            lcout => \current_shift_inst.control_input_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__47623\,
            in1 => \N__48243\,
            in2 => \N__42248\,
            in3 => \N__43256\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100111"
        )
    port map (
            in0 => \N__38432\,
            in1 => \N__38076\,
            in2 => \N__38067\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.control_input_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110011"
        )
    port map (
            in0 => \N__38040\,
            in1 => \N__38031\,
            in2 => \_gnd_net_\,
            in3 => \N__38429\,
            lcout => \current_shift_inst.control_input_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47619\,
            in1 => \N__48244\,
            in2 => \N__43163\,
            in3 => \N__42176\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110011"
        )
    port map (
            in0 => \N__38276\,
            in1 => \N__48228\,
            in2 => \N__42318\,
            in3 => \N__47863\,
            lcout => \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48235\,
            in1 => \N__47862\,
            in2 => \N__42960\,
            in3 => \N__42458\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48227\,
            in1 => \N__40220\,
            in2 => \N__47879\,
            in3 => \N__42515\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111010001"
        )
    port map (
            in0 => \N__43484\,
            in1 => \N__48225\,
            in2 => \N__43452\,
            in3 => \N__47857\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__48226\,
            in1 => \N__42085\,
            in2 => \N__47878\,
            in3 => \N__40325\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47861\,
            in1 => \N__48234\,
            in2 => \N__43209\,
            in3 => \N__42657\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47848\,
            in1 => \N__48236\,
            in2 => \N__42912\,
            in3 => \N__42418\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48237\,
            in1 => \N__47849\,
            in2 => \N__43533\,
            in3 => \N__42352\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40008\,
            lcout => \current_shift_inst.un4_control_input_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41575\,
            in1 => \N__41559\,
            in2 => \_gnd_net_\,
            in3 => \N__46955\,
            lcout => \elapsed_time_ns_1_RNI14DN9_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40203\,
            lcout => \current_shift_inst.un4_control_input_1_axb_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_0_c_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38249\,
            in2 => \N__46554\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_21_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38803\,
            in2 => \N__48486\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_0\,
            carryout => \current_shift_inst.un10_control_input_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39477\,
            in2 => \N__38849\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_1\,
            carryout => \current_shift_inst.un10_control_input_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38807\,
            in2 => \N__39816\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_2\,
            carryout => \current_shift_inst.un10_control_input_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39762\,
            in2 => \N__38850\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_3\,
            carryout => \current_shift_inst.un10_control_input_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38811\,
            in2 => \N__39711\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_4\,
            carryout => \current_shift_inst.un10_control_input_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39801\,
            in2 => \N__38851\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_5\,
            carryout => \current_shift_inst.un10_control_input_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_7_c_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38815\,
            in2 => \N__39492\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_6\,
            carryout => \current_shift_inst.un10_control_input_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38693\,
            in2 => \N__39888\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_22_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39828\,
            in2 => \N__38749\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_8\,
            carryout => \current_shift_inst.un10_control_input_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38681\,
            in2 => \N__39843\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_9\,
            carryout => \current_shift_inst.un10_control_input_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43314\,
            in2 => \N__38746\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_10\,
            carryout => \current_shift_inst.un10_control_input_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38685\,
            in2 => \N__39981\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_11\,
            carryout => \current_shift_inst.un10_control_input_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43392\,
            in2 => \N__38747\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_12\,
            carryout => \current_shift_inst.un10_control_input_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38689\,
            in2 => \N__43407\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_13\,
            carryout => \current_shift_inst.un10_control_input_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39726\,
            in2 => \N__38748\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_14\,
            carryout => \current_shift_inst.un10_control_input_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39870\,
            in2 => \N__38759\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_23_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38724\,
            in2 => \N__40518\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_16\,
            carryout => \current_shift_inst.un10_control_input_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_LC_15_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40332\,
            in2 => \N__38760\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_17\,
            carryout => \current_shift_inst.un10_control_input_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38728\,
            in2 => \N__40347\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_18\,
            carryout => \current_shift_inst.un10_control_input_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_LC_15_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40107\,
            in2 => \N__38761\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_19\,
            carryout => \current_shift_inst.un10_control_input_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_LC_15_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38732\,
            in2 => \N__40293\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_20\,
            carryout => \current_shift_inst.un10_control_input_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39858\,
            in2 => \N__38762\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_21\,
            carryout => \current_shift_inst.un10_control_input_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_LC_15_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38736\,
            in2 => \N__39924\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_22\,
            carryout => \current_shift_inst.un10_control_input_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38816\,
            in2 => \N__39954\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_24_0_\,
            carryout => \current_shift_inst.un10_control_input_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40500\,
            in2 => \N__38852\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_24\,
            carryout => \current_shift_inst.un10_control_input_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38820\,
            in2 => \N__40284\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_25\,
            carryout => \current_shift_inst.un10_control_input_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40338\,
            in2 => \N__38853\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_26\,
            carryout => \current_shift_inst.un10_control_input_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38824\,
            in2 => \N__40494\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_27\,
            carryout => \current_shift_inst.un10_control_input_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40485\,
            in2 => \N__38854\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_28\,
            carryout => \current_shift_inst.un10_control_input_cry_29\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_LC_15_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38828\,
            in2 => \N__40509\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \current_shift_inst.un10_control_input_cry_29\,
            carryout => \current_shift_inst.un10_control_input_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__48242\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38502\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.time_passed_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010001011100010"
        )
    port map (
            in0 => \N__38316\,
            in1 => \N__39060\,
            in2 => \N__39027\,
            in3 => \N__39372\,
            lcout => \phase_controller_inst2.hc_time_passed\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49293\
        );

    \phase_controller_inst2.stoper_hc.running_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111000101110"
        )
    port map (
            in0 => \N__38292\,
            in1 => \N__39059\,
            in2 => \N__39026\,
            in3 => \N__39371\,
            lcout => \phase_controller_inst2.stoper_hc.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49942\,
            ce => 'H',
            sr => \N__49293\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNIFU8H_30_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39018\,
            in2 => \_gnd_net_\,
            in3 => \N__39370\,
            lcout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i\,
            ltout => \phase_controller_inst2.stoper_hc.running_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38280\,
            in3 => \N__39061\,
            lcout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_1_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__39063\,
            in1 => \N__41215\,
            in2 => \N__39039\,
            in3 => \N__40418\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49932\,
            ce => 'H',
            sr => \N__49298\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1_30_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39062\,
            in2 => \_gnd_net_\,
            in3 => \N__39035\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNI7COB1Z0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.start_latched_RNIHS8D_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__38985\,
            lcout => \phase_controller_inst2.stoper_hc.start_latched_RNIHS8DZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_1_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45117\,
            in2 => \N__38949\,
            in3 => \N__40414\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_1\,
            ltout => OPEN,
            carryin => \bfn_16_7_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_2_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40397\,
            in1 => \N__38937\,
            in2 => \N__38931\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_3_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40373\,
            in1 => \N__38922\,
            in2 => \N__38916\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_4_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38904\,
            in2 => \N__38898\,
            in3 => \N__40682\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_5_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38889\,
            in2 => \N__38883\,
            in3 => \N__40667\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_6_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45396\,
            in2 => \N__38871\,
            in3 => \N__40652\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_7_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45321\,
            in2 => \N__39147\,
            in3 => \N__40637\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_8_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39138\,
            in2 => \N__39123\,
            in3 => \N__40622\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_7\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_9_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40607\,
            in1 => \N__40881\,
            in2 => \N__39114\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_9\,
            ltout => OPEN,
            carryin => \bfn_16_8_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_10_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40971\,
            in2 => \N__39105\,
            in3 => \N__40592\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_11_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39096\,
            in2 => \N__40905\,
            in3 => \N__40577\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_12_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40893\,
            in2 => \N__39090\,
            in3 => \N__40802\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_13_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45225\,
            in2 => \N__39081\,
            in3 => \N__40787\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_14_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40772\,
            in1 => \N__44502\,
            in2 => \N__39072\,
            in3 => \_gnd_net_\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_inv_15_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39228\,
            in2 => \N__45159\,
            in3 => \N__40757\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_time_i_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_16_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44490\,
            in2 => \N__44433\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_15\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_18_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39222\,
            in2 => \N__39210\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_20_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44889\,
            in2 => \N__45531\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_22_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41037\,
            in2 => \N__41097\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_24_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45105\,
            in2 => \N__45051\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_26_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44898\,
            in2 => \N__44961\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_28_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39201\,
            in2 => \N__39186\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_30_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39171\,
            in2 => \N__39162\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un4_running_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un4_running_cry_30\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_LUT4_0_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39375\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_30_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45272\,
            in2 => \N__50355\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45248\,
            in2 => \N__45306\,
            in3 => \N__39321\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45273\,
            in2 => \N__45815\,
            in3 => \N__39282\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45249\,
            in2 => \N__45785\,
            in3 => \N__39279\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45755\,
            in2 => \N__45816\,
            in3 => \N__39276\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45731\,
            in2 => \N__45786\,
            in3 => \N__39234\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45756\,
            in2 => \N__45707\,
            in3 => \N__39231\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45732\,
            in2 => \N__45668\,
            in3 => \N__39402\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9\,
            clk => \N__49885\,
            ce => \N__50238\,
            sr => \N__49329\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45626\,
            in2 => \N__45708\,
            in3 => \N__39399\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11\,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45599\,
            in2 => \N__45669\,
            in3 => \N__39396\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46085\,
            in2 => \N__45630\,
            in3 => \N__39393\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45600\,
            in2 => \N__46058\,
            in3 => \N__39390\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46025\,
            in2 => \N__46089\,
            in3 => \N__39387\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45998\,
            in2 => \N__46059\,
            in3 => \N__39384\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45971\,
            in2 => \N__46029\,
            in3 => \N__39381\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45999\,
            in2 => \N__45938\,
            in3 => \N__39378\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17\,
            clk => \N__49875\,
            ce => \N__50233\,
            sr => \N__49337\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45902\,
            in2 => \N__45975\,
            in3 => \N__39429\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19\,
            ltout => OPEN,
            carryin => \bfn_16_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45872\,
            in2 => \N__45939\,
            in3 => \N__39426\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45842\,
            in2 => \N__45906\,
            in3 => \N__39423\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46322\,
            in2 => \N__45876\,
            in3 => \N__39420\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46292\,
            in2 => \N__45846\,
            in3 => \N__39417\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46265\,
            in2 => \N__46326\,
            in3 => \N__39414\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46238\,
            in2 => \N__46296\,
            in3 => \N__39411\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46266\,
            in2 => \N__46205\,
            in3 => \N__39408\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25\,
            clk => \N__49864\,
            ce => \N__50234\,
            sr => \N__49346\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46166\,
            in2 => \N__46242\,
            in3 => \N__39405\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27\,
            ltout => OPEN,
            carryin => \bfn_16_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            clk => \N__49853\,
            ce => \N__50226\,
            sr => \N__49356\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46139\,
            in2 => \N__46206\,
            in3 => \N__39657\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            clk => \N__49853\,
            ce => \N__50226\,
            sr => \N__49356\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46167\,
            in2 => \N__46113\,
            in3 => \N__39615\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            clk => \N__49853\,
            ce => \N__50226\,
            sr => \N__49356\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46608\,
            in2 => \N__46143\,
            in3 => \N__39573\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28\,
            carryout => \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29\,
            clk => \N__49853\,
            ce => \N__50226\,
            sr => \N__49356\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39570\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => \N__50226\,
            sr => \N__49356\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45305\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49853\,
            ce => \N__50226\,
            sr => \N__49356\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48087\,
            in1 => \N__42859\,
            in2 => \N__47875\,
            in3 => \N__41744\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI00M61_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46529\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49841\,
            ce => \N__46411\,
            sr => \N__49363\
        );

    \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40027\,
            in1 => \N__48584\,
            in2 => \_gnd_net_\,
            in3 => \N__41995\,
            lcout => \current_shift_inst.un10_control_input_cry_7_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48580\,
            in1 => \N__40081\,
            in2 => \_gnd_net_\,
            in3 => \N__41767\,
            lcout => \current_shift_inst.un10_control_input_cry_2_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42866\,
            in1 => \N__48581\,
            in2 => \_gnd_net_\,
            in3 => \N__41743\,
            lcout => \current_shift_inst.un10_control_input_cry_3_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48583\,
            in1 => \_gnd_net_\,
            in2 => \N__42757\,
            in3 => \N__42040\,
            lcout => \current_shift_inst.un10_control_input_cry_6_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \N__47801\,
            in1 => \N__48091\,
            in2 => \N__42278\,
            in3 => \N__43103\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110100011"
        )
    port map (
            in0 => \N__41717\,
            in1 => \N__41837\,
            in2 => \N__48198\,
            in3 => \N__47799\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__41836\,
            in1 => \N__48582\,
            in2 => \_gnd_net_\,
            in3 => \N__41716\,
            lcout => \current_shift_inst.un10_control_input_cry_4_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010101"
        )
    port map (
            in0 => \N__42819\,
            in1 => \N__47800\,
            in2 => \N__41700\,
            in3 => \N__48092\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48186\,
            in1 => \N__47796\,
            in2 => \N__40166\,
            in3 => \N__41936\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43102\,
            in1 => \N__48624\,
            in2 => \_gnd_net_\,
            in3 => \N__42268\,
            lcout => \current_shift_inst.un10_control_input_cry_15_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48622\,
            in1 => \_gnd_net_\,
            in2 => \N__42817\,
            in3 => \N__41695\,
            lcout => \current_shift_inst.un10_control_input_cry_5_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100000011"
        )
    port map (
            in0 => \N__47798\,
            in1 => \N__48187\,
            in2 => \N__47918\,
            in3 => \N__47272\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40080\,
            lcout => \current_shift_inst.un4_control_input_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41827\,
            lcout => \current_shift_inst.un4_control_input_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48185\,
            in1 => \N__47797\,
            in2 => \N__42818\,
            in3 => \N__41696\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI68O61_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42697\,
            in1 => \N__48623\,
            in2 => \_gnd_net_\,
            in3 => \N__41965\,
            lcout => \current_shift_inst.un10_control_input_cry_8_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48628\,
            in1 => \N__43249\,
            in2 => \_gnd_net_\,
            in3 => \N__42235\,
            lcout => \current_shift_inst.un10_control_input_cry_16_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48638\,
            in1 => \N__40256\,
            in2 => \_gnd_net_\,
            in3 => \N__42550\,
            lcout => \current_shift_inst.un10_control_input_cry_22_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__48626\,
            in1 => \N__48352\,
            in2 => \_gnd_net_\,
            in3 => \N__48385\,
            lcout => \current_shift_inst.un10_control_input_cry_10_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__40159\,
            in1 => \N__41935\,
            in2 => \_gnd_net_\,
            in3 => \N__48625\,
            lcout => \current_shift_inst.un10_control_input_cry_9_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40158\,
            lcout => \current_shift_inst.un4_control_input_1_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48460\,
            in1 => \N__48627\,
            in2 => \_gnd_net_\,
            in3 => \N__48421\,
            lcout => \current_shift_inst.un10_control_input_cry_12_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48384\,
            lcout => \current_shift_inst.un4_control_input_1_axb_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43371\,
            lcout => \current_shift_inst.un4_control_input_1_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40317\,
            lcout => \current_shift_inst.un4_control_input_1_axb_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40249\,
            in1 => \N__48197\,
            in2 => \N__47877\,
            in3 => \N__42551\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40548\,
            lcout => \current_shift_inst.un4_control_input_1_axb_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48640\,
            in1 => \N__43048\,
            in2 => \_gnd_net_\,
            in3 => \N__42478\,
            lcout => \current_shift_inst.un10_control_input_cry_24_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__48196\,
            in1 => \N__47853\,
            in2 => \N__48291\,
            in3 => \N__48314\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48639\,
            in1 => \N__40213\,
            in2 => \_gnd_net_\,
            in3 => \N__42508\,
            lcout => \current_shift_inst.un10_control_input_cry_23_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48644\,
            in1 => \N__48313\,
            in2 => \_gnd_net_\,
            in3 => \N__48286\,
            lcout => \current_shift_inst.un10_control_input_cry_20_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__40248\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46490\,
            in2 => \N__43299\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_3\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46439\,
            in2 => \N__43805\,
            in3 => \N__40053\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43298\,
            in2 => \N__43775\,
            in3 => \N__40050\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43742\,
            in2 => \N__43806\,
            in3 => \N__40047\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43715\,
            in2 => \N__43776\,
            in3 => \N__40044\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43691\,
            in2 => \N__43746\,
            in3 => \N__39987\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43716\,
            in2 => \N__43667\,
            in3 => \N__39984\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43692\,
            in2 => \N__43635\,
            in3 => \N__40134\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9\,
            clk => \N__49816\,
            ce => \N__46410\,
            sr => \N__49388\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43592\,
            in2 => \N__43668\,
            in3 => \N__40131\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_11\,
            ltout => OPEN,
            carryin => \bfn_16_20_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43565\,
            in2 => \N__43634\,
            in3 => \N__40128\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44033\,
            in2 => \N__43596\,
            in3 => \N__40125\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43566\,
            in2 => \N__44009\,
            in3 => \N__40122\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44034\,
            in2 => \N__43979\,
            in3 => \N__40119\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43946\,
            in2 => \N__44010\,
            in3 => \N__40116\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43916\,
            in2 => \N__43980\,
            in3 => \N__40113\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43886\,
            in2 => \N__43950\,
            in3 => \N__40110\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17\,
            clk => \N__49815\,
            ce => \N__46409\,
            sr => \N__49392\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43853\,
            in2 => \N__43920\,
            in3 => \N__40275\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_19\,
            ltout => OPEN,
            carryin => \bfn_16_21_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43829\,
            in2 => \N__43890\,
            in3 => \N__40272\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43854\,
            in2 => \N__44288\,
            in3 => \N__40269\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43830\,
            in2 => \N__44258\,
            in3 => \N__40266\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44228\,
            in2 => \N__44289\,
            in3 => \N__40224\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44201\,
            in2 => \N__44259\,
            in3 => \N__40182\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44229\,
            in2 => \N__44174\,
            in3 => \N__40179\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44138\,
            in2 => \N__44205\,
            in3 => \N__40176\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25\,
            clk => \N__49813\,
            ce => \N__46408\,
            sr => \N__49396\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44102\,
            in2 => \N__44175\,
            in3 => \N__40173\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_27\,
            ltout => OPEN,
            carryin => \bfn_16_22_0_\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            clk => \N__49811\,
            ce => \N__46407\,
            sr => \N__49399\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44075\,
            in2 => \N__44142\,
            in3 => \N__40359\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            clk => \N__49811\,
            ce => \N__46407\,
            sr => \N__49399\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44052\,
            in2 => \N__44106\,
            in3 => \N__40356\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            clk => \N__49811\,
            ce => \N__46407\,
            sr => \N__49399\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44076\,
            in2 => \N__44736\,
            in3 => \N__40353\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28\,
            carryout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29\,
            clk => \N__49811\,
            ce => \N__46407\,
            sr => \N__49399\
        );

    \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40350\,
            lcout => \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42598\,
            in1 => \N__48647\,
            in2 => \_gnd_net_\,
            in3 => \N__42136\,
            lcout => \current_shift_inst.un10_control_input_cry_19_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42896\,
            in1 => \N__48184\,
            in2 => \_gnd_net_\,
            in3 => \N__42420\,
            lcout => \current_shift_inst.un10_control_input_cry_27_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48646\,
            in1 => \N__43150\,
            in2 => \_gnd_net_\,
            in3 => \N__42175\,
            lcout => \current_shift_inst.un10_control_input_cry_18_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__40324\,
            in1 => \N__48648\,
            in2 => \_gnd_net_\,
            in3 => \N__42089\,
            lcout => \current_shift_inst.un10_control_input_cry_21_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__42940\,
            in1 => \N__48183\,
            in2 => \_gnd_net_\,
            in3 => \N__42459\,
            lcout => \current_shift_inst.un10_control_input_cry_26_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48645\,
            in1 => \N__40552\,
            in2 => \_gnd_net_\,
            in3 => \N__42212\,
            lcout => \current_shift_inst.un10_control_input_cry_17_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48182\,
            in2 => \_gnd_net_\,
            in3 => \N__42314\,
            lcout => \current_shift_inst.un10_control_input_cry_30_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48179\,
            in1 => \N__43201\,
            in2 => \_gnd_net_\,
            in3 => \N__42656\,
            lcout => \current_shift_inst.un10_control_input_cry_25_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48180\,
            in1 => \N__42997\,
            in2 => \_gnd_net_\,
            in3 => \N__42388\,
            lcout => \current_shift_inst.un10_control_input_cry_28_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__43519\,
            in1 => \N__48181\,
            in2 => \_gnd_net_\,
            in3 => \N__42354\,
            lcout => \current_shift_inst.un10_control_input_cry_29_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_24_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40479\,
            in1 => \N__47047\,
            in2 => \_gnd_net_\,
            in3 => \N__40440\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49943\,
            ce => \N__47160\,
            sr => \N__49294\
        );

    \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0_0_c_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40425\,
            in2 => \N__40419\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_2_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41211\,
            in1 => \N__40398\,
            in2 => \_gnd_net_\,
            in3 => \N__40386\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_2\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_0\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_3_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__41263\,
            in1 => \N__40374\,
            in2 => \N__40383\,
            in3 => \N__40362\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_3\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_1\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_4_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41212\,
            in1 => \N__40683\,
            in2 => \_gnd_net_\,
            in3 => \N__40671\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_4\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_2\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_5_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41264\,
            in1 => \N__40668\,
            in2 => \_gnd_net_\,
            in3 => \N__40656\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_5\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_3\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_6_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41213\,
            in1 => \N__40653\,
            in2 => \_gnd_net_\,
            in3 => \N__40641\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_4\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_7_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41265\,
            in1 => \N__40638\,
            in2 => \_gnd_net_\,
            in3 => \N__40626\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_5\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_8_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41214\,
            in1 => \N__40623\,
            in2 => \_gnd_net_\,
            in3 => \N__40611\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_8\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_6\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_7\,
            clk => \N__49933\,
            ce => 'H',
            sr => \N__49299\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_9_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41253\,
            in1 => \N__40608\,
            in2 => \_gnd_net_\,
            in3 => \N__40596\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_8_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_10_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41242\,
            in1 => \N__40593\,
            in2 => \_gnd_net_\,
            in3 => \N__40581\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_8\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_11_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41250\,
            in1 => \N__40578\,
            in2 => \_gnd_net_\,
            in3 => \N__40566\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_9\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_12_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41243\,
            in1 => \N__40803\,
            in2 => \_gnd_net_\,
            in3 => \N__40791\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_10\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_13_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41251\,
            in1 => \N__40788\,
            in2 => \_gnd_net_\,
            in3 => \N__40776\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_11\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_14_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41244\,
            in1 => \N__40773\,
            in2 => \_gnd_net_\,
            in3 => \N__40761\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_12\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_15_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41252\,
            in1 => \N__40758\,
            in2 => \_gnd_net_\,
            in3 => \N__40746\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_13\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_16_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41245\,
            in1 => \N__44477\,
            in2 => \_gnd_net_\,
            in3 => \N__40743\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_14\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_15\,
            clk => \N__49921\,
            ce => 'H',
            sr => \N__49307\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_17_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41246\,
            in1 => \N__44459\,
            in2 => \_gnd_net_\,
            in3 => \N__40740\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_18_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41276\,
            in1 => \N__40727\,
            in2 => \_gnd_net_\,
            in3 => \N__40713\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_16\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_19_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41247\,
            in1 => \N__40703\,
            in2 => \_gnd_net_\,
            in3 => \N__40689\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_19\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_17\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_20_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41277\,
            in1 => \N__45546\,
            in2 => \_gnd_net_\,
            in3 => \N__40686\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_18\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_21_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41248\,
            in1 => \N__45563\,
            in2 => \_gnd_net_\,
            in3 => \N__40869\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_19\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_22_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41278\,
            in1 => \N__41056\,
            in2 => \_gnd_net_\,
            in3 => \N__40866\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_20\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_23_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41249\,
            in1 => \N__41077\,
            in2 => \_gnd_net_\,
            in3 => \N__40863\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_21\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_24_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41279\,
            in1 => \N__45066\,
            in2 => \_gnd_net_\,
            in3 => \N__40860\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_24\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_22\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_23\,
            clk => \N__49910\,
            ce => 'H',
            sr => \N__49314\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_25_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41269\,
            in1 => \N__45083\,
            in2 => \_gnd_net_\,
            in3 => \N__40857\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_26_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41273\,
            in1 => \N__44948\,
            in2 => \_gnd_net_\,
            in3 => \N__40854\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_24\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_27_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41270\,
            in1 => \N__44916\,
            in2 => \_gnd_net_\,
            in3 => \N__40851\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_25\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_28_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41274\,
            in1 => \N__40846\,
            in2 => \_gnd_net_\,
            in3 => \N__40830\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_28\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_26\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_29_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41271\,
            in1 => \N__40822\,
            in2 => \_gnd_net_\,
            in3 => \N__40806\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_29\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_27\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_30_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41275\,
            in1 => \N__41308\,
            in2 => \_gnd_net_\,
            in3 => \N__41289\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_30\,
            ltout => OPEN,
            carryin => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_28\,
            carryout => \phase_controller_inst2.stoper_hc.un1_accumulated_time_cry_29\,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.accumulated_time_31_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__41272\,
            in1 => \N__41119\,
            in2 => \_gnd_net_\,
            in3 => \N__41130\,
            lcout => \phase_controller_inst2.stoper_hc.accumulated_timeZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49899\,
            ce => 'H',
            sr => \N__49321\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_22_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000100"
        )
    port map (
            in0 => \N__41057\,
            in1 => \N__41640\,
            in2 => \N__41082\,
            in3 => \N__41526\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_22_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__41639\,
            in1 => \N__41081\,
            in2 => \N__41061\,
            in3 => \N__41525\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_10_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41028\,
            in1 => \N__40987\,
            in2 => \_gnd_net_\,
            in3 => \N__47021\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49886\,
            ce => \N__47155\,
            sr => \N__49330\
        );

    \phase_controller_inst2.stoper_hc.target_time_11_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47020\,
            in1 => \N__40947\,
            in2 => \_gnd_net_\,
            in3 => \N__40929\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49886\,
            ce => \N__47155\,
            sr => \N__49330\
        );

    \phase_controller_inst2.stoper_hc.target_time_12_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41367\,
            in1 => \N__41342\,
            in2 => \_gnd_net_\,
            in3 => \N__47022\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49886\,
            ce => \N__47155\,
            sr => \N__49330\
        );

    \phase_controller_inst2.stoper_hc.target_time_9_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47024\,
            in1 => \N__41395\,
            in2 => \_gnd_net_\,
            in3 => \N__41431\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => \N__47154\,
            sr => \N__49338\
        );

    \phase_controller_inst2.stoper_hc.target_time_22_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41678\,
            in1 => \N__47025\,
            in2 => \_gnd_net_\,
            in3 => \N__41655\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => \N__47154\,
            sr => \N__49338\
        );

    \phase_controller_inst2.stoper_hc.target_time_26_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47023\,
            in1 => \N__41623\,
            in2 => \_gnd_net_\,
            in3 => \N__41604\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => \N__47154\,
            sr => \N__49338\
        );

    \phase_controller_inst2.stoper_hc.target_time_23_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41586\,
            in1 => \N__41551\,
            in2 => \_gnd_net_\,
            in3 => \N__47026\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49876\,
            ce => \N__47154\,
            sr => \N__49338\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__46874\,
            in1 => \N__41461\,
            in2 => \_gnd_net_\,
            in3 => \N__41513\,
            lcout => \elapsed_time_ns_1_RNIF13T9_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__46464\,
            in1 => \N__48086\,
            in2 => \_gnd_net_\,
            in3 => \N__41892\,
            lcout => \current_shift_inst.un38_control_input_cry_0_s0_sf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44347\,
            in1 => \N__44320\,
            in2 => \_gnd_net_\,
            in3 => \N__46875\,
            lcout => \elapsed_time_ns_1_RNI02CN9_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45139\,
            in1 => \N__46880\,
            in2 => \_gnd_net_\,
            in3 => \N__50324\,
            lcout => \elapsed_time_ns_1_RNIDV2T9_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__41430\,
            in1 => \_gnd_net_\,
            in2 => \N__46991\,
            in3 => \N__41396\,
            lcout => \elapsed_time_ns_1_RNIL73T9_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__41341\,
            in1 => \N__41374\,
            in2 => \_gnd_net_\,
            in3 => \N__46879\,
            lcout => \elapsed_time_ns_1_RNIV0CN9_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46577\,
            lcout => \current_shift_inst.un4_control_input1_1\,
            ltout => \current_shift_inst.un4_control_input1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48008\,
            in2 => \N__41886\,
            in3 => \N__46460\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__48507\,
            in1 => \N__48524\,
            in2 => \N__46376\,
            in3 => \N__48009\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNITDHV_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48010\,
            in1 => \N__41838\,
            in2 => \N__47876\,
            in3 => \N__41718\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46383\,
            in2 => \N__46578\,
            in3 => \N__46576\,
            lcout => \current_shift_inst.un4_control_input1_2\,
            ltout => OPEN,
            carryin => \bfn_17_15_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41787\,
            in2 => \_gnd_net_\,
            in3 => \N__41754\,
            lcout => \current_shift_inst.un4_control_input1_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_1\,
            carryout => \current_shift_inst.un4_control_input_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42828\,
            in2 => \_gnd_net_\,
            in3 => \N__41727\,
            lcout => \current_shift_inst.un4_control_input1_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_2\,
            carryout => \current_shift_inst.un4_control_input_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41724\,
            in2 => \_gnd_net_\,
            in3 => \N__41703\,
            lcout => \current_shift_inst.un4_control_input1_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_3\,
            carryout => \current_shift_inst.un4_control_input_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42786\,
            in2 => \_gnd_net_\,
            in3 => \N__42057\,
            lcout => \current_shift_inst.un4_control_input1_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_4\,
            carryout => \current_shift_inst.un4_control_input_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42723\,
            in2 => \_gnd_net_\,
            in3 => \N__42024\,
            lcout => \current_shift_inst.un4_control_input1_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_5\,
            carryout => \current_shift_inst.un4_control_input_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42021\,
            in2 => \_gnd_net_\,
            in3 => \N__41979\,
            lcout => \current_shift_inst.un4_control_input1_8\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_6\,
            carryout => \current_shift_inst.un4_control_input_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42669\,
            in2 => \_gnd_net_\,
            in3 => \N__41952\,
            lcout => \current_shift_inst.un4_control_input1_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_7\,
            carryout => \current_shift_inst.un4_control_input_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41949\,
            in2 => \_gnd_net_\,
            in3 => \N__41919\,
            lcout => \current_shift_inst.un4_control_input1_10\,
            ltout => OPEN,
            carryin => \bfn_17_16_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41916\,
            in2 => \_gnd_net_\,
            in3 => \N__41910\,
            lcout => \current_shift_inst.un4_control_input1_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_9\,
            carryout => \current_shift_inst.un4_control_input_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41907\,
            in2 => \_gnd_net_\,
            in3 => \N__41901\,
            lcout => \current_shift_inst.un4_control_input1_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_10\,
            carryout => \current_shift_inst.un4_control_input_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42768\,
            in2 => \_gnd_net_\,
            in3 => \N__41898\,
            lcout => \current_shift_inst.un4_control_input1_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_11\,
            carryout => \current_shift_inst.un4_control_input_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42777\,
            in2 => \_gnd_net_\,
            in3 => \N__41895\,
            lcout => \current_shift_inst.un4_control_input1_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_12\,
            carryout => \current_shift_inst.un4_control_input_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43269\,
            in2 => \_gnd_net_\,
            in3 => \N__42282\,
            lcout => \current_shift_inst.un4_control_input1_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_13\,
            carryout => \current_shift_inst.un4_control_input_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43074\,
            in2 => \_gnd_net_\,
            in3 => \N__42252\,
            lcout => \current_shift_inst.un4_control_input1_16\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_14\,
            carryout => \current_shift_inst.un4_control_input_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43218\,
            in2 => \_gnd_net_\,
            in3 => \N__42222\,
            lcout => \current_shift_inst.un4_control_input1_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_15\,
            carryout => \current_shift_inst.un4_control_input_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42219\,
            in2 => \_gnd_net_\,
            in3 => \N__42183\,
            lcout => \current_shift_inst.un4_control_input1_18\,
            ltout => OPEN,
            carryin => \bfn_17_17_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_17\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43122\,
            in3 => \N__42144\,
            lcout => \current_shift_inst.un4_control_input1_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_17\,
            carryout => \current_shift_inst.un4_control_input_1_cry_18\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42573\,
            in2 => \_gnd_net_\,
            in3 => \N__42105\,
            lcout => \current_shift_inst.un4_control_input1_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_18\,
            carryout => \current_shift_inst.un4_control_input_1_cry_19\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43542\,
            in2 => \_gnd_net_\,
            in3 => \N__42102\,
            lcout => \current_shift_inst.un4_control_input1_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_19\,
            carryout => \current_shift_inst.un4_control_input_1_cry_20\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42099\,
            in2 => \_gnd_net_\,
            in3 => \N__42060\,
            lcout => \current_shift_inst.un4_control_input1_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_20\,
            carryout => \current_shift_inst.un4_control_input_1_cry_21\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42564\,
            in2 => \_gnd_net_\,
            in3 => \N__42534\,
            lcout => \current_shift_inst.un4_control_input1_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_21\,
            carryout => \current_shift_inst.un4_control_input_1_cry_22\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42531\,
            in2 => \_gnd_net_\,
            in3 => \N__42492\,
            lcout => \current_shift_inst.un4_control_input1_24\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_22\,
            carryout => \current_shift_inst.un4_control_input_1_cry_23\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43023\,
            in2 => \_gnd_net_\,
            in3 => \N__42465\,
            lcout => \current_shift_inst.un4_control_input1_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_23\,
            carryout => \current_shift_inst.un4_control_input_1_cry_24\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43173\,
            in2 => \_gnd_net_\,
            in3 => \N__42462\,
            lcout => \current_shift_inst.un4_control_input1_26\,
            ltout => OPEN,
            carryin => \bfn_17_18_0_\,
            carryout => \current_shift_inst.un4_control_input_1_cry_25\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42921\,
            in2 => \_gnd_net_\,
            in3 => \N__42423\,
            lcout => \current_shift_inst.un4_control_input1_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_25\,
            carryout => \current_shift_inst.un4_control_input_1_cry_26\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42879\,
            in2 => \_gnd_net_\,
            in3 => \N__42393\,
            lcout => \current_shift_inst.un4_control_input1_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_26\,
            carryout => \current_shift_inst.un4_control_input_1_cry_27\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42969\,
            in2 => \_gnd_net_\,
            in3 => \N__42357\,
            lcout => \current_shift_inst.un4_control_input1_29\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_27\,
            carryout => \current_shift_inst.un4_control_input_1_cry_28\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43494\,
            in2 => \_gnd_net_\,
            in3 => \N__42324\,
            lcout => \current_shift_inst.un4_control_input1_30\,
            ltout => OPEN,
            carryin => \current_shift_inst.un4_control_input_1_cry_28\,
            carryout => \current_shift_inst.un4_control_input1_31\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42321\,
            lcout => \current_shift_inst.un4_control_input1_31_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__42844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \current_shift_inst.un4_control_input_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42799\,
            lcout => \current_shift_inst.un4_control_input_1_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47901\,
            lcout => \current_shift_inst.un4_control_input_1_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48450\,
            lcout => \current_shift_inst.un4_control_input_1_axb_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42738\,
            lcout => \current_shift_inst.un4_control_input_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42687\,
            lcout => \current_shift_inst.un4_control_input_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__48254\,
            in1 => \N__42640\,
            in2 => \N__47880\,
            in3 => \N__43205\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNISV131_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42589\,
            lcout => \current_shift_inst.un4_control_input_1_axb_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43470\,
            lcout => \current_shift_inst.un4_control_input_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43239\,
            lcout => \current_shift_inst.un4_control_input_1_axb_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43191\,
            lcout => \current_shift_inst.un4_control_input_1_axb_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43140\,
            lcout => \current_shift_inst.un4_control_input_1_axb_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43092\,
            lcout => \current_shift_inst.un4_control_input_1_axb_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43039\,
            lcout => \current_shift_inst.un4_control_input_1_axb_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42987\,
            lcout => \current_shift_inst.un4_control_input_1_axb_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42939\,
            lcout => \current_shift_inst.un4_control_input_1_axb_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__42895\,
            lcout => \current_shift_inst.un4_control_input_1_axb_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48304\,
            lcout => \current_shift_inst.un4_control_input_1_axb_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_17_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43510\,
            lcout => \current_shift_inst.un4_control_input_1_axb_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48643\,
            in1 => \N__43480\,
            in2 => \_gnd_net_\,
            in3 => \N__43441\,
            lcout => \current_shift_inst.un10_control_input_cry_14_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__47911\,
            in1 => \N__48642\,
            in2 => \_gnd_net_\,
            in3 => \N__47277\,
            lcout => \current_shift_inst.un10_control_input_cry_13_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48641\,
            in1 => \N__43375\,
            in2 => \_gnd_net_\,
            in3 => \N__43336\,
            lcout => \current_shift_inst.un10_control_input_cry_11_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.counter_0_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44867\,
            in1 => \N__46483\,
            in2 => \_gnd_net_\,
            in3 => \N__43305\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_23_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_0\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_1_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44818\,
            in1 => \N__46432\,
            in2 => \_gnd_net_\,
            in3 => \N__43302\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_0\,
            carryout => \current_shift_inst.timer_s1.counter_cry_1\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_2_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44868\,
            in1 => \N__43288\,
            in2 => \_gnd_net_\,
            in3 => \N__43272\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_1\,
            carryout => \current_shift_inst.timer_s1.counter_cry_2\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_3_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44819\,
            in1 => \N__43793\,
            in2 => \_gnd_net_\,
            in3 => \N__43779\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_2\,
            carryout => \current_shift_inst.timer_s1.counter_cry_3\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_4_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44869\,
            in1 => \N__43763\,
            in2 => \_gnd_net_\,
            in3 => \N__43749\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_3\,
            carryout => \current_shift_inst.timer_s1.counter_cry_4\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_5_LC_17_23_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44820\,
            in1 => \N__43735\,
            in2 => \_gnd_net_\,
            in3 => \N__43719\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_4\,
            carryout => \current_shift_inst.timer_s1.counter_cry_5\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_6_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44870\,
            in1 => \N__43709\,
            in2 => \_gnd_net_\,
            in3 => \N__43695\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_5\,
            carryout => \current_shift_inst.timer_s1.counter_cry_6\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_7_LC_17_23_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44821\,
            in1 => \N__43685\,
            in2 => \_gnd_net_\,
            in3 => \N__43671\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_6\,
            carryout => \current_shift_inst.timer_s1.counter_cry_7\,
            clk => \N__49812\,
            ce => \N__44714\,
            sr => \N__49400\
        );

    \current_shift_inst.timer_s1.counter_8_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44849\,
            in1 => \N__43654\,
            in2 => \_gnd_net_\,
            in3 => \N__43638\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_17_24_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_8\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_9_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44853\,
            in1 => \N__43618\,
            in2 => \_gnd_net_\,
            in3 => \N__43599\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_8\,
            carryout => \current_shift_inst.timer_s1.counter_cry_9\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_10_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44846\,
            in1 => \N__43585\,
            in2 => \_gnd_net_\,
            in3 => \N__43569\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_9\,
            carryout => \current_shift_inst.timer_s1.counter_cry_10\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_11_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44850\,
            in1 => \N__43559\,
            in2 => \_gnd_net_\,
            in3 => \N__43545\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_10\,
            carryout => \current_shift_inst.timer_s1.counter_cry_11\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_12_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44847\,
            in1 => \N__44027\,
            in2 => \_gnd_net_\,
            in3 => \N__44013\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_11\,
            carryout => \current_shift_inst.timer_s1.counter_cry_12\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_13_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44851\,
            in1 => \N__43997\,
            in2 => \_gnd_net_\,
            in3 => \N__43983\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_12\,
            carryout => \current_shift_inst.timer_s1.counter_cry_13\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_14_LC_17_24_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44848\,
            in1 => \N__43967\,
            in2 => \_gnd_net_\,
            in3 => \N__43953\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_13\,
            carryout => \current_shift_inst.timer_s1.counter_cry_14\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_15_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44852\,
            in1 => \N__43939\,
            in2 => \_gnd_net_\,
            in3 => \N__43923\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_14\,
            carryout => \current_shift_inst.timer_s1.counter_cry_15\,
            clk => \N__49810\,
            ce => \N__44706\,
            sr => \N__49406\
        );

    \current_shift_inst.timer_s1.counter_16_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44863\,
            in1 => \N__43909\,
            in2 => \_gnd_net_\,
            in3 => \N__43893\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_17_25_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_16\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_17_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44871\,
            in1 => \N__43879\,
            in2 => \_gnd_net_\,
            in3 => \N__43857\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_16\,
            carryout => \current_shift_inst.timer_s1.counter_cry_17\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_18_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44864\,
            in1 => \N__43847\,
            in2 => \_gnd_net_\,
            in3 => \N__43833\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_17\,
            carryout => \current_shift_inst.timer_s1.counter_cry_18\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_19_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44872\,
            in1 => \N__43823\,
            in2 => \_gnd_net_\,
            in3 => \N__43809\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_18\,
            carryout => \current_shift_inst.timer_s1.counter_cry_19\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_20_LC_17_25_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44865\,
            in1 => \N__44276\,
            in2 => \_gnd_net_\,
            in3 => \N__44262\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_19\,
            carryout => \current_shift_inst.timer_s1.counter_cry_20\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_21_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44873\,
            in1 => \N__44246\,
            in2 => \_gnd_net_\,
            in3 => \N__44232\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_20\,
            carryout => \current_shift_inst.timer_s1.counter_cry_21\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_22_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44866\,
            in1 => \N__44222\,
            in2 => \_gnd_net_\,
            in3 => \N__44208\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_21\,
            carryout => \current_shift_inst.timer_s1.counter_cry_22\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_23_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44874\,
            in1 => \N__44194\,
            in2 => \_gnd_net_\,
            in3 => \N__44178\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_22\,
            carryout => \current_shift_inst.timer_s1.counter_cry_23\,
            clk => \N__49807\,
            ce => \N__44715\,
            sr => \N__49409\
        );

    \current_shift_inst.timer_s1.counter_24_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44822\,
            in1 => \N__44161\,
            in2 => \_gnd_net_\,
            in3 => \N__44145\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_17_26_0_\,
            carryout => \current_shift_inst.timer_s1.counter_cry_24\,
            clk => \N__49804\,
            ce => \N__44713\,
            sr => \N__49413\
        );

    \current_shift_inst.timer_s1.counter_25_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44826\,
            in1 => \N__44131\,
            in2 => \_gnd_net_\,
            in3 => \N__44109\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_24\,
            carryout => \current_shift_inst.timer_s1.counter_cry_25\,
            clk => \N__49804\,
            ce => \N__44713\,
            sr => \N__49413\
        );

    \current_shift_inst.timer_s1.counter_26_LC_17_26_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44823\,
            in1 => \N__44095\,
            in2 => \_gnd_net_\,
            in3 => \N__44079\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_25\,
            carryout => \current_shift_inst.timer_s1.counter_cry_26\,
            clk => \N__49804\,
            ce => \N__44713\,
            sr => \N__49413\
        );

    \current_shift_inst.timer_s1.counter_27_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44827\,
            in1 => \N__44069\,
            in2 => \_gnd_net_\,
            in3 => \N__44055\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_26\,
            carryout => \current_shift_inst.timer_s1.counter_cry_27\,
            clk => \N__49804\,
            ce => \N__44713\,
            sr => \N__49413\
        );

    \current_shift_inst.timer_s1.counter_28_LC_17_26_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__44824\,
            in1 => \N__44048\,
            in2 => \_gnd_net_\,
            in3 => \N__44877\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \current_shift_inst.timer_s1.counter_cry_27\,
            carryout => \current_shift_inst.timer_s1.counter_cry_28\,
            clk => \N__49804\,
            ce => \N__44713\,
            sr => \N__49413\
        );

    \current_shift_inst.timer_s1.counter_29_LC_17_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__44729\,
            in1 => \N__44825\,
            in2 => \_gnd_net_\,
            in3 => \N__44739\,
            lcout => \current_shift_inst.timer_s1.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49804\,
            ce => \N__44713\,
            sr => \N__49413\
        );

    \phase_controller_inst2.stoper_hc.target_time_20_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47040\,
            in1 => \N__44667\,
            in2 => \_gnd_net_\,
            in3 => \N__44631\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => \N__47161\,
            sr => \N__49295\
        );

    \phase_controller_inst2.stoper_hc.target_time_17_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44613\,
            in1 => \N__44588\,
            in2 => \_gnd_net_\,
            in3 => \N__47042\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => \N__47161\,
            sr => \N__49295\
        );

    \phase_controller_inst2.stoper_hc.target_time_14_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44547\,
            in1 => \N__44517\,
            in2 => \_gnd_net_\,
            in3 => \N__47041\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49944\,
            ce => \N__47161\,
            sr => \N__49295\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_16_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010101110"
        )
    port map (
            in0 => \N__44442\,
            in1 => \N__44364\,
            in2 => \N__44478\,
            in3 => \N__44458\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_16_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100001011"
        )
    port map (
            in0 => \N__44363\,
            in1 => \N__44476\,
            in2 => \N__44460\,
            in3 => \N__44441\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_16_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44418\,
            in1 => \N__47044\,
            in2 => \_gnd_net_\,
            in3 => \N__44382\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => \N__47159\,
            sr => \N__49300\
        );

    \phase_controller_inst2.stoper_hc.target_time_13_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44355\,
            in1 => \N__44325\,
            in2 => \_gnd_net_\,
            in3 => \N__47045\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => \N__47159\,
            sr => \N__49300\
        );

    \phase_controller_inst2.stoper_hc.target_time_15_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45216\,
            in1 => \N__45192\,
            in2 => \_gnd_net_\,
            in3 => \N__47046\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => \N__47159\,
            sr => \N__49300\
        );

    \phase_controller_inst2.stoper_hc.target_time_1_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47043\,
            in1 => \N__45147\,
            in2 => \_gnd_net_\,
            in3 => \N__50323\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49934\,
            ce => \N__47159\,
            sr => \N__49300\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_24_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__45065\,
            in1 => \N__45096\,
            in2 => \N__44973\,
            in3 => \N__45082\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_24_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__45095\,
            in1 => \N__44972\,
            in2 => \N__45084\,
            in3 => \N__45064\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_25_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__45039\,
            in1 => \N__45013\,
            in2 => \_gnd_net_\,
            in3 => \N__47032\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49922\,
            ce => \N__47158\,
            sr => \N__49308\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_26_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100100011"
        )
    port map (
            in0 => \N__44927\,
            in1 => \N__44914\,
            in2 => \N__44949\,
            in3 => \N__47174\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_26_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__44947\,
            in1 => \N__44928\,
            in2 => \N__47178\,
            in3 => \N__44915\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_0_20_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110100"
        )
    port map (
            in0 => \N__45545\,
            in1 => \N__45576\,
            in2 => \N__45456\,
            in3 => \N__45562\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_lt20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_20_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111011001111"
        )
    port map (
            in0 => \N__45575\,
            in1 => \N__45455\,
            in2 => \N__45564\,
            in3 => \N__45544\,
            lcout => \phase_controller_inst2.stoper_hc.un4_running_cry_c_RNO_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_21_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45515\,
            in1 => \N__47056\,
            in2 => \_gnd_net_\,
            in3 => \N__45474\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49911\,
            ce => \N__47157\,
            sr => \N__49315\
        );

    \phase_controller_inst2.stoper_hc.target_time_6_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__47055\,
            in1 => \N__45441\,
            in2 => \_gnd_net_\,
            in3 => \N__45414\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49911\,
            ce => \N__47157\,
            sr => \N__49315\
        );

    \phase_controller_inst2.stoper_hc.target_time_7_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45384\,
            in1 => \N__47057\,
            in2 => \_gnd_net_\,
            in3 => \N__45352\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49911\,
            ce => \N__47157\,
            sr => \N__49315\
        );

    \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50177\,
            in1 => \N__50344\,
            in2 => \_gnd_net_\,
            in3 => \N__45309\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_18_11_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50173\,
            in1 => \N__45295\,
            in2 => \_gnd_net_\,
            in3 => \N__45276\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_0\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50178\,
            in1 => \N__45266\,
            in2 => \_gnd_net_\,
            in3 => \N__45252\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_1\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50174\,
            in1 => \N__45242\,
            in2 => \_gnd_net_\,
            in3 => \N__45228\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_2\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50179\,
            in1 => \N__45803\,
            in2 => \_gnd_net_\,
            in3 => \N__45789\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_3\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50175\,
            in1 => \N__45773\,
            in2 => \_gnd_net_\,
            in3 => \N__45759\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_4\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50180\,
            in1 => \N__45749\,
            in2 => \_gnd_net_\,
            in3 => \N__45735\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_5\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50176\,
            in1 => \N__45725\,
            in2 => \_gnd_net_\,
            in3 => \N__45711\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_6\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_7\,
            clk => \N__49900\,
            ce => \N__50283\,
            sr => \N__49322\
        );

    \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50166\,
            in1 => \N__45694\,
            in2 => \_gnd_net_\,
            in3 => \N__45672\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50162\,
            in1 => \N__45655\,
            in2 => \_gnd_net_\,
            in3 => \N__45633\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_8\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50163\,
            in1 => \N__45619\,
            in2 => \_gnd_net_\,
            in3 => \N__45603\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_9\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50159\,
            in1 => \N__45593\,
            in2 => \_gnd_net_\,
            in3 => \N__45579\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_10\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50164\,
            in1 => \N__46078\,
            in2 => \_gnd_net_\,
            in3 => \N__46062\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_11\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50160\,
            in1 => \N__46046\,
            in2 => \_gnd_net_\,
            in3 => \N__46032\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_12\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50165\,
            in1 => \N__46018\,
            in2 => \_gnd_net_\,
            in3 => \N__46002\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_13\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50161\,
            in1 => \N__45997\,
            in2 => \_gnd_net_\,
            in3 => \N__45978\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_14\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_15\,
            clk => \N__49887\,
            ce => \N__50278\,
            sr => \N__49331\
        );

    \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50146\,
            in1 => \N__45964\,
            in2 => \_gnd_net_\,
            in3 => \N__45942\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50181\,
            in1 => \N__45925\,
            in2 => \_gnd_net_\,
            in3 => \N__45909\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_16\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50147\,
            in1 => \N__45895\,
            in2 => \_gnd_net_\,
            in3 => \N__45879\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_17\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50182\,
            in1 => \N__45865\,
            in2 => \_gnd_net_\,
            in3 => \N__45849\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_18\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50148\,
            in1 => \N__45835\,
            in2 => \_gnd_net_\,
            in3 => \N__45819\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_19\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50183\,
            in1 => \N__46315\,
            in2 => \_gnd_net_\,
            in3 => \N__46299\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_20\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50149\,
            in1 => \N__46285\,
            in2 => \_gnd_net_\,
            in3 => \N__46269\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_21\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50184\,
            in1 => \N__46259\,
            in2 => \_gnd_net_\,
            in3 => \N__46245\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_22\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_23\,
            clk => \N__49877\,
            ce => \N__50277\,
            sr => \N__49339\
        );

    \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50167\,
            in1 => \N__46237\,
            in2 => \_gnd_net_\,
            in3 => \N__46209\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            clk => \N__49865\,
            ce => \N__50279\,
            sr => \N__49347\
        );

    \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50171\,
            in1 => \N__46192\,
            in2 => \_gnd_net_\,
            in3 => \N__46170\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_24\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            clk => \N__49865\,
            ce => \N__50279\,
            sr => \N__49347\
        );

    \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50168\,
            in1 => \N__46160\,
            in2 => \_gnd_net_\,
            in3 => \N__46146\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_25\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            clk => \N__49865\,
            ce => \N__50279\,
            sr => \N__49347\
        );

    \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50172\,
            in1 => \N__46132\,
            in2 => \_gnd_net_\,
            in3 => \N__46116\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_26\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            clk => \N__49865\,
            ce => \N__50279\,
            sr => \N__49347\
        );

    \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__50169\,
            in1 => \N__46106\,
            in2 => \_gnd_net_\,
            in3 => \N__46092\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \delay_measurement_inst.delay_hc_timer.counter_cry_27\,
            carryout => \delay_measurement_inst.delay_hc_timer.counter_cry_28\,
            clk => \N__49865\,
            ce => \N__50279\,
            sr => \N__49347\
        );

    \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__46604\,
            in1 => \N__50170\,
            in2 => \_gnd_net_\,
            in3 => \N__46611\,
            lcout => \delay_measurement_inst.delay_hc_timer.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49865\,
            ce => \N__50279\,
            sr => \N__49347\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48206\,
            in2 => \_gnd_net_\,
            in3 => \N__47768\,
            lcout => \current_shift_inst.un38_control_input_axb_31_s0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46458\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_i_1\,
            ltout => \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__46459\,
            in1 => \_gnd_net_\,
            in2 => \N__46557\,
            in3 => \N__48550\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNINRRH_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46530\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_31_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => \N__46413\,
            sr => \N__49357\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46494\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49854\,
            ce => \N__46413\,
            sr => \N__49357\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46440\,
            lcout => \current_shift_inst.elapsed_time_ns_s1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49842\,
            ce => \N__46412\,
            sr => \N__49364\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48501\,
            lcout => \current_shift_inst.un4_control_input_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__48503\,
            in1 => \N__48205\,
            in2 => \N__46377\,
            in3 => \N__48525\,
            lcout => \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__48551\,
            in1 => \N__48523\,
            in2 => \_gnd_net_\,
            in3 => \N__48502\,
            lcout => \current_shift_inst.un10_control_input_cry_1_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48239\,
            in1 => \N__48468\,
            in2 => \N__47865\,
            in3 => \N__48425\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48238\,
            in1 => \N__48392\,
            in2 => \N__47864\,
            in3 => \N__48353\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__48241\,
            in1 => \N__47791\,
            in2 => \N__48321\,
            in3 => \N__48287\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__48240\,
            in1 => \N__47919\,
            in2 => \N__47866\,
            in3 => \N__47273\,
            lcout => \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \phase_controller_inst2.stoper_hc.target_time_18_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__47244\,
            in1 => \N__47069\,
            in2 => \_gnd_net_\,
            in3 => \N__47211\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49949\,
            ce => \N__47163\,
            sr => \N__49301\
        );

    \phase_controller_inst2.stoper_hc.target_time_27_LC_20_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__47120\,
            in1 => \N__50371\,
            in2 => \_gnd_net_\,
            in3 => \N__47070\,
            lcout => \phase_controller_inst2.stoper_hc.target_timeZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49945\,
            ce => \N__47162\,
            sr => \N__49309\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50375\,
            in1 => \N__47113\,
            in2 => \_gnd_net_\,
            in3 => \N__47048\,
            lcout => \elapsed_time_ns_1_RNI58DN9_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50351\,
            lcout => \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49923\,
            ce => \N__50214\,
            sr => \N__49323\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__49972\,
            in1 => \_gnd_net_\,
            in2 => \N__50042\,
            in3 => \N__50006\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_164_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49973\,
            in2 => \_gnd_net_\,
            in3 => \N__50035\,
            lcout => \delay_measurement_inst.delay_hc_timer.N_163_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49971\,
            lcout => \delay_measurement_inst.delay_hc_timer.running_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_measurement_inst.delay_hc_timer.running_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__49974\,
            in1 => \N__50043\,
            in2 => \_gnd_net_\,
            in3 => \N__50010\,
            lcout => \delay_measurement_inst.delay_hc_timer.runningZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__49889\,
            ce => 'H',
            sr => \N__49348\
        );

    \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofx_LC_24_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__48954\,
            in1 => \N__48881\,
            in2 => \_gnd_net_\,
            in3 => \N__48868\,
            lcout => \pwm_generator_inst.un2_threshold_add_1_axb_15_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
