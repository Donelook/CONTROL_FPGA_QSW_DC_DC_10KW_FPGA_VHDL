// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Sep 25 2024 17:56:48

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "MAIN" view "INTERFACE"

module MAIN (
    s3_phy,
    il_min_comp2,
    il_max_comp1,
    error_pin,
    s1_phy,
    reset,
    il_min_comp1,
    delay_tr_input,
    s4_phy,
    start_stop,
    s2_phy,
    pwm_output,
    il_max_comp2,
    delay_hc_input);

    output s3_phy;
    input il_min_comp2;
    input il_max_comp1;
    input error_pin;
    output s1_phy;
    input reset;
    input il_min_comp1;
    input delay_tr_input;
    output s4_phy;
    input start_stop;
    output s2_phy;
    output pwm_output;
    input il_max_comp2;
    input delay_hc_input;

    wire N__53311;
    wire N__53310;
    wire N__53309;
    wire N__53300;
    wire N__53299;
    wire N__53298;
    wire N__53291;
    wire N__53290;
    wire N__53289;
    wire N__53282;
    wire N__53281;
    wire N__53280;
    wire N__53273;
    wire N__53272;
    wire N__53271;
    wire N__53264;
    wire N__53263;
    wire N__53262;
    wire N__53255;
    wire N__53254;
    wire N__53253;
    wire N__53246;
    wire N__53245;
    wire N__53244;
    wire N__53237;
    wire N__53236;
    wire N__53235;
    wire N__53228;
    wire N__53227;
    wire N__53226;
    wire N__53219;
    wire N__53218;
    wire N__53217;
    wire N__53210;
    wire N__53209;
    wire N__53208;
    wire N__53201;
    wire N__53200;
    wire N__53199;
    wire N__53182;
    wire N__53179;
    wire N__53176;
    wire N__53175;
    wire N__53172;
    wire N__53169;
    wire N__53168;
    wire N__53163;
    wire N__53160;
    wire N__53155;
    wire N__53152;
    wire N__53149;
    wire N__53146;
    wire N__53143;
    wire N__53140;
    wire N__53137;
    wire N__53134;
    wire N__53131;
    wire N__53128;
    wire N__53125;
    wire N__53124;
    wire N__53121;
    wire N__53118;
    wire N__53113;
    wire N__53112;
    wire N__53111;
    wire N__53108;
    wire N__53105;
    wire N__53104;
    wire N__53099;
    wire N__53096;
    wire N__53093;
    wire N__53090;
    wire N__53085;
    wire N__53082;
    wire N__53079;
    wire N__53076;
    wire N__53073;
    wire N__53070;
    wire N__53067;
    wire N__53062;
    wire N__53059;
    wire N__53056;
    wire N__53053;
    wire N__53052;
    wire N__53051;
    wire N__53048;
    wire N__53045;
    wire N__53042;
    wire N__53039;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53023;
    wire N__53020;
    wire N__53017;
    wire N__53014;
    wire N__53011;
    wire N__53008;
    wire N__53005;
    wire N__53004;
    wire N__53003;
    wire N__52998;
    wire N__52995;
    wire N__52990;
    wire N__52987;
    wire N__52984;
    wire N__52983;
    wire N__52980;
    wire N__52977;
    wire N__52976;
    wire N__52971;
    wire N__52968;
    wire N__52965;
    wire N__52962;
    wire N__52957;
    wire N__52954;
    wire N__52951;
    wire N__52948;
    wire N__52945;
    wire N__52942;
    wire N__52939;
    wire N__52938;
    wire N__52935;
    wire N__52932;
    wire N__52927;
    wire N__52924;
    wire N__52921;
    wire N__52920;
    wire N__52919;
    wire N__52918;
    wire N__52917;
    wire N__52916;
    wire N__52911;
    wire N__52908;
    wire N__52901;
    wire N__52900;
    wire N__52897;
    wire N__52894;
    wire N__52891;
    wire N__52888;
    wire N__52885;
    wire N__52882;
    wire N__52877;
    wire N__52876;
    wire N__52875;
    wire N__52874;
    wire N__52871;
    wire N__52868;
    wire N__52865;
    wire N__52858;
    wire N__52855;
    wire N__52852;
    wire N__52849;
    wire N__52846;
    wire N__52837;
    wire N__52834;
    wire N__52833;
    wire N__52832;
    wire N__52831;
    wire N__52830;
    wire N__52829;
    wire N__52824;
    wire N__52823;
    wire N__52816;
    wire N__52813;
    wire N__52810;
    wire N__52807;
    wire N__52802;
    wire N__52797;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52779;
    wire N__52774;
    wire N__52771;
    wire N__52770;
    wire N__52767;
    wire N__52764;
    wire N__52761;
    wire N__52758;
    wire N__52757;
    wire N__52754;
    wire N__52751;
    wire N__52748;
    wire N__52745;
    wire N__52742;
    wire N__52739;
    wire N__52732;
    wire N__52729;
    wire N__52728;
    wire N__52727;
    wire N__52726;
    wire N__52723;
    wire N__52722;
    wire N__52719;
    wire N__52718;
    wire N__52715;
    wire N__52710;
    wire N__52705;
    wire N__52702;
    wire N__52701;
    wire N__52700;
    wire N__52697;
    wire N__52692;
    wire N__52687;
    wire N__52684;
    wire N__52675;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52657;
    wire N__52656;
    wire N__52655;
    wire N__52654;
    wire N__52653;
    wire N__52652;
    wire N__52651;
    wire N__52650;
    wire N__52649;
    wire N__52648;
    wire N__52647;
    wire N__52646;
    wire N__52645;
    wire N__52644;
    wire N__52643;
    wire N__52642;
    wire N__52641;
    wire N__52640;
    wire N__52639;
    wire N__52638;
    wire N__52637;
    wire N__52636;
    wire N__52635;
    wire N__52634;
    wire N__52633;
    wire N__52632;
    wire N__52631;
    wire N__52630;
    wire N__52629;
    wire N__52628;
    wire N__52627;
    wire N__52626;
    wire N__52625;
    wire N__52624;
    wire N__52623;
    wire N__52622;
    wire N__52621;
    wire N__52620;
    wire N__52619;
    wire N__52618;
    wire N__52617;
    wire N__52616;
    wire N__52615;
    wire N__52614;
    wire N__52613;
    wire N__52612;
    wire N__52611;
    wire N__52610;
    wire N__52609;
    wire N__52608;
    wire N__52607;
    wire N__52606;
    wire N__52605;
    wire N__52604;
    wire N__52603;
    wire N__52602;
    wire N__52601;
    wire N__52600;
    wire N__52599;
    wire N__52598;
    wire N__52597;
    wire N__52596;
    wire N__52595;
    wire N__52594;
    wire N__52593;
    wire N__52592;
    wire N__52591;
    wire N__52590;
    wire N__52589;
    wire N__52588;
    wire N__52587;
    wire N__52586;
    wire N__52585;
    wire N__52584;
    wire N__52583;
    wire N__52582;
    wire N__52581;
    wire N__52580;
    wire N__52579;
    wire N__52578;
    wire N__52577;
    wire N__52576;
    wire N__52575;
    wire N__52574;
    wire N__52573;
    wire N__52572;
    wire N__52571;
    wire N__52570;
    wire N__52569;
    wire N__52568;
    wire N__52567;
    wire N__52566;
    wire N__52565;
    wire N__52564;
    wire N__52563;
    wire N__52562;
    wire N__52561;
    wire N__52560;
    wire N__52559;
    wire N__52558;
    wire N__52557;
    wire N__52556;
    wire N__52555;
    wire N__52554;
    wire N__52553;
    wire N__52552;
    wire N__52551;
    wire N__52550;
    wire N__52549;
    wire N__52548;
    wire N__52547;
    wire N__52546;
    wire N__52545;
    wire N__52544;
    wire N__52543;
    wire N__52542;
    wire N__52541;
    wire N__52540;
    wire N__52539;
    wire N__52538;
    wire N__52297;
    wire N__52294;
    wire N__52293;
    wire N__52292;
    wire N__52291;
    wire N__52290;
    wire N__52287;
    wire N__52284;
    wire N__52281;
    wire N__52278;
    wire N__52275;
    wire N__52272;
    wire N__52271;
    wire N__52270;
    wire N__52269;
    wire N__52268;
    wire N__52267;
    wire N__52266;
    wire N__52265;
    wire N__52264;
    wire N__52263;
    wire N__52262;
    wire N__52261;
    wire N__52260;
    wire N__52259;
    wire N__52258;
    wire N__52257;
    wire N__52256;
    wire N__52255;
    wire N__52254;
    wire N__52253;
    wire N__52252;
    wire N__52251;
    wire N__52250;
    wire N__52249;
    wire N__52248;
    wire N__52247;
    wire N__52246;
    wire N__52245;
    wire N__52244;
    wire N__52243;
    wire N__52242;
    wire N__52241;
    wire N__52240;
    wire N__52239;
    wire N__52238;
    wire N__52237;
    wire N__52236;
    wire N__52235;
    wire N__52234;
    wire N__52233;
    wire N__52232;
    wire N__52231;
    wire N__52230;
    wire N__52229;
    wire N__52226;
    wire N__52225;
    wire N__52224;
    wire N__52223;
    wire N__52222;
    wire N__52221;
    wire N__52220;
    wire N__52219;
    wire N__52218;
    wire N__52217;
    wire N__52216;
    wire N__52215;
    wire N__52214;
    wire N__52213;
    wire N__52212;
    wire N__52211;
    wire N__52210;
    wire N__52209;
    wire N__52208;
    wire N__52207;
    wire N__52206;
    wire N__52203;
    wire N__52200;
    wire N__52199;
    wire N__52198;
    wire N__52197;
    wire N__52196;
    wire N__52195;
    wire N__52194;
    wire N__52193;
    wire N__52192;
    wire N__52191;
    wire N__52190;
    wire N__52189;
    wire N__52188;
    wire N__52187;
    wire N__52184;
    wire N__52183;
    wire N__52182;
    wire N__52181;
    wire N__52180;
    wire N__52179;
    wire N__52178;
    wire N__52177;
    wire N__52176;
    wire N__52175;
    wire N__52174;
    wire N__52173;
    wire N__52172;
    wire N__52171;
    wire N__52170;
    wire N__52169;
    wire N__52168;
    wire N__51973;
    wire N__51970;
    wire N__51967;
    wire N__51964;
    wire N__51961;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51949;
    wire N__51946;
    wire N__51945;
    wire N__51942;
    wire N__51939;
    wire N__51936;
    wire N__51933;
    wire N__51930;
    wire N__51925;
    wire N__51922;
    wire N__51919;
    wire N__51916;
    wire N__51913;
    wire N__51910;
    wire N__51907;
    wire N__51904;
    wire N__51903;
    wire N__51900;
    wire N__51897;
    wire N__51894;
    wire N__51891;
    wire N__51890;
    wire N__51887;
    wire N__51884;
    wire N__51881;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51865;
    wire N__51862;
    wire N__51859;
    wire N__51858;
    wire N__51857;
    wire N__51856;
    wire N__51855;
    wire N__51854;
    wire N__51853;
    wire N__51852;
    wire N__51851;
    wire N__51850;
    wire N__51849;
    wire N__51848;
    wire N__51847;
    wire N__51846;
    wire N__51845;
    wire N__51844;
    wire N__51827;
    wire N__51810;
    wire N__51805;
    wire N__51802;
    wire N__51801;
    wire N__51800;
    wire N__51799;
    wire N__51798;
    wire N__51797;
    wire N__51794;
    wire N__51789;
    wire N__51782;
    wire N__51779;
    wire N__51774;
    wire N__51769;
    wire N__51766;
    wire N__51763;
    wire N__51760;
    wire N__51757;
    wire N__51754;
    wire N__51751;
    wire N__51748;
    wire N__51745;
    wire N__51742;
    wire N__51739;
    wire N__51736;
    wire N__51733;
    wire N__51730;
    wire N__51727;
    wire N__51724;
    wire N__51721;
    wire N__51718;
    wire N__51715;
    wire N__51712;
    wire N__51711;
    wire N__51708;
    wire N__51705;
    wire N__51704;
    wire N__51701;
    wire N__51698;
    wire N__51695;
    wire N__51688;
    wire N__51685;
    wire N__51682;
    wire N__51679;
    wire N__51676;
    wire N__51673;
    wire N__51670;
    wire N__51667;
    wire N__51664;
    wire N__51661;
    wire N__51660;
    wire N__51659;
    wire N__51656;
    wire N__51653;
    wire N__51650;
    wire N__51649;
    wire N__51648;
    wire N__51647;
    wire N__51646;
    wire N__51645;
    wire N__51644;
    wire N__51643;
    wire N__51642;
    wire N__51635;
    wire N__51632;
    wire N__51629;
    wire N__51626;
    wire N__51623;
    wire N__51622;
    wire N__51621;
    wire N__51620;
    wire N__51619;
    wire N__51616;
    wire N__51611;
    wire N__51608;
    wire N__51607;
    wire N__51606;
    wire N__51605;
    wire N__51604;
    wire N__51601;
    wire N__51592;
    wire N__51591;
    wire N__51590;
    wire N__51589;
    wire N__51588;
    wire N__51587;
    wire N__51586;
    wire N__51585;
    wire N__51584;
    wire N__51583;
    wire N__51582;
    wire N__51581;
    wire N__51580;
    wire N__51579;
    wire N__51578;
    wire N__51577;
    wire N__51574;
    wire N__51569;
    wire N__51566;
    wire N__51559;
    wire N__51556;
    wire N__51553;
    wire N__51550;
    wire N__51547;
    wire N__51544;
    wire N__51541;
    wire N__51538;
    wire N__51535;
    wire N__51532;
    wire N__51529;
    wire N__51526;
    wire N__51523;
    wire N__51520;
    wire N__51517;
    wire N__51514;
    wire N__51511;
    wire N__51508;
    wire N__51505;
    wire N__51504;
    wire N__51503;
    wire N__51502;
    wire N__51501;
    wire N__51500;
    wire N__51499;
    wire N__51498;
    wire N__51497;
    wire N__51496;
    wire N__51495;
    wire N__51494;
    wire N__51489;
    wire N__51486;
    wire N__51479;
    wire N__51476;
    wire N__51475;
    wire N__51474;
    wire N__51473;
    wire N__51472;
    wire N__51471;
    wire N__51470;
    wire N__51469;
    wire N__51468;
    wire N__51467;
    wire N__51466;
    wire N__51465;
    wire N__51464;
    wire N__51463;
    wire N__51454;
    wire N__51449;
    wire N__51440;
    wire N__51431;
    wire N__51422;
    wire N__51421;
    wire N__51420;
    wire N__51419;
    wire N__51418;
    wire N__51417;
    wire N__51414;
    wire N__51413;
    wire N__51410;
    wire N__51409;
    wire N__51406;
    wire N__51405;
    wire N__51402;
    wire N__51401;
    wire N__51398;
    wire N__51397;
    wire N__51394;
    wire N__51393;
    wire N__51390;
    wire N__51389;
    wire N__51388;
    wire N__51387;
    wire N__51386;
    wire N__51383;
    wire N__51380;
    wire N__51377;
    wire N__51376;
    wire N__51375;
    wire N__51374;
    wire N__51373;
    wire N__51372;
    wire N__51371;
    wire N__51370;
    wire N__51369;
    wire N__51366;
    wire N__51361;
    wire N__51360;
    wire N__51359;
    wire N__51358;
    wire N__51357;
    wire N__51356;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51346;
    wire N__51345;
    wire N__51344;
    wire N__51343;
    wire N__51342;
    wire N__51341;
    wire N__51340;
    wire N__51339;
    wire N__51338;
    wire N__51335;
    wire N__51332;
    wire N__51329;
    wire N__51326;
    wire N__51323;
    wire N__51320;
    wire N__51317;
    wire N__51314;
    wire N__51311;
    wire N__51308;
    wire N__51305;
    wire N__51302;
    wire N__51301;
    wire N__51300;
    wire N__51299;
    wire N__51298;
    wire N__51297;
    wire N__51296;
    wire N__51295;
    wire N__51294;
    wire N__51293;
    wire N__51292;
    wire N__51291;
    wire N__51290;
    wire N__51289;
    wire N__51286;
    wire N__51277;
    wire N__51274;
    wire N__51271;
    wire N__51268;
    wire N__51265;
    wire N__51250;
    wire N__51233;
    wire N__51232;
    wire N__51229;
    wire N__51228;
    wire N__51225;
    wire N__51224;
    wire N__51221;
    wire N__51220;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51204;
    wire N__51201;
    wire N__51192;
    wire N__51189;
    wire N__51186;
    wire N__51183;
    wire N__51172;
    wire N__51171;
    wire N__51170;
    wire N__51169;
    wire N__51168;
    wire N__51161;
    wire N__51152;
    wire N__51143;
    wire N__51142;
    wire N__51133;
    wire N__51124;
    wire N__51115;
    wire N__51112;
    wire N__51109;
    wire N__51106;
    wire N__51103;
    wire N__51100;
    wire N__51097;
    wire N__51094;
    wire N__51091;
    wire N__51090;
    wire N__51087;
    wire N__51086;
    wire N__51085;
    wire N__51084;
    wire N__51081;
    wire N__51080;
    wire N__51079;
    wire N__51078;
    wire N__51077;
    wire N__51076;
    wire N__51075;
    wire N__51074;
    wire N__51071;
    wire N__51070;
    wire N__51067;
    wire N__51066;
    wire N__51063;
    wire N__51062;
    wire N__51061;
    wire N__51060;
    wire N__51055;
    wire N__51050;
    wire N__51045;
    wire N__51040;
    wire N__51025;
    wire N__51022;
    wire N__51013;
    wire N__51010;
    wire N__51001;
    wire N__50998;
    wire N__50993;
    wire N__50990;
    wire N__50989;
    wire N__50982;
    wire N__50979;
    wire N__50976;
    wire N__50971;
    wire N__50962;
    wire N__50957;
    wire N__50952;
    wire N__50949;
    wire N__50946;
    wire N__50939;
    wire N__50936;
    wire N__50927;
    wire N__50922;
    wire N__50907;
    wire N__50904;
    wire N__50901;
    wire N__50900;
    wire N__50893;
    wire N__50888;
    wire N__50885;
    wire N__50882;
    wire N__50871;
    wire N__50868;
    wire N__50863;
    wire N__50852;
    wire N__50849;
    wire N__50844;
    wire N__50837;
    wire N__50834;
    wire N__50827;
    wire N__50824;
    wire N__50821;
    wire N__50818;
    wire N__50815;
    wire N__50810;
    wire N__50805;
    wire N__50800;
    wire N__50797;
    wire N__50794;
    wire N__50791;
    wire N__50786;
    wire N__50783;
    wire N__50778;
    wire N__50771;
    wire N__50766;
    wire N__50755;
    wire N__50754;
    wire N__50751;
    wire N__50750;
    wire N__50749;
    wire N__50748;
    wire N__50745;
    wire N__50744;
    wire N__50741;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50722;
    wire N__50719;
    wire N__50716;
    wire N__50713;
    wire N__50708;
    wire N__50703;
    wire N__50698;
    wire N__50695;
    wire N__50694;
    wire N__50691;
    wire N__50688;
    wire N__50685;
    wire N__50682;
    wire N__50677;
    wire N__50676;
    wire N__50673;
    wire N__50670;
    wire N__50667;
    wire N__50664;
    wire N__50661;
    wire N__50656;
    wire N__50653;
    wire N__50650;
    wire N__50647;
    wire N__50646;
    wire N__50645;
    wire N__50638;
    wire N__50635;
    wire N__50632;
    wire N__50629;
    wire N__50626;
    wire N__50623;
    wire N__50620;
    wire N__50619;
    wire N__50616;
    wire N__50613;
    wire N__50610;
    wire N__50605;
    wire N__50602;
    wire N__50599;
    wire N__50596;
    wire N__50593;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50583;
    wire N__50580;
    wire N__50575;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50563;
    wire N__50560;
    wire N__50559;
    wire N__50556;
    wire N__50553;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50541;
    wire N__50540;
    wire N__50539;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50533;
    wire N__50532;
    wire N__50531;
    wire N__50530;
    wire N__50529;
    wire N__50528;
    wire N__50527;
    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50523;
    wire N__50522;
    wire N__50519;
    wire N__50518;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50510;
    wire N__50505;
    wire N__50502;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50486;
    wire N__50485;
    wire N__50484;
    wire N__50481;
    wire N__50480;
    wire N__50479;
    wire N__50478;
    wire N__50477;
    wire N__50474;
    wire N__50469;
    wire N__50464;
    wire N__50461;
    wire N__50452;
    wire N__50447;
    wire N__50444;
    wire N__50439;
    wire N__50430;
    wire N__50427;
    wire N__50422;
    wire N__50417;
    wire N__50414;
    wire N__50407;
    wire N__50398;
    wire N__50391;
    wire N__50380;
    wire N__50379;
    wire N__50376;
    wire N__50373;
    wire N__50368;
    wire N__50365;
    wire N__50362;
    wire N__50359;
    wire N__50358;
    wire N__50357;
    wire N__50354;
    wire N__50349;
    wire N__50344;
    wire N__50343;
    wire N__50342;
    wire N__50341;
    wire N__50336;
    wire N__50333;
    wire N__50332;
    wire N__50329;
    wire N__50328;
    wire N__50323;
    wire N__50320;
    wire N__50317;
    wire N__50314;
    wire N__50311;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50297;
    wire N__50296;
    wire N__50293;
    wire N__50290;
    wire N__50287;
    wire N__50282;
    wire N__50279;
    wire N__50276;
    wire N__50269;
    wire N__50268;
    wire N__50267;
    wire N__50266;
    wire N__50263;
    wire N__50256;
    wire N__50253;
    wire N__50248;
    wire N__50245;
    wire N__50244;
    wire N__50243;
    wire N__50240;
    wire N__50239;
    wire N__50234;
    wire N__50231;
    wire N__50228;
    wire N__50223;
    wire N__50218;
    wire N__50217;
    wire N__50214;
    wire N__50211;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50179;
    wire N__50176;
    wire N__50173;
    wire N__50170;
    wire N__50167;
    wire N__50164;
    wire N__50161;
    wire N__50158;
    wire N__50155;
    wire N__50152;
    wire N__50149;
    wire N__50146;
    wire N__50143;
    wire N__50140;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50113;
    wire N__50112;
    wire N__50109;
    wire N__50106;
    wire N__50105;
    wire N__50104;
    wire N__50101;
    wire N__50100;
    wire N__50097;
    wire N__50096;
    wire N__50093;
    wire N__50092;
    wire N__50091;
    wire N__50090;
    wire N__50089;
    wire N__50088;
    wire N__50087;
    wire N__50086;
    wire N__50085;
    wire N__50084;
    wire N__50083;
    wire N__50082;
    wire N__50081;
    wire N__50080;
    wire N__50079;
    wire N__50078;
    wire N__50077;
    wire N__50076;
    wire N__50075;
    wire N__50074;
    wire N__50073;
    wire N__50070;
    wire N__50069;
    wire N__50068;
    wire N__50067;
    wire N__50066;
    wire N__50063;
    wire N__50062;
    wire N__50061;
    wire N__50058;
    wire N__50057;
    wire N__50056;
    wire N__50055;
    wire N__50054;
    wire N__50053;
    wire N__50052;
    wire N__50051;
    wire N__50050;
    wire N__50049;
    wire N__50048;
    wire N__50047;
    wire N__50046;
    wire N__50043;
    wire N__50038;
    wire N__50037;
    wire N__50034;
    wire N__50033;
    wire N__50032;
    wire N__50029;
    wire N__50026;
    wire N__50023;
    wire N__50020;
    wire N__50019;
    wire N__50018;
    wire N__50015;
    wire N__50014;
    wire N__50013;
    wire N__50012;
    wire N__50011;
    wire N__50008;
    wire N__50007;
    wire N__50006;
    wire N__50005;
    wire N__50004;
    wire N__50003;
    wire N__50002;
    wire N__50001;
    wire N__50000;
    wire N__49999;
    wire N__49998;
    wire N__49997;
    wire N__49994;
    wire N__49979;
    wire N__49974;
    wire N__49965;
    wire N__49964;
    wire N__49963;
    wire N__49960;
    wire N__49959;
    wire N__49956;
    wire N__49955;
    wire N__49952;
    wire N__49951;
    wire N__49950;
    wire N__49949;
    wire N__49948;
    wire N__49947;
    wire N__49944;
    wire N__49941;
    wire N__49930;
    wire N__49923;
    wire N__49922;
    wire N__49919;
    wire N__49918;
    wire N__49915;
    wire N__49914;
    wire N__49911;
    wire N__49910;
    wire N__49907;
    wire N__49906;
    wire N__49903;
    wire N__49902;
    wire N__49899;
    wire N__49898;
    wire N__49895;
    wire N__49894;
    wire N__49893;
    wire N__49892;
    wire N__49891;
    wire N__49890;
    wire N__49889;
    wire N__49888;
    wire N__49887;
    wire N__49886;
    wire N__49885;
    wire N__49884;
    wire N__49883;
    wire N__49882;
    wire N__49881;
    wire N__49878;
    wire N__49877;
    wire N__49874;
    wire N__49861;
    wire N__49850;
    wire N__49833;
    wire N__49830;
    wire N__49829;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49821;
    wire N__49818;
    wire N__49817;
    wire N__49814;
    wire N__49805;
    wire N__49800;
    wire N__49797;
    wire N__49780;
    wire N__49779;
    wire N__49776;
    wire N__49775;
    wire N__49772;
    wire N__49771;
    wire N__49768;
    wire N__49767;
    wire N__49764;
    wire N__49761;
    wire N__49754;
    wire N__49739;
    wire N__49722;
    wire N__49719;
    wire N__49718;
    wire N__49715;
    wire N__49714;
    wire N__49711;
    wire N__49710;
    wire N__49707;
    wire N__49706;
    wire N__49703;
    wire N__49702;
    wire N__49699;
    wire N__49698;
    wire N__49695;
    wire N__49694;
    wire N__49691;
    wire N__49690;
    wire N__49689;
    wire N__49688;
    wire N__49685;
    wire N__49684;
    wire N__49681;
    wire N__49680;
    wire N__49679;
    wire N__49676;
    wire N__49675;
    wire N__49672;
    wire N__49671;
    wire N__49668;
    wire N__49665;
    wire N__49662;
    wire N__49653;
    wire N__49650;
    wire N__49633;
    wire N__49628;
    wire N__49623;
    wire N__49606;
    wire N__49597;
    wire N__49580;
    wire N__49563;
    wire N__49560;
    wire N__49549;
    wire N__49536;
    wire N__49507;
    wire N__49506;
    wire N__49505;
    wire N__49504;
    wire N__49503;
    wire N__49502;
    wire N__49501;
    wire N__49500;
    wire N__49499;
    wire N__49498;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49483;
    wire N__49480;
    wire N__49473;
    wire N__49472;
    wire N__49471;
    wire N__49470;
    wire N__49469;
    wire N__49468;
    wire N__49467;
    wire N__49466;
    wire N__49465;
    wire N__49460;
    wire N__49457;
    wire N__49454;
    wire N__49453;
    wire N__49452;
    wire N__49449;
    wire N__49448;
    wire N__49447;
    wire N__49446;
    wire N__49439;
    wire N__49422;
    wire N__49419;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49413;
    wire N__49412;
    wire N__49411;
    wire N__49410;
    wire N__49409;
    wire N__49408;
    wire N__49405;
    wire N__49400;
    wire N__49397;
    wire N__49390;
    wire N__49381;
    wire N__49380;
    wire N__49379;
    wire N__49378;
    wire N__49377;
    wire N__49376;
    wire N__49375;
    wire N__49374;
    wire N__49373;
    wire N__49372;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49368;
    wire N__49367;
    wire N__49366;
    wire N__49365;
    wire N__49364;
    wire N__49363;
    wire N__49362;
    wire N__49361;
    wire N__49360;
    wire N__49355;
    wire N__49354;
    wire N__49353;
    wire N__49352;
    wire N__49351;
    wire N__49350;
    wire N__49349;
    wire N__49348;
    wire N__49347;
    wire N__49346;
    wire N__49345;
    wire N__49334;
    wire N__49333;
    wire N__49332;
    wire N__49331;
    wire N__49328;
    wire N__49327;
    wire N__49326;
    wire N__49321;
    wire N__49316;
    wire N__49313;
    wire N__49304;
    wire N__49291;
    wire N__49274;
    wire N__49267;
    wire N__49264;
    wire N__49249;
    wire N__49242;
    wire N__49239;
    wire N__49226;
    wire N__49221;
    wire N__49198;
    wire N__49195;
    wire N__49192;
    wire N__49189;
    wire N__49186;
    wire N__49183;
    wire N__49180;
    wire N__49177;
    wire N__49174;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49166;
    wire N__49165;
    wire N__49164;
    wire N__49163;
    wire N__49162;
    wire N__49161;
    wire N__49160;
    wire N__49159;
    wire N__49158;
    wire N__49157;
    wire N__49156;
    wire N__49155;
    wire N__49150;
    wire N__49145;
    wire N__49142;
    wire N__49137;
    wire N__49122;
    wire N__49121;
    wire N__49120;
    wire N__49119;
    wire N__49118;
    wire N__49117;
    wire N__49116;
    wire N__49115;
    wire N__49114;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49108;
    wire N__49107;
    wire N__49106;
    wire N__49105;
    wire N__49104;
    wire N__49101;
    wire N__49098;
    wire N__49091;
    wire N__49080;
    wire N__49063;
    wire N__49052;
    wire N__49039;
    wire N__49036;
    wire N__49033;
    wire N__49030;
    wire N__49027;
    wire N__49024;
    wire N__49023;
    wire N__49020;
    wire N__49017;
    wire N__49012;
    wire N__49009;
    wire N__49006;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48979;
    wire N__48976;
    wire N__48973;
    wire N__48970;
    wire N__48967;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48952;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48940;
    wire N__48937;
    wire N__48934;
    wire N__48931;
    wire N__48928;
    wire N__48925;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48895;
    wire N__48892;
    wire N__48889;
    wire N__48886;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48868;
    wire N__48865;
    wire N__48862;
    wire N__48859;
    wire N__48856;
    wire N__48853;
    wire N__48850;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48838;
    wire N__48835;
    wire N__48832;
    wire N__48829;
    wire N__48826;
    wire N__48823;
    wire N__48820;
    wire N__48817;
    wire N__48814;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48802;
    wire N__48799;
    wire N__48796;
    wire N__48793;
    wire N__48790;
    wire N__48787;
    wire N__48784;
    wire N__48781;
    wire N__48778;
    wire N__48775;
    wire N__48772;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48727;
    wire N__48724;
    wire N__48721;
    wire N__48718;
    wire N__48715;
    wire N__48712;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48697;
    wire N__48694;
    wire N__48691;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48673;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48658;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48637;
    wire N__48634;
    wire N__48631;
    wire N__48628;
    wire N__48625;
    wire N__48622;
    wire N__48619;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48598;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48568;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48544;
    wire N__48541;
    wire N__48538;
    wire N__48535;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48523;
    wire N__48520;
    wire N__48517;
    wire N__48514;
    wire N__48511;
    wire N__48508;
    wire N__48505;
    wire N__48502;
    wire N__48499;
    wire N__48496;
    wire N__48493;
    wire N__48490;
    wire N__48487;
    wire N__48484;
    wire N__48481;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48463;
    wire N__48460;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48442;
    wire N__48439;
    wire N__48436;
    wire N__48433;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48418;
    wire N__48415;
    wire N__48412;
    wire N__48409;
    wire N__48406;
    wire N__48403;
    wire N__48400;
    wire N__48397;
    wire N__48394;
    wire N__48393;
    wire N__48390;
    wire N__48387;
    wire N__48386;
    wire N__48381;
    wire N__48378;
    wire N__48373;
    wire N__48372;
    wire N__48369;
    wire N__48366;
    wire N__48361;
    wire N__48360;
    wire N__48357;
    wire N__48354;
    wire N__48351;
    wire N__48350;
    wire N__48347;
    wire N__48344;
    wire N__48341;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48327;
    wire N__48326;
    wire N__48323;
    wire N__48318;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48303;
    wire N__48302;
    wire N__48301;
    wire N__48298;
    wire N__48291;
    wire N__48286;
    wire N__48283;
    wire N__48280;
    wire N__48277;
    wire N__48274;
    wire N__48273;
    wire N__48268;
    wire N__48265;
    wire N__48264;
    wire N__48261;
    wire N__48258;
    wire N__48253;
    wire N__48250;
    wire N__48249;
    wire N__48244;
    wire N__48243;
    wire N__48242;
    wire N__48239;
    wire N__48234;
    wire N__48231;
    wire N__48228;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48214;
    wire N__48213;
    wire N__48210;
    wire N__48207;
    wire N__48206;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48196;
    wire N__48193;
    wire N__48184;
    wire N__48181;
    wire N__48178;
    wire N__48175;
    wire N__48172;
    wire N__48169;
    wire N__48166;
    wire N__48163;
    wire N__48160;
    wire N__48157;
    wire N__48154;
    wire N__48151;
    wire N__48148;
    wire N__48145;
    wire N__48142;
    wire N__48139;
    wire N__48136;
    wire N__48133;
    wire N__48130;
    wire N__48127;
    wire N__48124;
    wire N__48121;
    wire N__48118;
    wire N__48117;
    wire N__48116;
    wire N__48115;
    wire N__48112;
    wire N__48109;
    wire N__48104;
    wire N__48097;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48083;
    wire N__48078;
    wire N__48075;
    wire N__48070;
    wire N__48067;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48059;
    wire N__48054;
    wire N__48051;
    wire N__48050;
    wire N__48045;
    wire N__48042;
    wire N__48037;
    wire N__48034;
    wire N__48033;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48020;
    wire N__48017;
    wire N__48010;
    wire N__48007;
    wire N__48006;
    wire N__48005;
    wire N__48002;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47986;
    wire N__47983;
    wire N__47980;
    wire N__47977;
    wire N__47974;
    wire N__47965;
    wire N__47964;
    wire N__47961;
    wire N__47960;
    wire N__47957;
    wire N__47954;
    wire N__47951;
    wire N__47948;
    wire N__47945;
    wire N__47938;
    wire N__47935;
    wire N__47934;
    wire N__47931;
    wire N__47930;
    wire N__47927;
    wire N__47924;
    wire N__47921;
    wire N__47914;
    wire N__47911;
    wire N__47910;
    wire N__47907;
    wire N__47904;
    wire N__47901;
    wire N__47898;
    wire N__47897;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47887;
    wire N__47884;
    wire N__47879;
    wire N__47876;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47862;
    wire N__47859;
    wire N__47858;
    wire N__47855;
    wire N__47852;
    wire N__47849;
    wire N__47846;
    wire N__47841;
    wire N__47838;
    wire N__47835;
    wire N__47830;
    wire N__47829;
    wire N__47826;
    wire N__47825;
    wire N__47822;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47806;
    wire N__47803;
    wire N__47802;
    wire N__47801;
    wire N__47798;
    wire N__47795;
    wire N__47792;
    wire N__47789;
    wire N__47786;
    wire N__47783;
    wire N__47776;
    wire N__47775;
    wire N__47772;
    wire N__47769;
    wire N__47768;
    wire N__47765;
    wire N__47762;
    wire N__47759;
    wire N__47758;
    wire N__47755;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47738;
    wire N__47731;
    wire N__47728;
    wire N__47727;
    wire N__47724;
    wire N__47721;
    wire N__47720;
    wire N__47719;
    wire N__47716;
    wire N__47713;
    wire N__47710;
    wire N__47707;
    wire N__47698;
    wire N__47695;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47678;
    wire N__47671;
    wire N__47668;
    wire N__47665;
    wire N__47664;
    wire N__47661;
    wire N__47660;
    wire N__47657;
    wire N__47654;
    wire N__47651;
    wire N__47644;
    wire N__47641;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47633;
    wire N__47630;
    wire N__47627;
    wire N__47624;
    wire N__47623;
    wire N__47620;
    wire N__47615;
    wire N__47612;
    wire N__47605;
    wire N__47604;
    wire N__47601;
    wire N__47598;
    wire N__47593;
    wire N__47590;
    wire N__47587;
    wire N__47584;
    wire N__47581;
    wire N__47580;
    wire N__47577;
    wire N__47574;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47564;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47552;
    wire N__47549;
    wire N__47546;
    wire N__47539;
    wire N__47536;
    wire N__47535;
    wire N__47534;
    wire N__47531;
    wire N__47528;
    wire N__47525;
    wire N__47524;
    wire N__47519;
    wire N__47514;
    wire N__47511;
    wire N__47506;
    wire N__47503;
    wire N__47502;
    wire N__47501;
    wire N__47498;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47470;
    wire N__47469;
    wire N__47468;
    wire N__47467;
    wire N__47464;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47452;
    wire N__47447;
    wire N__47444;
    wire N__47437;
    wire N__47434;
    wire N__47433;
    wire N__47430;
    wire N__47427;
    wire N__47426;
    wire N__47421;
    wire N__47418;
    wire N__47413;
    wire N__47412;
    wire N__47409;
    wire N__47406;
    wire N__47401;
    wire N__47400;
    wire N__47397;
    wire N__47394;
    wire N__47393;
    wire N__47390;
    wire N__47387;
    wire N__47384;
    wire N__47379;
    wire N__47376;
    wire N__47371;
    wire N__47368;
    wire N__47367;
    wire N__47364;
    wire N__47361;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47353;
    wire N__47350;
    wire N__47345;
    wire N__47342;
    wire N__47339;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47320;
    wire N__47319;
    wire N__47316;
    wire N__47315;
    wire N__47312;
    wire N__47309;
    wire N__47306;
    wire N__47299;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47285;
    wire N__47282;
    wire N__47279;
    wire N__47276;
    wire N__47275;
    wire N__47270;
    wire N__47267;
    wire N__47264;
    wire N__47257;
    wire N__47256;
    wire N__47255;
    wire N__47254;
    wire N__47253;
    wire N__47252;
    wire N__47251;
    wire N__47250;
    wire N__47249;
    wire N__47248;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47243;
    wire N__47242;
    wire N__47241;
    wire N__47240;
    wire N__47239;
    wire N__47238;
    wire N__47237;
    wire N__47236;
    wire N__47235;
    wire N__47234;
    wire N__47233;
    wire N__47232;
    wire N__47231;
    wire N__47230;
    wire N__47229;
    wire N__47228;
    wire N__47219;
    wire N__47210;
    wire N__47201;
    wire N__47192;
    wire N__47183;
    wire N__47174;
    wire N__47169;
    wire N__47160;
    wire N__47157;
    wire N__47146;
    wire N__47137;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47127;
    wire N__47124;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47114;
    wire N__47107;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47094;
    wire N__47089;
    wire N__47088;
    wire N__47087;
    wire N__47084;
    wire N__47079;
    wire N__47074;
    wire N__47071;
    wire N__47070;
    wire N__47067;
    wire N__47064;
    wire N__47063;
    wire N__47058;
    wire N__47055;
    wire N__47054;
    wire N__47051;
    wire N__47048;
    wire N__47045;
    wire N__47038;
    wire N__47037;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47027;
    wire N__47022;
    wire N__47017;
    wire N__47014;
    wire N__47011;
    wire N__47008;
    wire N__47005;
    wire N__47002;
    wire N__46999;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46989;
    wire N__46986;
    wire N__46983;
    wire N__46978;
    wire N__46975;
    wire N__46972;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46960;
    wire N__46957;
    wire N__46954;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46942;
    wire N__46939;
    wire N__46938;
    wire N__46935;
    wire N__46932;
    wire N__46927;
    wire N__46924;
    wire N__46921;
    wire N__46920;
    wire N__46917;
    wire N__46914;
    wire N__46909;
    wire N__46908;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46894;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46882;
    wire N__46879;
    wire N__46876;
    wire N__46873;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46863;
    wire N__46862;
    wire N__46861;
    wire N__46858;
    wire N__46855;
    wire N__46852;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46832;
    wire N__46829;
    wire N__46826;
    wire N__46821;
    wire N__46816;
    wire N__46813;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46803;
    wire N__46800;
    wire N__46795;
    wire N__46794;
    wire N__46791;
    wire N__46788;
    wire N__46787;
    wire N__46784;
    wire N__46781;
    wire N__46778;
    wire N__46771;
    wire N__46770;
    wire N__46765;
    wire N__46764;
    wire N__46761;
    wire N__46758;
    wire N__46753;
    wire N__46750;
    wire N__46747;
    wire N__46744;
    wire N__46741;
    wire N__46738;
    wire N__46737;
    wire N__46734;
    wire N__46731;
    wire N__46726;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46708;
    wire N__46705;
    wire N__46702;
    wire N__46699;
    wire N__46698;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46681;
    wire N__46678;
    wire N__46675;
    wire N__46672;
    wire N__46669;
    wire N__46666;
    wire N__46663;
    wire N__46660;
    wire N__46659;
    wire N__46656;
    wire N__46653;
    wire N__46648;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46632;
    wire N__46627;
    wire N__46624;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46612;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46600;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46590;
    wire N__46587;
    wire N__46584;
    wire N__46581;
    wire N__46576;
    wire N__46573;
    wire N__46570;
    wire N__46569;
    wire N__46566;
    wire N__46563;
    wire N__46558;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46522;
    wire N__46521;
    wire N__46520;
    wire N__46519;
    wire N__46518;
    wire N__46509;
    wire N__46508;
    wire N__46507;
    wire N__46506;
    wire N__46505;
    wire N__46504;
    wire N__46503;
    wire N__46502;
    wire N__46501;
    wire N__46500;
    wire N__46499;
    wire N__46490;
    wire N__46487;
    wire N__46478;
    wire N__46469;
    wire N__46468;
    wire N__46467;
    wire N__46466;
    wire N__46465;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46461;
    wire N__46460;
    wire N__46459;
    wire N__46458;
    wire N__46457;
    wire N__46452;
    wire N__46443;
    wire N__46434;
    wire N__46425;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46403;
    wire N__46396;
    wire N__46393;
    wire N__46392;
    wire N__46389;
    wire N__46386;
    wire N__46385;
    wire N__46380;
    wire N__46377;
    wire N__46374;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46362;
    wire N__46359;
    wire N__46356;
    wire N__46355;
    wire N__46350;
    wire N__46347;
    wire N__46344;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46318;
    wire N__46315;
    wire N__46312;
    wire N__46311;
    wire N__46308;
    wire N__46305;
    wire N__46302;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46290;
    wire N__46287;
    wire N__46284;
    wire N__46279;
    wire N__46276;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46264;
    wire N__46263;
    wire N__46260;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46231;
    wire N__46228;
    wire N__46225;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46213;
    wire N__46210;
    wire N__46209;
    wire N__46206;
    wire N__46203;
    wire N__46198;
    wire N__46197;
    wire N__46194;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46180;
    wire N__46177;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46165;
    wire N__46164;
    wire N__46159;
    wire N__46158;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46144;
    wire N__46141;
    wire N__46140;
    wire N__46139;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46123;
    wire N__46120;
    wire N__46119;
    wire N__46116;
    wire N__46113;
    wire N__46112;
    wire N__46107;
    wire N__46104;
    wire N__46101;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46089;
    wire N__46086;
    wire N__46085;
    wire N__46082;
    wire N__46079;
    wire N__46076;
    wire N__46071;
    wire N__46066;
    wire N__46063;
    wire N__46062;
    wire N__46061;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46045;
    wire N__46042;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46034;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46011;
    wire N__46010;
    wire N__46007;
    wire N__46004;
    wire N__46001;
    wire N__45998;
    wire N__45995;
    wire N__45990;
    wire N__45987;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45972;
    wire N__45971;
    wire N__45968;
    wire N__45965;
    wire N__45962;
    wire N__45959;
    wire N__45956;
    wire N__45949;
    wire N__45946;
    wire N__45943;
    wire N__45942;
    wire N__45941;
    wire N__45938;
    wire N__45935;
    wire N__45932;
    wire N__45929;
    wire N__45926;
    wire N__45921;
    wire N__45918;
    wire N__45913;
    wire N__45910;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45902;
    wire N__45897;
    wire N__45894;
    wire N__45891;
    wire N__45886;
    wire N__45883;
    wire N__45882;
    wire N__45877;
    wire N__45876;
    wire N__45873;
    wire N__45870;
    wire N__45867;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45848;
    wire N__45843;
    wire N__45840;
    wire N__45837;
    wire N__45832;
    wire N__45829;
    wire N__45826;
    wire N__45825;
    wire N__45822;
    wire N__45821;
    wire N__45818;
    wire N__45815;
    wire N__45812;
    wire N__45807;
    wire N__45802;
    wire N__45799;
    wire N__45798;
    wire N__45797;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45781;
    wire N__45778;
    wire N__45777;
    wire N__45774;
    wire N__45771;
    wire N__45770;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45754;
    wire N__45751;
    wire N__45748;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45731;
    wire N__45726;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45711;
    wire N__45710;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45698;
    wire N__45695;
    wire N__45688;
    wire N__45685;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45663;
    wire N__45658;
    wire N__45655;
    wire N__45652;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45644;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45628;
    wire N__45625;
    wire N__45624;
    wire N__45623;
    wire N__45618;
    wire N__45615;
    wire N__45612;
    wire N__45607;
    wire N__45604;
    wire N__45603;
    wire N__45600;
    wire N__45597;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45587;
    wire N__45582;
    wire N__45577;
    wire N__45574;
    wire N__45573;
    wire N__45570;
    wire N__45567;
    wire N__45562;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45552;
    wire N__45547;
    wire N__45544;
    wire N__45543;
    wire N__45542;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45512;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45496;
    wire N__45493;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45471;
    wire N__45466;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45430;
    wire N__45427;
    wire N__45424;
    wire N__45421;
    wire N__45418;
    wire N__45415;
    wire N__45412;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45379;
    wire N__45376;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45358;
    wire N__45355;
    wire N__45352;
    wire N__45349;
    wire N__45346;
    wire N__45343;
    wire N__45340;
    wire N__45337;
    wire N__45334;
    wire N__45331;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45319;
    wire N__45316;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45304;
    wire N__45303;
    wire N__45300;
    wire N__45297;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45280;
    wire N__45277;
    wire N__45274;
    wire N__45271;
    wire N__45268;
    wire N__45265;
    wire N__45262;
    wire N__45259;
    wire N__45256;
    wire N__45253;
    wire N__45250;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45232;
    wire N__45229;
    wire N__45226;
    wire N__45223;
    wire N__45220;
    wire N__45217;
    wire N__45214;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45199;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45187;
    wire N__45184;
    wire N__45181;
    wire N__45178;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45157;
    wire N__45154;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45142;
    wire N__45139;
    wire N__45136;
    wire N__45133;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45118;
    wire N__45115;
    wire N__45112;
    wire N__45109;
    wire N__45106;
    wire N__45103;
    wire N__45100;
    wire N__45097;
    wire N__45094;
    wire N__45091;
    wire N__45088;
    wire N__45085;
    wire N__45082;
    wire N__45079;
    wire N__45076;
    wire N__45073;
    wire N__45070;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45046;
    wire N__45043;
    wire N__45040;
    wire N__45037;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44980;
    wire N__44977;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44962;
    wire N__44959;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44947;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44935;
    wire N__44932;
    wire N__44929;
    wire N__44926;
    wire N__44923;
    wire N__44920;
    wire N__44917;
    wire N__44914;
    wire N__44911;
    wire N__44908;
    wire N__44905;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44875;
    wire N__44872;
    wire N__44869;
    wire N__44866;
    wire N__44863;
    wire N__44860;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44848;
    wire N__44845;
    wire N__44842;
    wire N__44839;
    wire N__44836;
    wire N__44833;
    wire N__44830;
    wire N__44827;
    wire N__44824;
    wire N__44821;
    wire N__44818;
    wire N__44815;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44803;
    wire N__44800;
    wire N__44797;
    wire N__44794;
    wire N__44791;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44773;
    wire N__44770;
    wire N__44767;
    wire N__44766;
    wire N__44765;
    wire N__44762;
    wire N__44761;
    wire N__44756;
    wire N__44753;
    wire N__44750;
    wire N__44747;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44731;
    wire N__44730;
    wire N__44727;
    wire N__44724;
    wire N__44723;
    wire N__44720;
    wire N__44717;
    wire N__44714;
    wire N__44707;
    wire N__44706;
    wire N__44705;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44683;
    wire N__44682;
    wire N__44677;
    wire N__44676;
    wire N__44673;
    wire N__44670;
    wire N__44669;
    wire N__44664;
    wire N__44661;
    wire N__44656;
    wire N__44655;
    wire N__44654;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44640;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44614;
    wire N__44611;
    wire N__44608;
    wire N__44605;
    wire N__44602;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44581;
    wire N__44578;
    wire N__44575;
    wire N__44574;
    wire N__44569;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44561;
    wire N__44556;
    wire N__44553;
    wire N__44548;
    wire N__44547;
    wire N__44544;
    wire N__44543;
    wire N__44540;
    wire N__44535;
    wire N__44532;
    wire N__44527;
    wire N__44526;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44513;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44503;
    wire N__44498;
    wire N__44495;
    wire N__44492;
    wire N__44485;
    wire N__44484;
    wire N__44481;
    wire N__44478;
    wire N__44477;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44461;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44443;
    wire N__44440;
    wire N__44435;
    wire N__44432;
    wire N__44425;
    wire N__44422;
    wire N__44421;
    wire N__44418;
    wire N__44415;
    wire N__44414;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44398;
    wire N__44395;
    wire N__44392;
    wire N__44391;
    wire N__44390;
    wire N__44387;
    wire N__44384;
    wire N__44381;
    wire N__44378;
    wire N__44375;
    wire N__44372;
    wire N__44371;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44353;
    wire N__44350;
    wire N__44349;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44334;
    wire N__44329;
    wire N__44328;
    wire N__44325;
    wire N__44324;
    wire N__44321;
    wire N__44320;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44299;
    wire N__44296;
    wire N__44293;
    wire N__44292;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44277;
    wire N__44272;
    wire N__44271;
    wire N__44266;
    wire N__44265;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44248;
    wire N__44247;
    wire N__44244;
    wire N__44243;
    wire N__44238;
    wire N__44235;
    wire N__44230;
    wire N__44227;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44197;
    wire N__44196;
    wire N__44195;
    wire N__44194;
    wire N__44193;
    wire N__44192;
    wire N__44191;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44166;
    wire N__44161;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44149;
    wire N__44148;
    wire N__44147;
    wire N__44144;
    wire N__44139;
    wire N__44136;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44126;
    wire N__44119;
    wire N__44118;
    wire N__44115;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44078;
    wire N__44077;
    wire N__44072;
    wire N__44067;
    wire N__44062;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44045;
    wire N__44044;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44026;
    wire N__44023;
    wire N__44022;
    wire N__44021;
    wire N__44018;
    wire N__44015;
    wire N__44012;
    wire N__44005;
    wire N__44002;
    wire N__43999;
    wire N__43996;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43978;
    wire N__43975;
    wire N__43972;
    wire N__43971;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43963;
    wire N__43960;
    wire N__43959;
    wire N__43956;
    wire N__43953;
    wire N__43950;
    wire N__43947;
    wire N__43944;
    wire N__43941;
    wire N__43938;
    wire N__43935;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43921;
    wire N__43918;
    wire N__43909;
    wire N__43906;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43878;
    wire N__43875;
    wire N__43872;
    wire N__43867;
    wire N__43864;
    wire N__43863;
    wire N__43860;
    wire N__43857;
    wire N__43852;
    wire N__43849;
    wire N__43848;
    wire N__43845;
    wire N__43842;
    wire N__43839;
    wire N__43836;
    wire N__43833;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43821;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43801;
    wire N__43798;
    wire N__43795;
    wire N__43792;
    wire N__43789;
    wire N__43786;
    wire N__43783;
    wire N__43780;
    wire N__43777;
    wire N__43774;
    wire N__43771;
    wire N__43768;
    wire N__43765;
    wire N__43762;
    wire N__43759;
    wire N__43756;
    wire N__43753;
    wire N__43752;
    wire N__43747;
    wire N__43744;
    wire N__43741;
    wire N__43738;
    wire N__43737;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43725;
    wire N__43722;
    wire N__43719;
    wire N__43714;
    wire N__43711;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43660;
    wire N__43657;
    wire N__43656;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43630;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43620;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43610;
    wire N__43605;
    wire N__43602;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43567;
    wire N__43564;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43522;
    wire N__43519;
    wire N__43516;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43501;
    wire N__43500;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43490;
    wire N__43489;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43471;
    wire N__43468;
    wire N__43467;
    wire N__43464;
    wire N__43461;
    wire N__43460;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43448;
    wire N__43443;
    wire N__43438;
    wire N__43435;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43420;
    wire N__43419;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43396;
    wire N__43389;
    wire N__43386;
    wire N__43381;
    wire N__43380;
    wire N__43379;
    wire N__43376;
    wire N__43373;
    wire N__43370;
    wire N__43365;
    wire N__43362;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43303;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43282;
    wire N__43279;
    wire N__43276;
    wire N__43273;
    wire N__43270;
    wire N__43267;
    wire N__43264;
    wire N__43261;
    wire N__43258;
    wire N__43255;
    wire N__43252;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43240;
    wire N__43237;
    wire N__43236;
    wire N__43235;
    wire N__43234;
    wire N__43233;
    wire N__43232;
    wire N__43231;
    wire N__43230;
    wire N__43229;
    wire N__43224;
    wire N__43223;
    wire N__43222;
    wire N__43221;
    wire N__43220;
    wire N__43219;
    wire N__43218;
    wire N__43207;
    wire N__43202;
    wire N__43199;
    wire N__43192;
    wire N__43185;
    wire N__43184;
    wire N__43183;
    wire N__43182;
    wire N__43181;
    wire N__43180;
    wire N__43179;
    wire N__43178;
    wire N__43177;
    wire N__43176;
    wire N__43175;
    wire N__43170;
    wire N__43163;
    wire N__43154;
    wire N__43147;
    wire N__43144;
    wire N__43139;
    wire N__43126;
    wire N__43123;
    wire N__43120;
    wire N__43117;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43102;
    wire N__43099;
    wire N__43096;
    wire N__43093;
    wire N__43090;
    wire N__43089;
    wire N__43086;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43071;
    wire N__43066;
    wire N__43063;
    wire N__43060;
    wire N__43057;
    wire N__43054;
    wire N__43051;
    wire N__43048;
    wire N__43045;
    wire N__43042;
    wire N__43039;
    wire N__43036;
    wire N__43033;
    wire N__43030;
    wire N__43027;
    wire N__43024;
    wire N__43021;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42949;
    wire N__42946;
    wire N__42943;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42922;
    wire N__42919;
    wire N__42916;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42883;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42850;
    wire N__42847;
    wire N__42844;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42817;
    wire N__42814;
    wire N__42811;
    wire N__42808;
    wire N__42805;
    wire N__42802;
    wire N__42799;
    wire N__42796;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42766;
    wire N__42763;
    wire N__42760;
    wire N__42757;
    wire N__42754;
    wire N__42751;
    wire N__42748;
    wire N__42745;
    wire N__42742;
    wire N__42739;
    wire N__42736;
    wire N__42733;
    wire N__42730;
    wire N__42727;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42712;
    wire N__42709;
    wire N__42706;
    wire N__42703;
    wire N__42700;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42688;
    wire N__42685;
    wire N__42682;
    wire N__42679;
    wire N__42676;
    wire N__42673;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42652;
    wire N__42649;
    wire N__42646;
    wire N__42643;
    wire N__42640;
    wire N__42639;
    wire N__42636;
    wire N__42635;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42597;
    wire N__42594;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42580;
    wire N__42577;
    wire N__42574;
    wire N__42571;
    wire N__42568;
    wire N__42565;
    wire N__42562;
    wire N__42559;
    wire N__42556;
    wire N__42555;
    wire N__42552;
    wire N__42549;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42525;
    wire N__42522;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42502;
    wire N__42499;
    wire N__42498;
    wire N__42495;
    wire N__42492;
    wire N__42487;
    wire N__42484;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42472;
    wire N__42469;
    wire N__42466;
    wire N__42463;
    wire N__42460;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42442;
    wire N__42439;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42420;
    wire N__42417;
    wire N__42414;
    wire N__42409;
    wire N__42406;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42382;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42370;
    wire N__42367;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42355;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42343;
    wire N__42340;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42328;
    wire N__42325;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42313;
    wire N__42310;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42298;
    wire N__42295;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42277;
    wire N__42274;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42244;
    wire N__42241;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42220;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42193;
    wire N__42190;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42178;
    wire N__42175;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42163;
    wire N__42160;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42148;
    wire N__42145;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42133;
    wire N__42130;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42112;
    wire N__42109;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42097;
    wire N__42094;
    wire N__42091;
    wire N__42088;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42076;
    wire N__42073;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42061;
    wire N__42058;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42046;
    wire N__42043;
    wire N__42040;
    wire N__42039;
    wire N__42038;
    wire N__42037;
    wire N__42034;
    wire N__42033;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42022;
    wire N__42019;
    wire N__42016;
    wire N__42013;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41996;
    wire N__41993;
    wire N__41990;
    wire N__41983;
    wire N__41978;
    wire N__41973;
    wire N__41968;
    wire N__41965;
    wire N__41962;
    wire N__41959;
    wire N__41956;
    wire N__41953;
    wire N__41952;
    wire N__41949;
    wire N__41948;
    wire N__41947;
    wire N__41944;
    wire N__41941;
    wire N__41938;
    wire N__41935;
    wire N__41934;
    wire N__41933;
    wire N__41932;
    wire N__41929;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41915;
    wire N__41912;
    wire N__41905;
    wire N__41902;
    wire N__41899;
    wire N__41896;
    wire N__41893;
    wire N__41890;
    wire N__41887;
    wire N__41884;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41848;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41832;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41809;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41796;
    wire N__41793;
    wire N__41790;
    wire N__41785;
    wire N__41782;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41770;
    wire N__41767;
    wire N__41764;
    wire N__41761;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41740;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41719;
    wire N__41716;
    wire N__41715;
    wire N__41710;
    wire N__41707;
    wire N__41704;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41692;
    wire N__41689;
    wire N__41688;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41674;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41661;
    wire N__41658;
    wire N__41655;
    wire N__41650;
    wire N__41647;
    wire N__41646;
    wire N__41643;
    wire N__41640;
    wire N__41635;
    wire N__41632;
    wire N__41629;
    wire N__41626;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41607;
    wire N__41604;
    wire N__41601;
    wire N__41598;
    wire N__41595;
    wire N__41590;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41572;
    wire N__41569;
    wire N__41566;
    wire N__41563;
    wire N__41560;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41550;
    wire N__41547;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41533;
    wire N__41530;
    wire N__41527;
    wire N__41524;
    wire N__41521;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41479;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41434;
    wire N__41431;
    wire N__41428;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41398;
    wire N__41395;
    wire N__41392;
    wire N__41389;
    wire N__41386;
    wire N__41383;
    wire N__41380;
    wire N__41377;
    wire N__41374;
    wire N__41371;
    wire N__41368;
    wire N__41365;
    wire N__41362;
    wire N__41359;
    wire N__41356;
    wire N__41353;
    wire N__41350;
    wire N__41347;
    wire N__41344;
    wire N__41341;
    wire N__41338;
    wire N__41335;
    wire N__41332;
    wire N__41329;
    wire N__41326;
    wire N__41323;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41308;
    wire N__41305;
    wire N__41302;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41290;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41269;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41257;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41245;
    wire N__41244;
    wire N__41243;
    wire N__41240;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41217;
    wire N__41214;
    wire N__41211;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41175;
    wire N__41172;
    wire N__41169;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41146;
    wire N__41143;
    wire N__41140;
    wire N__41137;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41100;
    wire N__41097;
    wire N__41094;
    wire N__41089;
    wire N__41086;
    wire N__41083;
    wire N__41080;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41038;
    wire N__41035;
    wire N__41032;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41008;
    wire N__41005;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40992;
    wire N__40989;
    wire N__40986;
    wire N__40981;
    wire N__40978;
    wire N__40977;
    wire N__40974;
    wire N__40971;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40957;
    wire N__40956;
    wire N__40953;
    wire N__40950;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40933;
    wire N__40930;
    wire N__40927;
    wire N__40924;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40912;
    wire N__40909;
    wire N__40906;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40864;
    wire N__40861;
    wire N__40858;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40840;
    wire N__40837;
    wire N__40834;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40816;
    wire N__40813;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40803;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40771;
    wire N__40768;
    wire N__40765;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40636;
    wire N__40633;
    wire N__40630;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40549;
    wire N__40546;
    wire N__40543;
    wire N__40540;
    wire N__40537;
    wire N__40534;
    wire N__40531;
    wire N__40528;
    wire N__40525;
    wire N__40522;
    wire N__40519;
    wire N__40516;
    wire N__40513;
    wire N__40510;
    wire N__40507;
    wire N__40504;
    wire N__40503;
    wire N__40500;
    wire N__40497;
    wire N__40494;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40468;
    wire N__40467;
    wire N__40464;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40450;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40426;
    wire N__40423;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40411;
    wire N__40408;
    wire N__40407;
    wire N__40402;
    wire N__40399;
    wire N__40396;
    wire N__40393;
    wire N__40392;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40377;
    wire N__40372;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40360;
    wire N__40357;
    wire N__40354;
    wire N__40351;
    wire N__40348;
    wire N__40345;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40327;
    wire N__40324;
    wire N__40321;
    wire N__40318;
    wire N__40315;
    wire N__40312;
    wire N__40309;
    wire N__40306;
    wire N__40303;
    wire N__40300;
    wire N__40297;
    wire N__40294;
    wire N__40291;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40273;
    wire N__40270;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40252;
    wire N__40249;
    wire N__40246;
    wire N__40243;
    wire N__40240;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40228;
    wire N__40225;
    wire N__40222;
    wire N__40219;
    wire N__40216;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40204;
    wire N__40201;
    wire N__40198;
    wire N__40195;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40183;
    wire N__40180;
    wire N__40177;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40123;
    wire N__40120;
    wire N__40117;
    wire N__40114;
    wire N__40111;
    wire N__40108;
    wire N__40105;
    wire N__40102;
    wire N__40099;
    wire N__40096;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40084;
    wire N__40081;
    wire N__40078;
    wire N__40075;
    wire N__40072;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40006;
    wire N__40003;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39973;
    wire N__39970;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39950;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39934;
    wire N__39931;
    wire N__39930;
    wire N__39925;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39910;
    wire N__39907;
    wire N__39904;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39896;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39880;
    wire N__39877;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39855;
    wire N__39850;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39840;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39825;
    wire N__39820;
    wire N__39817;
    wire N__39816;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39802;
    wire N__39799;
    wire N__39798;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39783;
    wire N__39778;
    wire N__39775;
    wire N__39772;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39757;
    wire N__39754;
    wire N__39753;
    wire N__39752;
    wire N__39749;
    wire N__39746;
    wire N__39743;
    wire N__39738;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39726;
    wire N__39723;
    wire N__39720;
    wire N__39719;
    wire N__39714;
    wire N__39711;
    wire N__39708;
    wire N__39703;
    wire N__39700;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39688;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39673;
    wire N__39670;
    wire N__39667;
    wire N__39666;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39651;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39636;
    wire N__39635;
    wire N__39632;
    wire N__39629;
    wire N__39626;
    wire N__39621;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39606;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39591;
    wire N__39586;
    wire N__39583;
    wire N__39582;
    wire N__39581;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39565;
    wire N__39562;
    wire N__39561;
    wire N__39560;
    wire N__39555;
    wire N__39552;
    wire N__39549;
    wire N__39544;
    wire N__39541;
    wire N__39540;
    wire N__39537;
    wire N__39534;
    wire N__39533;
    wire N__39528;
    wire N__39525;
    wire N__39522;
    wire N__39517;
    wire N__39514;
    wire N__39513;
    wire N__39508;
    wire N__39507;
    wire N__39504;
    wire N__39501;
    wire N__39498;
    wire N__39493;
    wire N__39490;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39482;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39466;
    wire N__39463;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39451;
    wire N__39450;
    wire N__39447;
    wire N__39444;
    wire N__39441;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39422;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39399;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39384;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39370;
    wire N__39369;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39359;
    wire N__39354;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39342;
    wire N__39339;
    wire N__39336;
    wire N__39335;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39319;
    wire N__39316;
    wire N__39315;
    wire N__39310;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39295;
    wire N__39292;
    wire N__39291;
    wire N__39286;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39271;
    wire N__39268;
    wire N__39265;
    wire N__39262;
    wire N__39259;
    wire N__39256;
    wire N__39253;
    wire N__39250;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39238;
    wire N__39237;
    wire N__39234;
    wire N__39231;
    wire N__39228;
    wire N__39223;
    wire N__39220;
    wire N__39219;
    wire N__39216;
    wire N__39213;
    wire N__39210;
    wire N__39209;
    wire N__39204;
    wire N__39201;
    wire N__39198;
    wire N__39193;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39181;
    wire N__39178;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39145;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39135;
    wire N__39134;
    wire N__39131;
    wire N__39126;
    wire N__39121;
    wire N__39120;
    wire N__39115;
    wire N__39112;
    wire N__39111;
    wire N__39110;
    wire N__39107;
    wire N__39102;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39088;
    wire N__39085;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39048;
    wire N__39047;
    wire N__39044;
    wire N__39039;
    wire N__39034;
    wire N__39033;
    wire N__39028;
    wire N__39025;
    wire N__39024;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39009;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38994;
    wire N__38989;
    wire N__38986;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38976;
    wire N__38971;
    wire N__38968;
    wire N__38967;
    wire N__38966;
    wire N__38963;
    wire N__38958;
    wire N__38953;
    wire N__38952;
    wire N__38951;
    wire N__38948;
    wire N__38945;
    wire N__38942;
    wire N__38937;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38919;
    wire N__38914;
    wire N__38911;
    wire N__38908;
    wire N__38905;
    wire N__38902;
    wire N__38901;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38886;
    wire N__38883;
    wire N__38878;
    wire N__38875;
    wire N__38872;
    wire N__38871;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38859;
    wire N__38854;
    wire N__38853;
    wire N__38852;
    wire N__38849;
    wire N__38844;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38824;
    wire N__38821;
    wire N__38818;
    wire N__38817;
    wire N__38816;
    wire N__38813;
    wire N__38812;
    wire N__38809;
    wire N__38808;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38798;
    wire N__38791;
    wire N__38786;
    wire N__38779;
    wire N__38776;
    wire N__38775;
    wire N__38772;
    wire N__38769;
    wire N__38764;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38752;
    wire N__38751;
    wire N__38748;
    wire N__38745;
    wire N__38742;
    wire N__38737;
    wire N__38736;
    wire N__38735;
    wire N__38732;
    wire N__38727;
    wire N__38722;
    wire N__38721;
    wire N__38720;
    wire N__38717;
    wire N__38714;
    wire N__38711;
    wire N__38706;
    wire N__38701;
    wire N__38698;
    wire N__38695;
    wire N__38692;
    wire N__38691;
    wire N__38686;
    wire N__38683;
    wire N__38682;
    wire N__38677;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38647;
    wire N__38644;
    wire N__38641;
    wire N__38638;
    wire N__38635;
    wire N__38632;
    wire N__38629;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38611;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38593;
    wire N__38590;
    wire N__38587;
    wire N__38586;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38572;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38562;
    wire N__38559;
    wire N__38556;
    wire N__38553;
    wire N__38548;
    wire N__38545;
    wire N__38542;
    wire N__38539;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38515;
    wire N__38514;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38478;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38446;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38434;
    wire N__38431;
    wire N__38428;
    wire N__38425;
    wire N__38422;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38412;
    wire N__38407;
    wire N__38404;
    wire N__38401;
    wire N__38398;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38373;
    wire N__38370;
    wire N__38367;
    wire N__38364;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38287;
    wire N__38284;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38262;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38247;
    wire N__38244;
    wire N__38241;
    wire N__38238;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38161;
    wire N__38158;
    wire N__38155;
    wire N__38154;
    wire N__38151;
    wire N__38150;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38136;
    wire N__38131;
    wire N__38128;
    wire N__38127;
    wire N__38126;
    wire N__38123;
    wire N__38118;
    wire N__38115;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38071;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37918;
    wire N__37915;
    wire N__37912;
    wire N__37909;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37893;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37879;
    wire N__37878;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37864;
    wire N__37861;
    wire N__37858;
    wire N__37855;
    wire N__37852;
    wire N__37849;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37828;
    wire N__37825;
    wire N__37822;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37807;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37788;
    wire N__37785;
    wire N__37782;
    wire N__37779;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37758;
    wire N__37753;
    wire N__37750;
    wire N__37749;
    wire N__37744;
    wire N__37741;
    wire N__37740;
    wire N__37735;
    wire N__37732;
    wire N__37731;
    wire N__37728;
    wire N__37723;
    wire N__37720;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37700;
    wire N__37697;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37672;
    wire N__37671;
    wire N__37668;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37658;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37633;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37597;
    wire N__37594;
    wire N__37585;
    wire N__37584;
    wire N__37581;
    wire N__37580;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37561;
    wire N__37558;
    wire N__37555;
    wire N__37552;
    wire N__37543;
    wire N__37540;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37513;
    wire N__37510;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37462;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37444;
    wire N__37441;
    wire N__37438;
    wire N__37435;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37420;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37405;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37390;
    wire N__37387;
    wire N__37384;
    wire N__37381;
    wire N__37378;
    wire N__37375;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37360;
    wire N__37357;
    wire N__37354;
    wire N__37351;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37327;
    wire N__37324;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37297;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37273;
    wire N__37270;
    wire N__37267;
    wire N__37264;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37210;
    wire N__37207;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37183;
    wire N__37180;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37165;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37041;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36970;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36943;
    wire N__36940;
    wire N__36939;
    wire N__36938;
    wire N__36937;
    wire N__36936;
    wire N__36935;
    wire N__36934;
    wire N__36933;
    wire N__36932;
    wire N__36931;
    wire N__36930;
    wire N__36929;
    wire N__36928;
    wire N__36927;
    wire N__36926;
    wire N__36925;
    wire N__36924;
    wire N__36923;
    wire N__36922;
    wire N__36921;
    wire N__36920;
    wire N__36919;
    wire N__36918;
    wire N__36917;
    wire N__36916;
    wire N__36915;
    wire N__36914;
    wire N__36913;
    wire N__36912;
    wire N__36911;
    wire N__36910;
    wire N__36909;
    wire N__36900;
    wire N__36891;
    wire N__36882;
    wire N__36875;
    wire N__36866;
    wire N__36857;
    wire N__36848;
    wire N__36837;
    wire N__36820;
    wire N__36817;
    wire N__36816;
    wire N__36815;
    wire N__36814;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36799;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36781;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36772;
    wire N__36771;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36757;
    wire N__36754;
    wire N__36751;
    wire N__36742;
    wire N__36741;
    wire N__36740;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36728;
    wire N__36725;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36703;
    wire N__36700;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36677;
    wire N__36674;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36640;
    wire N__36637;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36625;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36617;
    wire N__36616;
    wire N__36611;
    wire N__36608;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36595;
    wire N__36594;
    wire N__36593;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36565;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36553;
    wire N__36550;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36515;
    wire N__36512;
    wire N__36509;
    wire N__36502;
    wire N__36499;
    wire N__36498;
    wire N__36497;
    wire N__36496;
    wire N__36493;
    wire N__36486;
    wire N__36483;
    wire N__36478;
    wire N__36477;
    wire N__36476;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36421;
    wire N__36418;
    wire N__36409;
    wire N__36406;
    wire N__36405;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36395;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36376;
    wire N__36375;
    wire N__36374;
    wire N__36371;
    wire N__36366;
    wire N__36361;
    wire N__36358;
    wire N__36357;
    wire N__36356;
    wire N__36355;
    wire N__36354;
    wire N__36353;
    wire N__36346;
    wire N__36339;
    wire N__36334;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36307;
    wire N__36304;
    wire N__36301;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36293;
    wire N__36292;
    wire N__36289;
    wire N__36286;
    wire N__36281;
    wire N__36274;
    wire N__36273;
    wire N__36272;
    wire N__36269;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36257;
    wire N__36250;
    wire N__36249;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36213;
    wire N__36210;
    wire N__36209;
    wire N__36206;
    wire N__36205;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36172;
    wire N__36169;
    wire N__36166;
    wire N__36165;
    wire N__36164;
    wire N__36161;
    wire N__36156;
    wire N__36151;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36143;
    wire N__36138;
    wire N__36133;
    wire N__36130;
    wire N__36129;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36105;
    wire N__36104;
    wire N__36101;
    wire N__36096;
    wire N__36091;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36078;
    wire N__36077;
    wire N__36072;
    wire N__36069;
    wire N__36066;
    wire N__36061;
    wire N__36058;
    wire N__36057;
    wire N__36054;
    wire N__36051;
    wire N__36046;
    wire N__36045;
    wire N__36042;
    wire N__36039;
    wire N__36036;
    wire N__36031;
    wire N__36028;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35989;
    wire N__35986;
    wire N__35983;
    wire N__35982;
    wire N__35977;
    wire N__35974;
    wire N__35971;
    wire N__35968;
    wire N__35965;
    wire N__35962;
    wire N__35959;
    wire N__35956;
    wire N__35953;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35942;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35932;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35913;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35898;
    wire N__35897;
    wire N__35894;
    wire N__35893;
    wire N__35890;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35876;
    wire N__35869;
    wire N__35866;
    wire N__35865;
    wire N__35864;
    wire N__35863;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35858;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35852;
    wire N__35845;
    wire N__35842;
    wire N__35833;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35825;
    wire N__35824;
    wire N__35823;
    wire N__35822;
    wire N__35821;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35817;
    wire N__35816;
    wire N__35815;
    wire N__35814;
    wire N__35813;
    wire N__35812;
    wire N__35811;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35792;
    wire N__35789;
    wire N__35774;
    wire N__35771;
    wire N__35762;
    wire N__35749;
    wire N__35744;
    wire N__35737;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35672;
    wire N__35665;
    wire N__35662;
    wire N__35659;
    wire N__35656;
    wire N__35653;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35645;
    wire N__35644;
    wire N__35639;
    wire N__35636;
    wire N__35633;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35616;
    wire N__35613;
    wire N__35612;
    wire N__35611;
    wire N__35608;
    wire N__35605;
    wire N__35602;
    wire N__35597;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35577;
    wire N__35576;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35564;
    wire N__35557;
    wire N__35554;
    wire N__35551;
    wire N__35548;
    wire N__35547;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35537;
    wire N__35536;
    wire N__35531;
    wire N__35526;
    wire N__35521;
    wire N__35518;
    wire N__35515;
    wire N__35514;
    wire N__35511;
    wire N__35508;
    wire N__35505;
    wire N__35504;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35462;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35394;
    wire N__35391;
    wire N__35388;
    wire N__35383;
    wire N__35380;
    wire N__35377;
    wire N__35374;
    wire N__35371;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35363;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35331;
    wire N__35326;
    wire N__35323;
    wire N__35320;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35307;
    wire N__35304;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35278;
    wire N__35275;
    wire N__35272;
    wire N__35269;
    wire N__35266;
    wire N__35265;
    wire N__35262;
    wire N__35261;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35248;
    wire N__35245;
    wire N__35240;
    wire N__35237;
    wire N__35232;
    wire N__35229;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35202;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35150;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35094;
    wire N__35091;
    wire N__35090;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35080;
    wire N__35077;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35052;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35042;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34998;
    wire N__34997;
    wire N__34994;
    wire N__34991;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34971;
    wire N__34966;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34950;
    wire N__34947;
    wire N__34946;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34936;
    wire N__34933;
    wire N__34924;
    wire N__34921;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34913;
    wire N__34910;
    wire N__34909;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34888;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34861;
    wire N__34860;
    wire N__34859;
    wire N__34856;
    wire N__34855;
    wire N__34852;
    wire N__34849;
    wire N__34846;
    wire N__34843;
    wire N__34840;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34824;
    wire N__34823;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34810;
    wire N__34803;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34780;
    wire N__34777;
    wire N__34774;
    wire N__34771;
    wire N__34770;
    wire N__34767;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34759;
    wire N__34756;
    wire N__34753;
    wire N__34750;
    wire N__34747;
    wire N__34744;
    wire N__34741;
    wire N__34732;
    wire N__34729;
    wire N__34726;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34701;
    wire N__34698;
    wire N__34697;
    wire N__34694;
    wire N__34693;
    wire N__34690;
    wire N__34685;
    wire N__34682;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34657;
    wire N__34656;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34624;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34585;
    wire N__34582;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34558;
    wire N__34557;
    wire N__34556;
    wire N__34553;
    wire N__34548;
    wire N__34543;
    wire N__34542;
    wire N__34541;
    wire N__34538;
    wire N__34533;
    wire N__34528;
    wire N__34525;
    wire N__34522;
    wire N__34519;
    wire N__34516;
    wire N__34513;
    wire N__34510;
    wire N__34507;
    wire N__34504;
    wire N__34503;
    wire N__34502;
    wire N__34499;
    wire N__34494;
    wire N__34489;
    wire N__34486;
    wire N__34485;
    wire N__34484;
    wire N__34483;
    wire N__34474;
    wire N__34471;
    wire N__34470;
    wire N__34469;
    wire N__34466;
    wire N__34461;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34444;
    wire N__34441;
    wire N__34440;
    wire N__34437;
    wire N__34436;
    wire N__34435;
    wire N__34434;
    wire N__34431;
    wire N__34430;
    wire N__34427;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34399;
    wire N__34398;
    wire N__34397;
    wire N__34396;
    wire N__34395;
    wire N__34392;
    wire N__34387;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34368;
    wire N__34363;
    wire N__34360;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34335;
    wire N__34330;
    wire N__34327;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34315;
    wire N__34312;
    wire N__34311;
    wire N__34310;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34291;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34270;
    wire N__34267;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34255;
    wire N__34254;
    wire N__34251;
    wire N__34248;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34183;
    wire N__34180;
    wire N__34177;
    wire N__34174;
    wire N__34171;
    wire N__34168;
    wire N__34167;
    wire N__34164;
    wire N__34161;
    wire N__34156;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34137;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34123;
    wire N__34120;
    wire N__34117;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34096;
    wire N__34093;
    wire N__34090;
    wire N__34087;
    wire N__34084;
    wire N__34081;
    wire N__34078;
    wire N__34077;
    wire N__34076;
    wire N__34073;
    wire N__34068;
    wire N__34063;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34055;
    wire N__34052;
    wire N__34047;
    wire N__34044;
    wire N__34039;
    wire N__34036;
    wire N__34035;
    wire N__34034;
    wire N__34033;
    wire N__34032;
    wire N__34029;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34009;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33990;
    wire N__33989;
    wire N__33986;
    wire N__33981;
    wire N__33976;
    wire N__33973;
    wire N__33972;
    wire N__33969;
    wire N__33968;
    wire N__33965;
    wire N__33960;
    wire N__33955;
    wire N__33952;
    wire N__33951;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33937;
    wire N__33934;
    wire N__33933;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33919;
    wire N__33916;
    wire N__33913;
    wire N__33912;
    wire N__33911;
    wire N__33910;
    wire N__33901;
    wire N__33898;
    wire N__33897;
    wire N__33896;
    wire N__33893;
    wire N__33888;
    wire N__33883;
    wire N__33882;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33865;
    wire N__33862;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33817;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33796;
    wire N__33793;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33778;
    wire N__33777;
    wire N__33776;
    wire N__33773;
    wire N__33772;
    wire N__33771;
    wire N__33770;
    wire N__33769;
    wire N__33768;
    wire N__33767;
    wire N__33762;
    wire N__33759;
    wire N__33754;
    wire N__33753;
    wire N__33752;
    wire N__33751;
    wire N__33750;
    wire N__33749;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33730;
    wire N__33729;
    wire N__33728;
    wire N__33727;
    wire N__33726;
    wire N__33725;
    wire N__33724;
    wire N__33723;
    wire N__33714;
    wire N__33711;
    wire N__33710;
    wire N__33709;
    wire N__33704;
    wire N__33699;
    wire N__33696;
    wire N__33695;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33691;
    wire N__33686;
    wire N__33683;
    wire N__33682;
    wire N__33681;
    wire N__33672;
    wire N__33667;
    wire N__33662;
    wire N__33659;
    wire N__33654;
    wire N__33649;
    wire N__33642;
    wire N__33639;
    wire N__33632;
    wire N__33627;
    wire N__33610;
    wire N__33607;
    wire N__33604;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33570;
    wire N__33565;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33544;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33532;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33484;
    wire N__33483;
    wire N__33478;
    wire N__33475;
    wire N__33474;
    wire N__33473;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33457;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33445;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33430;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33414;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33393;
    wire N__33392;
    wire N__33389;
    wire N__33384;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33374;
    wire N__33369;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33348;
    wire N__33343;
    wire N__33340;
    wire N__33339;
    wire N__33334;
    wire N__33331;
    wire N__33330;
    wire N__33325;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33319;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33279;
    wire N__33274;
    wire N__33271;
    wire N__33270;
    wire N__33265;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33238;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33213;
    wire N__33208;
    wire N__33205;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33190;
    wire N__33189;
    wire N__33186;
    wire N__33185;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33171;
    wire N__33166;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33140;
    wire N__33137;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33109;
    wire N__33108;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33025;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32950;
    wire N__32947;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32926;
    wire N__32925;
    wire N__32924;
    wire N__32919;
    wire N__32918;
    wire N__32917;
    wire N__32916;
    wire N__32915;
    wire N__32914;
    wire N__32913;
    wire N__32912;
    wire N__32911;
    wire N__32910;
    wire N__32909;
    wire N__32908;
    wire N__32907;
    wire N__32906;
    wire N__32905;
    wire N__32904;
    wire N__32903;
    wire N__32902;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32883;
    wire N__32882;
    wire N__32881;
    wire N__32880;
    wire N__32879;
    wire N__32878;
    wire N__32877;
    wire N__32874;
    wire N__32871;
    wire N__32858;
    wire N__32843;
    wire N__32838;
    wire N__32835;
    wire N__32830;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32814;
    wire N__32811;
    wire N__32808;
    wire N__32803;
    wire N__32796;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32755;
    wire N__32754;
    wire N__32751;
    wire N__32748;
    wire N__32743;
    wire N__32742;
    wire N__32741;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32725;
    wire N__32724;
    wire N__32719;
    wire N__32716;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32708;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32692;
    wire N__32689;
    wire N__32686;
    wire N__32683;
    wire N__32680;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32668;
    wire N__32667;
    wire N__32662;
    wire N__32659;
    wire N__32658;
    wire N__32657;
    wire N__32656;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32623;
    wire N__32620;
    wire N__32619;
    wire N__32616;
    wire N__32615;
    wire N__32612;
    wire N__32609;
    wire N__32606;
    wire N__32603;
    wire N__32600;
    wire N__32597;
    wire N__32596;
    wire N__32593;
    wire N__32582;
    wire N__32579;
    wire N__32576;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32560;
    wire N__32557;
    wire N__32556;
    wire N__32555;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32545;
    wire N__32544;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32530;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32516;
    wire N__32509;
    wire N__32508;
    wire N__32507;
    wire N__32506;
    wire N__32505;
    wire N__32504;
    wire N__32503;
    wire N__32502;
    wire N__32501;
    wire N__32500;
    wire N__32499;
    wire N__32498;
    wire N__32497;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32493;
    wire N__32492;
    wire N__32491;
    wire N__32490;
    wire N__32489;
    wire N__32488;
    wire N__32487;
    wire N__32486;
    wire N__32485;
    wire N__32484;
    wire N__32483;
    wire N__32482;
    wire N__32481;
    wire N__32480;
    wire N__32479;
    wire N__32478;
    wire N__32471;
    wire N__32462;
    wire N__32453;
    wire N__32442;
    wire N__32433;
    wire N__32424;
    wire N__32415;
    wire N__32406;
    wire N__32403;
    wire N__32398;
    wire N__32395;
    wire N__32390;
    wire N__32381;
    wire N__32374;
    wire N__32371;
    wire N__32368;
    wire N__32367;
    wire N__32362;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32335;
    wire N__32334;
    wire N__32333;
    wire N__32332;
    wire N__32331;
    wire N__32330;
    wire N__32329;
    wire N__32328;
    wire N__32327;
    wire N__32326;
    wire N__32325;
    wire N__32324;
    wire N__32323;
    wire N__32322;
    wire N__32321;
    wire N__32320;
    wire N__32319;
    wire N__32318;
    wire N__32317;
    wire N__32316;
    wire N__32315;
    wire N__32314;
    wire N__32313;
    wire N__32312;
    wire N__32303;
    wire N__32294;
    wire N__32285;
    wire N__32276;
    wire N__32275;
    wire N__32274;
    wire N__32273;
    wire N__32272;
    wire N__32271;
    wire N__32270;
    wire N__32269;
    wire N__32268;
    wire N__32259;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32229;
    wire N__32220;
    wire N__32215;
    wire N__32210;
    wire N__32205;
    wire N__32194;
    wire N__32191;
    wire N__32190;
    wire N__32189;
    wire N__32188;
    wire N__32179;
    wire N__32176;
    wire N__32173;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32143;
    wire N__32142;
    wire N__32137;
    wire N__32134;
    wire N__32133;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32114;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32098;
    wire N__32097;
    wire N__32096;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32080;
    wire N__32077;
    wire N__32074;
    wire N__32071;
    wire N__32068;
    wire N__32067;
    wire N__32066;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32050;
    wire N__32047;
    wire N__32046;
    wire N__32045;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32013;
    wire N__32008;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31993;
    wire N__31990;
    wire N__31989;
    wire N__31984;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31969;
    wire N__31966;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31954;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31918;
    wire N__31915;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31903;
    wire N__31900;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31888;
    wire N__31885;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31873;
    wire N__31870;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31858;
    wire N__31855;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31843;
    wire N__31840;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31828;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31813;
    wire N__31810;
    wire N__31809;
    wire N__31804;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31789;
    wire N__31786;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31774;
    wire N__31771;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31759;
    wire N__31756;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31744;
    wire N__31741;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31729;
    wire N__31726;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31711;
    wire N__31708;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31696;
    wire N__31693;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31678;
    wire N__31675;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31663;
    wire N__31660;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31639;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31623;
    wire N__31622;
    wire N__31621;
    wire N__31620;
    wire N__31619;
    wire N__31618;
    wire N__31617;
    wire N__31616;
    wire N__31615;
    wire N__31614;
    wire N__31613;
    wire N__31612;
    wire N__31611;
    wire N__31610;
    wire N__31609;
    wire N__31608;
    wire N__31607;
    wire N__31606;
    wire N__31605;
    wire N__31604;
    wire N__31603;
    wire N__31602;
    wire N__31601;
    wire N__31600;
    wire N__31599;
    wire N__31598;
    wire N__31597;
    wire N__31590;
    wire N__31579;
    wire N__31578;
    wire N__31577;
    wire N__31576;
    wire N__31575;
    wire N__31566;
    wire N__31557;
    wire N__31548;
    wire N__31539;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31515;
    wire N__31500;
    wire N__31495;
    wire N__31492;
    wire N__31491;
    wire N__31490;
    wire N__31489;
    wire N__31486;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31460;
    wire N__31457;
    wire N__31452;
    wire N__31447;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31432;
    wire N__31429;
    wire N__31426;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31414;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31401;
    wire N__31400;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31384;
    wire N__31381;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31373;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31357;
    wire N__31354;
    wire N__31353;
    wire N__31350;
    wire N__31345;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31330;
    wire N__31327;
    wire N__31326;
    wire N__31323;
    wire N__31318;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31261;
    wire N__31258;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31243;
    wire N__31240;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31225;
    wire N__31222;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31207;
    wire N__31204;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31189;
    wire N__31186;
    wire N__31183;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31168;
    wire N__31165;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31150;
    wire N__31147;
    wire N__31144;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31129;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31116;
    wire N__31113;
    wire N__31110;
    wire N__31107;
    wire N__31102;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31087;
    wire N__31084;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31069;
    wire N__31066;
    wire N__31065;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31051;
    wire N__31048;
    wire N__31047;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31027;
    wire N__31024;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31009;
    wire N__31006;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30991;
    wire N__30988;
    wire N__30987;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30973;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30958;
    wire N__30955;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30938;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30922;
    wire N__30919;
    wire N__30916;
    wire N__30913;
    wire N__30910;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30808;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30781;
    wire N__30778;
    wire N__30775;
    wire N__30774;
    wire N__30773;
    wire N__30772;
    wire N__30771;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30766;
    wire N__30765;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30749;
    wire N__30746;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30728;
    wire N__30725;
    wire N__30718;
    wire N__30709;
    wire N__30704;
    wire N__30699;
    wire N__30696;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30580;
    wire N__30577;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30550;
    wire N__30547;
    wire N__30544;
    wire N__30541;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30445;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30385;
    wire N__30382;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30355;
    wire N__30352;
    wire N__30349;
    wire N__30346;
    wire N__30343;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30298;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30255;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30202;
    wire N__30199;
    wire N__30196;
    wire N__30193;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30172;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30130;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30106;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30091;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30076;
    wire N__30073;
    wire N__30070;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30058;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30043;
    wire N__30042;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30028;
    wire N__30025;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30004;
    wire N__30003;
    wire N__30000;
    wire N__29997;
    wire N__29992;
    wire N__29989;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29971;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29914;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29901;
    wire N__29898;
    wire N__29895;
    wire N__29890;
    wire N__29887;
    wire N__29884;
    wire N__29881;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29863;
    wire N__29860;
    wire N__29857;
    wire N__29854;
    wire N__29851;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29839;
    wire N__29836;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29828;
    wire N__29825;
    wire N__29822;
    wire N__29819;
    wire N__29812;
    wire N__29809;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29794;
    wire N__29791;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29783;
    wire N__29780;
    wire N__29777;
    wire N__29774;
    wire N__29767;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29752;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29740;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29728;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29653;
    wire N__29652;
    wire N__29651;
    wire N__29648;
    wire N__29643;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29584;
    wire N__29581;
    wire N__29578;
    wire N__29575;
    wire N__29572;
    wire N__29569;
    wire N__29566;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29551;
    wire N__29548;
    wire N__29545;
    wire N__29542;
    wire N__29539;
    wire N__29536;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29524;
    wire N__29523;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29466;
    wire N__29465;
    wire N__29462;
    wire N__29459;
    wire N__29456;
    wire N__29451;
    wire N__29446;
    wire N__29443;
    wire N__29442;
    wire N__29441;
    wire N__29438;
    wire N__29433;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29409;
    wire N__29406;
    wire N__29405;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29390;
    wire N__29387;
    wire N__29380;
    wire N__29377;
    wire N__29376;
    wire N__29375;
    wire N__29372;
    wire N__29367;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29331;
    wire N__29328;
    wire N__29327;
    wire N__29324;
    wire N__29323;
    wire N__29320;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29302;
    wire N__29299;
    wire N__29298;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29286;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29268;
    wire N__29267;
    wire N__29266;
    wire N__29265;
    wire N__29264;
    wire N__29261;
    wire N__29258;
    wire N__29255;
    wire N__29248;
    wire N__29239;
    wire N__29238;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29158;
    wire N__29155;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29137;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29068;
    wire N__29065;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28969;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28957;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28939;
    wire N__28936;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28915;
    wire N__28912;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28900;
    wire N__28897;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28882;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28834;
    wire N__28831;
    wire N__28828;
    wire N__28825;
    wire N__28822;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28810;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28789;
    wire N__28786;
    wire N__28783;
    wire N__28780;
    wire N__28777;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28762;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28726;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28714;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28669;
    wire N__28668;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28645;
    wire N__28644;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28621;
    wire N__28620;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28558;
    wire N__28555;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28504;
    wire N__28501;
    wire N__28498;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28444;
    wire N__28441;
    wire N__28438;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28414;
    wire N__28413;
    wire N__28412;
    wire N__28411;
    wire N__28410;
    wire N__28409;
    wire N__28406;
    wire N__28405;
    wire N__28402;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28388;
    wire N__28385;
    wire N__28376;
    wire N__28373;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28355;
    wire N__28352;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28264;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28156;
    wire N__28153;
    wire N__28150;
    wire N__28147;
    wire N__28144;
    wire N__28141;
    wire N__28138;
    wire N__28135;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28066;
    wire N__28063;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28012;
    wire N__28009;
    wire N__28006;
    wire N__28003;
    wire N__28000;
    wire N__27997;
    wire N__27994;
    wire N__27991;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27979;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27913;
    wire N__27910;
    wire N__27909;
    wire N__27906;
    wire N__27903;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27885;
    wire N__27882;
    wire N__27879;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27847;
    wire N__27844;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27822;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27799;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27786;
    wire N__27781;
    wire N__27778;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27763;
    wire N__27760;
    wire N__27757;
    wire N__27754;
    wire N__27751;
    wire N__27748;
    wire N__27745;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27735;
    wire N__27730;
    wire N__27727;
    wire N__27724;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27712;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27604;
    wire N__27601;
    wire N__27600;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27580;
    wire N__27577;
    wire N__27574;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27562;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27550;
    wire N__27547;
    wire N__27544;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27499;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27478;
    wire N__27475;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27463;
    wire N__27460;
    wire N__27457;
    wire N__27454;
    wire N__27451;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27424;
    wire N__27421;
    wire N__27418;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27283;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27232;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27177;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27160;
    wire N__27157;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27135;
    wire N__27130;
    wire N__27127;
    wire N__27126;
    wire N__27123;
    wire N__27120;
    wire N__27115;
    wire N__27112;
    wire N__27109;
    wire N__27106;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27094;
    wire N__27091;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27079;
    wire N__27076;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27043;
    wire N__27040;
    wire N__27037;
    wire N__27034;
    wire N__27031;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27019;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26980;
    wire N__26977;
    wire N__26976;
    wire N__26971;
    wire N__26968;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26956;
    wire N__26953;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26941;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26923;
    wire N__26922;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26899;
    wire N__26896;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26886;
    wire N__26883;
    wire N__26878;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26870;
    wire N__26869;
    wire N__26862;
    wire N__26859;
    wire N__26854;
    wire N__26851;
    wire N__26848;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26797;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26782;
    wire N__26779;
    wire N__26776;
    wire N__26773;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26689;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26668;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26620;
    wire N__26617;
    wire N__26614;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26602;
    wire N__26599;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26587;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26566;
    wire N__26563;
    wire N__26560;
    wire N__26557;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26491;
    wire N__26488;
    wire N__26485;
    wire N__26482;
    wire N__26479;
    wire N__26476;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26457;
    wire N__26452;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26437;
    wire N__26434;
    wire N__26433;
    wire N__26430;
    wire N__26427;
    wire N__26422;
    wire N__26421;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26407;
    wire N__26404;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26392;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26377;
    wire N__26374;
    wire N__26373;
    wire N__26368;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26353;
    wire N__26350;
    wire N__26349;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26332;
    wire N__26329;
    wire N__26328;
    wire N__26327;
    wire N__26324;
    wire N__26319;
    wire N__26314;
    wire N__26311;
    wire N__26310;
    wire N__26309;
    wire N__26306;
    wire N__26301;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26289;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26272;
    wire N__26271;
    wire N__26270;
    wire N__26269;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26253;
    wire N__26250;
    wire N__26247;
    wire N__26242;
    wire N__26239;
    wire N__26238;
    wire N__26233;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26218;
    wire N__26215;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26203;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26179;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26169;
    wire N__26164;
    wire N__26161;
    wire N__26160;
    wire N__26155;
    wire N__26154;
    wire N__26151;
    wire N__26148;
    wire N__26145;
    wire N__26140;
    wire N__26137;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26129;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26113;
    wire N__26110;
    wire N__26109;
    wire N__26108;
    wire N__26103;
    wire N__26100;
    wire N__26097;
    wire N__26092;
    wire N__26089;
    wire N__26088;
    wire N__26085;
    wire N__26082;
    wire N__26077;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26062;
    wire N__26059;
    wire N__26058;
    wire N__26053;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26038;
    wire N__26035;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26023;
    wire N__26020;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26008;
    wire N__26005;
    wire N__26004;
    wire N__26001;
    wire N__25998;
    wire N__25993;
    wire N__25990;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25978;
    wire N__25975;
    wire N__25974;
    wire N__25971;
    wire N__25968;
    wire N__25963;
    wire N__25960;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25948;
    wire N__25945;
    wire N__25944;
    wire N__25941;
    wire N__25938;
    wire N__25933;
    wire N__25930;
    wire N__25929;
    wire N__25926;
    wire N__25923;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25911;
    wire N__25908;
    wire N__25905;
    wire N__25902;
    wire N__25897;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25882;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25870;
    wire N__25867;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25840;
    wire N__25837;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25825;
    wire N__25822;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25810;
    wire N__25807;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25761;
    wire N__25758;
    wire N__25755;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25741;
    wire N__25738;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25708;
    wire N__25705;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25663;
    wire N__25660;
    wire N__25657;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25558;
    wire N__25555;
    wire N__25552;
    wire N__25549;
    wire N__25548;
    wire N__25547;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25531;
    wire N__25528;
    wire N__25525;
    wire N__25524;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25500;
    wire N__25499;
    wire N__25496;
    wire N__25493;
    wire N__25490;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25476;
    wire N__25475;
    wire N__25472;
    wire N__25469;
    wire N__25466;
    wire N__25459;
    wire N__25456;
    wire N__25453;
    wire N__25452;
    wire N__25451;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25428;
    wire N__25427;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25411;
    wire N__25408;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25396;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25382;
    wire N__25375;
    wire N__25372;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25360;
    wire N__25357;
    wire N__25356;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25330;
    wire N__25329;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25312;
    wire N__25309;
    wire N__25306;
    wire N__25305;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25281;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25264;
    wire N__25261;
    wire N__25258;
    wire N__25257;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25240;
    wire N__25237;
    wire N__25234;
    wire N__25233;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25216;
    wire N__25213;
    wire N__25212;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25188;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25178;
    wire N__25171;
    wire N__25168;
    wire N__25167;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25152;
    wire N__25147;
    wire N__25144;
    wire N__25141;
    wire N__25140;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25125;
    wire N__25120;
    wire N__25117;
    wire N__25114;
    wire N__25113;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25089;
    wire N__25088;
    wire N__25085;
    wire N__25082;
    wire N__25079;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25065;
    wire N__25064;
    wire N__25061;
    wire N__25058;
    wire N__25055;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25041;
    wire N__25040;
    wire N__25037;
    wire N__25034;
    wire N__25031;
    wire N__25024;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25016;
    wire N__25013;
    wire N__25010;
    wire N__25003;
    wire N__25000;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24979;
    wire N__24976;
    wire N__24975;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24960;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24903;
    wire N__24902;
    wire N__24899;
    wire N__24894;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24882;
    wire N__24881;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24865;
    wire N__24862;
    wire N__24859;
    wire N__24856;
    wire N__24853;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24799;
    wire N__24796;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24721;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24559;
    wire N__24556;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24502;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24457;
    wire N__24454;
    wire N__24451;
    wire N__24448;
    wire N__24445;
    wire N__24444;
    wire N__24439;
    wire N__24436;
    wire N__24435;
    wire N__24430;
    wire N__24427;
    wire N__24426;
    wire N__24421;
    wire N__24418;
    wire N__24417;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24372;
    wire N__24371;
    wire N__24370;
    wire N__24369;
    wire N__24368;
    wire N__24367;
    wire N__24366;
    wire N__24365;
    wire N__24364;
    wire N__24363;
    wire N__24362;
    wire N__24361;
    wire N__24360;
    wire N__24359;
    wire N__24358;
    wire N__24357;
    wire N__24356;
    wire N__24355;
    wire N__24354;
    wire N__24353;
    wire N__24352;
    wire N__24343;
    wire N__24342;
    wire N__24341;
    wire N__24340;
    wire N__24339;
    wire N__24338;
    wire N__24337;
    wire N__24336;
    wire N__24335;
    wire N__24330;
    wire N__24321;
    wire N__24312;
    wire N__24303;
    wire N__24294;
    wire N__24291;
    wire N__24282;
    wire N__24273;
    wire N__24268;
    wire N__24257;
    wire N__24254;
    wire N__24249;
    wire N__24244;
    wire N__24241;
    wire N__24238;
    wire N__24235;
    wire N__24232;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24216;
    wire N__24213;
    wire N__24210;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24193;
    wire N__24190;
    wire N__24187;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24175;
    wire N__24172;
    wire N__24169;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24148;
    wire N__24145;
    wire N__24142;
    wire N__24139;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24120;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24108;
    wire N__24103;
    wire N__24100;
    wire N__24097;
    wire N__24096;
    wire N__24091;
    wire N__24088;
    wire N__24085;
    wire N__24084;
    wire N__24079;
    wire N__24076;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24057;
    wire N__24052;
    wire N__24049;
    wire N__24048;
    wire N__24043;
    wire N__24040;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24028;
    wire N__24025;
    wire N__24024;
    wire N__24019;
    wire N__24016;
    wire N__24015;
    wire N__24010;
    wire N__24007;
    wire N__24006;
    wire N__24001;
    wire N__23998;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23986;
    wire N__23983;
    wire N__23982;
    wire N__23977;
    wire N__23974;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23963;
    wire N__23956;
    wire N__23953;
    wire N__23952;
    wire N__23951;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23935;
    wire N__23932;
    wire N__23931;
    wire N__23930;
    wire N__23927;
    wire N__23924;
    wire N__23921;
    wire N__23914;
    wire N__23911;
    wire N__23910;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23893;
    wire N__23890;
    wire N__23889;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23869;
    wire N__23866;
    wire N__23865;
    wire N__23864;
    wire N__23863;
    wire N__23862;
    wire N__23861;
    wire N__23860;
    wire N__23859;
    wire N__23858;
    wire N__23857;
    wire N__23852;
    wire N__23843;
    wire N__23834;
    wire N__23831;
    wire N__23824;
    wire N__23821;
    wire N__23820;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23760;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23743;
    wire N__23740;
    wire N__23739;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23722;
    wire N__23719;
    wire N__23718;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23696;
    wire N__23693;
    wire N__23690;
    wire N__23687;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23569;
    wire N__23566;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23482;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23470;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23458;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23448;
    wire N__23445;
    wire N__23440;
    wire N__23439;
    wire N__23436;
    wire N__23433;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23395;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23391;
    wire N__23388;
    wire N__23387;
    wire N__23386;
    wire N__23385;
    wire N__23384;
    wire N__23383;
    wire N__23380;
    wire N__23375;
    wire N__23368;
    wire N__23359;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23332;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23302;
    wire N__23299;
    wire N__23296;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23227;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23206;
    wire N__23203;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23011;
    wire N__23008;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22732;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22591;
    wire N__22590;
    wire N__22589;
    wire N__22588;
    wire N__22587;
    wire N__22584;
    wire N__22583;
    wire N__22580;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22562;
    wire N__22557;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22510;
    wire N__22507;
    wire N__22504;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22336;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22318;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22291;
    wire N__22288;
    wire N__22285;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22210;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22126;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22078;
    wire N__22075;
    wire N__22072;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22060;
    wire N__22057;
    wire N__22054;
    wire N__22051;
    wire N__22048;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21982;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire delay_tr_input_ibuf_gb_io_gb_input;
    wire delay_hc_input_ibuf_gb_io_gb_input;
    wire \pwm_generator_inst.O_0_1 ;
    wire \pwm_generator_inst.O_0_0 ;
    wire \pwm_generator_inst.O_0_5 ;
    wire \pwm_generator_inst.O_0_3 ;
    wire \pwm_generator_inst.O_0_4 ;
    wire \pwm_generator_inst.O_0_2 ;
    wire \pwm_generator_inst.O_0_6 ;
    wire GNDG0;
    wire VCCG0;
    wire \pwm_generator_inst.O_0 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_0 ;
    wire bfn_1_14_0_;
    wire \pwm_generator_inst.O_1 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_1 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_0 ;
    wire \pwm_generator_inst.O_2 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_2 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_1 ;
    wire \pwm_generator_inst.O_3 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_3 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_2 ;
    wire \pwm_generator_inst.O_4 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_4 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_3 ;
    wire \pwm_generator_inst.O_5 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_5 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_4 ;
    wire \pwm_generator_inst.O_6 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_6 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_5 ;
    wire \pwm_generator_inst.O_7 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_7 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_7 ;
    wire \pwm_generator_inst.O_8 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_8 ;
    wire bfn_1_15_0_;
    wire \pwm_generator_inst.O_9 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_9 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_8 ;
    wire \pwm_generator_inst.O_10 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_10 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_9 ;
    wire \pwm_generator_inst.O_11 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_11 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_10 ;
    wire \pwm_generator_inst.O_12 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_12 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_11 ;
    wire \pwm_generator_inst.O_13 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_13 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_12 ;
    wire \pwm_generator_inst.O_14 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_14 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_13 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_14 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_15 ;
    wire bfn_1_16_0_;
    wire \pwm_generator_inst.un18_threshold_1_cry_16 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_17 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_18 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_19 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_20 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_21 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_22 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_23 ;
    wire bfn_1_17_0_;
    wire \pwm_generator_inst.un18_threshold_1_cry_24 ;
    wire \pwm_generator_inst.un18_threshold_1_cry_25 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_19 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_21 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_22 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_23 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_17 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_25 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_20 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_24 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_18 ;
    wire \pwm_generator_inst.un5_threshold_2_0 ;
    wire \pwm_generator_inst.un5_threshold_1_15 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_15 ;
    wire bfn_1_19_0_;
    wire \pwm_generator_inst.un5_threshold_2_1 ;
    wire \pwm_generator_inst.un5_threshold_1_16 ;
    wire \pwm_generator_inst.un18_threshold_1_axb_16 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un5_threshold_2_2 ;
    wire \pwm_generator_inst.un5_threshold_1_17 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un5_threshold_2_3 ;
    wire \pwm_generator_inst.un5_threshold_1_18 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un5_threshold_1_19 ;
    wire \pwm_generator_inst.un5_threshold_2_4 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un5_threshold_1_20 ;
    wire \pwm_generator_inst.un5_threshold_2_5 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un5_threshold_1_21 ;
    wire \pwm_generator_inst.un5_threshold_2_6 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un5_threshold_1_22 ;
    wire \pwm_generator_inst.un5_threshold_2_7 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un5_threshold_1_23 ;
    wire \pwm_generator_inst.un5_threshold_2_8 ;
    wire bfn_1_20_0_;
    wire \pwm_generator_inst.un5_threshold_1_24 ;
    wire \pwm_generator_inst.un5_threshold_2_9 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un5_threshold_1_25 ;
    wire \pwm_generator_inst.un5_threshold_2_10 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un5_threshold_2_11 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un5_threshold_2_12 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un5_threshold_2_13 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_12 ;
    wire \pwm_generator_inst.un5_threshold_2_14 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_13 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_14 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_15 ;
    wire bfn_1_21_0_;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0 ;
    wire \pwm_generator_inst.un5_threshold_1_26 ;
    wire \pwm_generator_inst.un5_threshold_2_1_16 ;
    wire \pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_ ;
    wire \pwm_generator_inst.un5_threshold_2_1_15 ;
    wire \pwm_generator_inst.un5_threshold_add_1_axb_16 ;
    wire bfn_1_23_0_;
    wire \pwm_generator_inst.O_0_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_0 ;
    wire \pwm_generator_inst.O_0_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_1 ;
    wire \pwm_generator_inst.O_0_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_2 ;
    wire \pwm_generator_inst.O_0_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_3 ;
    wire \pwm_generator_inst.O_0_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_4 ;
    wire \pwm_generator_inst.O_0_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_5 ;
    wire \pwm_generator_inst.O_0_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_6 ;
    wire \pwm_generator_inst.un3_threshold_cry_7 ;
    wire \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0 ;
    wire bfn_1_24_0_;
    wire \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8 ;
    wire \pwm_generator_inst.un3_threshold_cry_9 ;
    wire \pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_10 ;
    wire \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_11 ;
    wire \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_13 ;
    wire \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_14 ;
    wire \pwm_generator_inst.un3_threshold_cry_15 ;
    wire \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7 ;
    wire bfn_1_25_0_;
    wire \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7 ;
    wire \pwm_generator_inst.un3_threshold_cry_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_17 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ;
    wire \pwm_generator_inst.un3_threshold_cry_18 ;
    wire \pwm_generator_inst.un2_threshold_2_12 ;
    wire \pwm_generator_inst.un3_threshold_cry_19 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ;
    wire bfn_2_17_0_;
    wire \pwm_generator_inst.un22_threshold_1_cry_0 ;
    wire \pwm_generator_inst.un18_threshold1_19 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_1 ;
    wire \pwm_generator_inst.un18_threshold1_20 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_2 ;
    wire \pwm_generator_inst.un18_threshold1_21 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_3 ;
    wire \pwm_generator_inst.un18_threshold1_22 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_4 ;
    wire \pwm_generator_inst.un18_threshold1_23 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_5 ;
    wire \pwm_generator_inst.un18_threshold1_24 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_6 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_7 ;
    wire bfn_2_18_0_;
    wire \pwm_generator_inst.un22_threshold_1_cry_8 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ;
    wire \pwm_generator_inst.un18_threshold1_25 ;
    wire \pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO ;
    wire \pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO ;
    wire \pwm_generator_inst.un18_threshold1_18 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ;
    wire \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ;
    wire \pwm_generator_inst.N_179_i ;
    wire \pwm_generator_inst.counter_i_0 ;
    wire bfn_3_17_0_;
    wire \pwm_generator_inst.N_180_i ;
    wire \pwm_generator_inst.counter_i_1 ;
    wire \pwm_generator_inst.un14_counter_cry_0 ;
    wire \pwm_generator_inst.N_181_i ;
    wire \pwm_generator_inst.counter_i_2 ;
    wire \pwm_generator_inst.un14_counter_cry_1 ;
    wire \pwm_generator_inst.N_182_i ;
    wire \pwm_generator_inst.counter_i_3 ;
    wire \pwm_generator_inst.un14_counter_cry_2 ;
    wire \pwm_generator_inst.N_183_i ;
    wire \pwm_generator_inst.counter_i_4 ;
    wire \pwm_generator_inst.un14_counter_cry_3 ;
    wire \pwm_generator_inst.N_184_i ;
    wire \pwm_generator_inst.counter_i_5 ;
    wire \pwm_generator_inst.un14_counter_cry_4 ;
    wire \pwm_generator_inst.N_185_i ;
    wire \pwm_generator_inst.counter_i_6 ;
    wire \pwm_generator_inst.un14_counter_cry_5 ;
    wire \pwm_generator_inst.N_186_i ;
    wire \pwm_generator_inst.counter_i_7 ;
    wire \pwm_generator_inst.un14_counter_cry_6 ;
    wire \pwm_generator_inst.un14_counter_cry_7 ;
    wire \pwm_generator_inst.N_187_i ;
    wire \pwm_generator_inst.counter_i_8 ;
    wire bfn_3_18_0_;
    wire \pwm_generator_inst.N_188_i ;
    wire \pwm_generator_inst.counter_i_9 ;
    wire \pwm_generator_inst.un14_counter_cry_8 ;
    wire \pwm_generator_inst.un14_counter_cry_9 ;
    wire pwm_output_c;
    wire \pwm_generator_inst.un1_counterlto2_0_cascade_ ;
    wire \pwm_generator_inst.un1_counterlto9_2 ;
    wire \pwm_generator_inst.un1_counterlt9_cascade_ ;
    wire \pwm_generator_inst.counterZ0Z_0 ;
    wire bfn_4_18_0_;
    wire \pwm_generator_inst.counterZ0Z_1 ;
    wire \pwm_generator_inst.counter_cry_0 ;
    wire \pwm_generator_inst.counterZ0Z_2 ;
    wire \pwm_generator_inst.counter_cry_1 ;
    wire \pwm_generator_inst.counterZ0Z_3 ;
    wire \pwm_generator_inst.counter_cry_2 ;
    wire \pwm_generator_inst.counterZ0Z_4 ;
    wire \pwm_generator_inst.counter_cry_3 ;
    wire \pwm_generator_inst.counterZ0Z_5 ;
    wire \pwm_generator_inst.counter_cry_4 ;
    wire \pwm_generator_inst.counterZ0Z_6 ;
    wire \pwm_generator_inst.counter_cry_5 ;
    wire \pwm_generator_inst.counterZ0Z_7 ;
    wire \pwm_generator_inst.counter_cry_6 ;
    wire \pwm_generator_inst.counter_cry_7 ;
    wire \pwm_generator_inst.counterZ0Z_8 ;
    wire bfn_4_19_0_;
    wire \pwm_generator_inst.un1_counter_0 ;
    wire \pwm_generator_inst.counter_cry_8 ;
    wire \pwm_generator_inst.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ;
    wire bfn_7_7_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_7 ;
    wire bfn_7_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_15 ;
    wire bfn_7_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_23 ;
    wire bfn_7_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counter_cry_28 ;
    wire elapsed_time_ns_1_RNI5GPBB_0_27;
    wire elapsed_time_ns_1_RNI5GPBB_0_27_cascade_;
    wire elapsed_time_ns_1_RNI7IPBB_0_29;
    wire elapsed_time_ns_1_RNI7IPBB_0_29_cascade_;
    wire elapsed_time_ns_1_RNIJI91B_0_7;
    wire elapsed_time_ns_1_RNIJI91B_0_7_cascade_;
    wire elapsed_time_ns_1_RNI1CPBB_0_23;
    wire \delay_measurement_inst.delay_tr_timer.running_i ;
    wire elapsed_time_ns_1_RNI6GOBB_0_19;
    wire elapsed_time_ns_1_RNI6GOBB_0_19_cascade_;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_0 ;
    wire bfn_7_17_0_;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_1 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_2 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_3 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_4 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_5 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_7 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_8 ;
    wire bfn_7_18_0_;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_9 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_10 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_11 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_12 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_13 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.counter_i_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ;
    wire bfn_7_19_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_30 ;
    wire bfn_7_20_0_;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt30 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_lt28 ;
    wire clk_12mhz;
    wire GB_BUFFER_clk_12mhz_THRU_CO;
    wire bfn_8_8_0_;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ;
    wire bfn_8_9_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ;
    wire bfn_8_10_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ;
    wire bfn_8_11_0_;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ;
    wire elapsed_time_ns_1_RNIT6OBB_0_10;
    wire elapsed_time_ns_1_RNI4FPBB_0_26;
    wire elapsed_time_ns_1_RNI4FPBB_0_26_cascade_;
    wire elapsed_time_ns_1_RNI2COBB_0_15;
    wire elapsed_time_ns_1_RNILK91B_0_9;
    wire elapsed_time_ns_1_RNILK91B_0_9_cascade_;
    wire elapsed_time_ns_1_RNI1BOBB_0_14;
    wire \phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ;
    wire bfn_8_13_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ;
    wire bfn_8_14_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_16;
    wire bfn_8_15_0_;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_17;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_18;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_19;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_21;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ;
    wire bfn_8_16_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.counter ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_0 ;
    wire bfn_8_17_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_0 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_2 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_1 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_2 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_4 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_3 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_5 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_4 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_5 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_7 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_6 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_7 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_8 ;
    wire bfn_8_18_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_9 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_8 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_10 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_9 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_11 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_10 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_12 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_11 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_13 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_12 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_13 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_15 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_14 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_15 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_16 ;
    wire bfn_8_19_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_17 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_16 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_18 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_17 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_19 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_18 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_20 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_19 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_21 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_20 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_22 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_21 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_22 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_23 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_24 ;
    wire bfn_8_20_0_;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_25 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_24 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_26 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_25 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_27 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_26 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_27 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_29 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_30 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_29 ;
    wire \phase_controller_inst2.stoper_tr.counter_cry_30 ;
    wire \phase_controller_inst2.stoper_tr.counterZ0Z_31 ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0_g ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_15 ;
    wire bfn_8_21_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_8 ;
    wire bfn_8_22_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ;
    wire \phase_controller_inst2.stateZ0Z_2 ;
    wire \phase_controller_inst2.hc_time_passed ;
    wire \phase_controller_inst2.start_timer_tr_0_sqmuxa ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ;
    wire elapsed_time_ns_1_RNI5FOBB_0_18;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ;
    wire elapsed_time_ns_1_RNIV8OBB_0_12;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ;
    wire elapsed_time_ns_1_RNI3DOBB_0_16;
    wire elapsed_time_ns_1_RNI3DOBB_0_16_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ;
    wire elapsed_time_ns_1_RNIHG91B_0_5;
    wire elapsed_time_ns_1_RNIHG91B_0_5_cascade_;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ;
    wire bfn_9_11_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ;
    wire bfn_9_12_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ;
    wire bfn_9_13_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ;
    wire bfn_9_14_0_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ;
    wire elapsed_time_ns_1_RNI6HPBB_0_28;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ;
    wire \pwm_generator_inst.un2_threshold_2_0 ;
    wire \pwm_generator_inst.un2_threshold_1_15 ;
    wire \pwm_generator_inst.un3_threshold_axbZ0Z_8 ;
    wire bfn_9_15_0_;
    wire \pwm_generator_inst.un2_threshold_2_1 ;
    wire \pwm_generator_inst.un2_threshold_1_16 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_0 ;
    wire \pwm_generator_inst.un2_threshold_1_17 ;
    wire \pwm_generator_inst.un2_threshold_2_2 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_1 ;
    wire \pwm_generator_inst.un2_threshold_1_18 ;
    wire \pwm_generator_inst.un2_threshold_2_3 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_2 ;
    wire \pwm_generator_inst.un2_threshold_2_4 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_3 ;
    wire \pwm_generator_inst.un2_threshold_2_5 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_4 ;
    wire \pwm_generator_inst.un2_threshold_2_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_5 ;
    wire \pwm_generator_inst.un2_threshold_2_7 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_6 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_7 ;
    wire \pwm_generator_inst.un2_threshold_2_8 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ;
    wire bfn_9_16_0_;
    wire \pwm_generator_inst.un2_threshold_2_9 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_8 ;
    wire \pwm_generator_inst.un2_threshold_2_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_9 ;
    wire \pwm_generator_inst.un2_threshold_1_19 ;
    wire \pwm_generator_inst.un2_threshold_2_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_10 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11 ;
    wire \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_24;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_25;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_26;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_27;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator ;
    wire bfn_9_18_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_2 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_3 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_2 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_4 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_5 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_6 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_8 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_7 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_8 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_9 ;
    wire bfn_9_19_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_10 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_9 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_11 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_10 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_12 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_13 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_12 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_14 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_16 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_15 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_17 ;
    wire bfn_9_20_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_18 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_19 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_20 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_21 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_22 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_24 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_23 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_25 ;
    wire bfn_9_21_0_;
    wire \current_shift_inst.PI_CTRL.integrator_1_26 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_27 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_28 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_29 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_30 ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ;
    wire \current_shift_inst.PI_CTRL.un1_integrator_cry_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ;
    wire s3_phy_c;
    wire s4_phy_c;
    wire \phase_controller_inst2.stoper_hc.runningZ0 ;
    wire il_min_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_1 ;
    wire il_max_comp2_c;
    wire \phase_controller_inst2.stateZ0Z_0 ;
    wire \phase_controller_inst2.state_ns_0_0_1_cascade_ ;
    wire \phase_controller_inst2.stateZ0Z_3 ;
    wire \phase_controller_inst2.stoper_tr.un4_start_0_cascade_ ;
    wire \phase_controller_inst2.tr_time_passed ;
    wire \phase_controller_inst2.stoper_tr.un2_start_0 ;
    wire \phase_controller_inst2.start_timer_trZ0 ;
    wire \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_tr.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ;
    wire elapsed_time_ns_1_RNIDC91B_0_1;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ;
    wire elapsed_time_ns_1_RNI4EOBB_0_17;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ;
    wire elapsed_time_ns_1_RNIU7OBB_0_11;
    wire elapsed_time_ns_1_RNIU7OBB_0_11_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ;
    wire \delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ;
    wire elapsed_time_ns_1_RNIED91B_0_2;
    wire elapsed_time_ns_1_RNIFE91B_0_3;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ;
    wire elapsed_time_ns_1_RNIIH91B_0_6;
    wire elapsed_time_ns_1_RNIIH91B_0_6_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ;
    wire elapsed_time_ns_1_RNIGF91B_0_4;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ;
    wire elapsed_time_ns_1_RNI2DPBB_0_24;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ;
    wire elapsed_time_ns_1_RNIKJ91B_0_8;
    wire elapsed_time_ns_1_RNIKJ91B_0_8_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ;
    wire elapsed_time_ns_1_RNI0BPBB_0_22;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ;
    wire elapsed_time_ns_1_RNIU8PBB_0_20;
    wire elapsed_time_ns_1_RNIU8PBB_0_20_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ;
    wire elapsed_time_ns_1_RNI3EPBB_0_25;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_1;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_6;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_5;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_13;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_7;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_4;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_2;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_3;
    wire \phase_controller_inst1.stoper_tr.counter_i_0 ;
    wire bfn_10_14_0_;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_1 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_2 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_3 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_4 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_5 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_7 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_8 ;
    wire bfn_10_15_0_;
    wire \phase_controller_inst1.stoper_tr.counter_i_9 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_11 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_12 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_13 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_i_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt16 ;
    wire bfn_10_16_0_;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_30 ;
    wire bfn_10_17_0_;
    wire \phase_controller_inst1.stoper_tr.un2_start_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ;
    wire \current_shift_inst.PI_CTRL.N_44_cascade_ ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_2_15 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_1_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_0 ;
    wire bfn_11_5_0_;
    wire \phase_controller_inst2.stoper_hc.counter_i_1 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_2 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_3 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_4 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_5 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_7 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_8 ;
    wire bfn_11_6_0_;
    wire \phase_controller_inst2.stoper_hc.counter_i_9 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_11 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_12 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_13 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.counter_i_15 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_15 ;
    wire bfn_11_7_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_30 ;
    wire bfn_11_8_0_;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt20 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ;
    wire \phase_controller_inst2.stoper_hc.counter ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_0 ;
    wire bfn_11_9_0_;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_0 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_1 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_2 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_3 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_4 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_5 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_6 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_7 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_8 ;
    wire bfn_11_10_0_;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_8 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_9 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_10 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_11 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_12 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_13 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_14 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_15 ;
    wire bfn_11_11_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_16 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_17 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_18 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_19 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_20 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_21 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_23 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_22 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_23 ;
    wire bfn_11_12_0_;
    wire \phase_controller_inst2.stoper_hc.counter_cry_24 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_25 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_26 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_27 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_28 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_29 ;
    wire \phase_controller_inst2.stoper_hc.start_latched_i_0 ;
    wire \phase_controller_inst2.stoper_hc.counter_cry_30 ;
    wire \phase_controller_inst2.stoper_hc.un2_start_0 ;
    wire \phase_controller_inst1.stoper_tr.counter ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_0 ;
    wire bfn_11_13_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_1 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_0 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_2 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_1 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_3 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_2 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_4 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_3 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_5 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_4 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_5 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_7 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_6 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_7 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_8 ;
    wire bfn_11_14_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_9 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_11 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_10 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_12 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_11 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_13 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_12 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_14 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_13 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_15 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_14 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_15 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_16 ;
    wire bfn_11_15_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_17 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_16 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_18 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_17 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_19 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_18 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_19 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_20 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_21 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_22 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_23 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_24 ;
    wire bfn_11_16_0_;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_25 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_24 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_26 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_25 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_27 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_26 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_27 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_29 ;
    wire \phase_controller_inst1.stoper_tr.start_latched_i_0 ;
    wire \phase_controller_inst1.stoper_tr.counter_cry_30 ;
    wire \phase_controller_inst1.stoper_tr.un2_start_0_g ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt20 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_20;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_21 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt22 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_22;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_23 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_22 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_23;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ;
    wire \phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ;
    wire \phase_controller_inst2.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_tr.start_latched_i_0 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_47 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_77 ;
    wire \current_shift_inst.PI_CTRL.N_43 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ;
    wire \current_shift_inst.PI_CTRL.N_46_16 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0 ;
    wire \current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_46_21 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ;
    wire \current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt16 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_16 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_18 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt24 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt26 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_26 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt28 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_29 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_31 ;
    wire \phase_controller_inst2.stoper_hc.counterZ0Z_30 ;
    wire \phase_controller_inst2.stoper_hc.un6_running_lt30 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ;
    wire elapsed_time_ns_1_RNI0AOBB_0_13;
    wire elapsed_time_ns_1_RNI0AOBB_0_13_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ;
    wire elapsed_time_ns_1_RNIV9PBB_0_21;
    wire \delay_measurement_inst.delay_tr_timer.delay_tr3 ;
    wire \delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ;
    wire elapsed_time_ns_1_RNIVAQBB_0_30;
    wire elapsed_time_ns_1_RNIVAQBB_0_30_cascade_;
    wire \phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ;
    wire \phase_controller_inst2.start_flagZ0 ;
    wire \phase_controller_inst2.stateZ0Z_4 ;
    wire start_stop_c;
    wire \phase_controller_inst1.stateZ0Z_4 ;
    wire \phase_controller_inst1.state_ns_0_0_1_cascade_ ;
    wire \phase_controller_inst1.start_flagZ0 ;
    wire \phase_controller_inst1.stoper_tr.un4_start_0_cascade_ ;
    wire \phase_controller_inst1.tr_time_passed ;
    wire \phase_controller_inst1.stateZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_tr.runningZ0 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_14;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_12;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_15;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_11;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_8;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_9;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_10;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt28 ;
    wire phase_controller_inst1_stoper_tr_target_ticks_1_i_28;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_29 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_30 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ;
    wire \phase_controller_inst1.stoper_tr.counterZ0Z_31 ;
    wire \phase_controller_inst1.stoper_tr.un6_running_lt30 ;
    wire \phase_controller_inst2.start_timer_hcZ0 ;
    wire \phase_controller_inst2.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst2.stoper_hc.un4_start_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_1 ;
    wire bfn_12_20_0_;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_2 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_3 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_4 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_5 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_6 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_9 ;
    wire bfn_12_21_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_17 ;
    wire bfn_12_22_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_25 ;
    wire bfn_12_23_0_;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ;
    wire GB_BUFFER_reset_c_g_THRU_CO;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ;
    wire bfn_13_7_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_7 ;
    wire bfn_13_8_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_15 ;
    wire bfn_13_9_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_19 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_23 ;
    wire bfn_13_10_0_;
    wire \phase_controller_inst1.stoper_hc.counter_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.counter_cry_30 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_31 ;
    wire elapsed_time_ns_1_RNI36DN9_0_25;
    wire elapsed_time_ns_1_RNI36DN9_0_25_cascade_;
    wire elapsed_time_ns_1_RNIV2EN9_0_30;
    wire elapsed_time_ns_1_RNI03DN9_0_22;
    wire elapsed_time_ns_1_RNI03DN9_0_22_cascade_;
    wire elapsed_time_ns_1_RNI7ADN9_0_29;
    wire elapsed_time_ns_1_RNI7ADN9_0_29_cascade_;
    wire \phase_controller_inst1.start_timer_tr_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un2_start_0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_168_i ;
    wire \delay_measurement_inst.delay_tr_timer.runningZ0 ;
    wire \delay_measurement_inst.delay_tr_timer.N_167_i ;
    wire il_max_comp1_c;
    wire \phase_controller_inst1.stoper_hc.runningZ0 ;
    wire \phase_controller_inst1.stoper_hc.un4_start_0_cascade_ ;
    wire \phase_controller_inst1.start_timer_hcZ0 ;
    wire il_min_comp1_c;
    wire \phase_controller_inst1.stateZ0Z_2 ;
    wire \phase_controller_inst1.hc_time_passed ;
    wire \phase_controller_inst1.stoper_hc.start_latched_i_0 ;
    wire \phase_controller_inst1.stoper_tr.start_latchedZ0 ;
    wire \phase_controller_inst1.start_timer_trZ0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ;
    wire elapsed_time_ns_1_RNI0CQBB_0_31;
    wire \phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ;
    wire \phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axb_0 ;
    wire bfn_13_17_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_1 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_2 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_3 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_4 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_5 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_6 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_7 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_8 ;
    wire bfn_13_18_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_8 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_9 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_10 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_11 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_12 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_14 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_15 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_16 ;
    wire bfn_13_19_0_;
    wire \current_shift_inst.PI_CTRL.prop_term_1_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_17 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_22 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_23 ;
    wire bfn_13_20_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_28 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_29 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_cry_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.integratorZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_18 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_24 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_22 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_23 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_23 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_20 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_21 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_30 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_29 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_27 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_26 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_31 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_31 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_25 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_25 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_28 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_28 ;
    wire \delay_measurement_inst.stop_timer_trZ0 ;
    wire \delay_measurement_inst.start_timer_trZ0 ;
    wire delay_tr_input_c_g;
    wire \phase_controller_inst1.stateZ0Z_1 ;
    wire s2_phy_c;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_0 ;
    wire bfn_14_5_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_1 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_0 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_2 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_3 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_4 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_5 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_7 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_8 ;
    wire bfn_14_6_0_;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_9 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_10 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_11 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_12 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_13 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.counter_i_15 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_15 ;
    wire bfn_14_7_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt30 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30 ;
    wire bfn_14_8_0_;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt16 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_17 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_16 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ;
    wire elapsed_time_ns_1_RNIG23T9_0_4;
    wire elapsed_time_ns_1_RNIG23T9_0_4_cascade_;
    wire \phase_controller_inst1.stoper_hc.start_latchedZ0 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ;
    wire \phase_controller_inst1.stoper_hc.counter ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt20 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt22 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt24 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_lt26 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_27 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.counterZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ;
    wire bfn_14_11_0_;
    wire \current_shift_inst.timer_s1.counter_cry_0 ;
    wire \current_shift_inst.timer_s1.counter_cry_1 ;
    wire \current_shift_inst.timer_s1.counter_cry_2 ;
    wire \current_shift_inst.timer_s1.counter_cry_3 ;
    wire \current_shift_inst.timer_s1.counter_cry_4 ;
    wire \current_shift_inst.timer_s1.counter_cry_5 ;
    wire \current_shift_inst.timer_s1.counter_cry_6 ;
    wire \current_shift_inst.timer_s1.counter_cry_7 ;
    wire bfn_14_12_0_;
    wire \current_shift_inst.timer_s1.counter_cry_8 ;
    wire \current_shift_inst.timer_s1.counter_cry_9 ;
    wire \current_shift_inst.timer_s1.counter_cry_10 ;
    wire \current_shift_inst.timer_s1.counter_cry_11 ;
    wire \current_shift_inst.timer_s1.counter_cry_12 ;
    wire \current_shift_inst.timer_s1.counter_cry_13 ;
    wire \current_shift_inst.timer_s1.counter_cry_14 ;
    wire \current_shift_inst.timer_s1.counter_cry_15 ;
    wire bfn_14_13_0_;
    wire \current_shift_inst.timer_s1.counter_cry_16 ;
    wire \current_shift_inst.timer_s1.counter_cry_17 ;
    wire \current_shift_inst.timer_s1.counter_cry_18 ;
    wire \current_shift_inst.timer_s1.counter_cry_19 ;
    wire \current_shift_inst.timer_s1.counter_cry_20 ;
    wire \current_shift_inst.timer_s1.counter_cry_21 ;
    wire \current_shift_inst.timer_s1.counter_cry_22 ;
    wire \current_shift_inst.timer_s1.counter_cry_23 ;
    wire bfn_14_14_0_;
    wire \current_shift_inst.timer_s1.counter_cry_24 ;
    wire \current_shift_inst.timer_s1.counter_cry_25 ;
    wire \current_shift_inst.timer_s1.counter_cry_26 ;
    wire \current_shift_inst.timer_s1.counter_cry_27 ;
    wire \current_shift_inst.timer_s1.counter_cry_28 ;
    wire bfn_14_15_0_;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_2 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_3 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_4 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_5 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_6 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_7 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_8 ;
    wire bfn_14_16_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_9 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_11 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_12 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_13 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_14 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_15 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_16 ;
    wire bfn_14_17_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_17 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_18 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_19 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_20 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_21 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_22 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_23 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_24 ;
    wire bfn_14_18_0_;
    wire \current_shift_inst.timer_s1.counterZ0Z_25 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_28 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_26 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_29 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_27 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_fast_31 ;
    wire \current_shift_inst.control_input_1 ;
    wire bfn_14_19_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ;
    wire \current_shift_inst.control_input_cry_0 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ;
    wire \current_shift_inst.control_input_cry_1 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ;
    wire \current_shift_inst.control_input_cry_2 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ;
    wire \current_shift_inst.control_input_cry_3 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ;
    wire \current_shift_inst.control_input_cry_4 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ;
    wire \current_shift_inst.control_input_cry_5 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ;
    wire \current_shift_inst.control_input_cry_6 ;
    wire \current_shift_inst.control_input_cry_7 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ;
    wire bfn_14_20_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ;
    wire \current_shift_inst.control_input_cry_8 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ;
    wire \current_shift_inst.control_input_cry_9 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ;
    wire \current_shift_inst.control_input_cry_10 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ;
    wire \current_shift_inst.control_input_cry_11 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ;
    wire \current_shift_inst.control_input_cry_12 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ;
    wire \current_shift_inst.control_input_cry_13 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ;
    wire \current_shift_inst.control_input_cry_14 ;
    wire \current_shift_inst.control_input_cry_15 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ;
    wire bfn_14_21_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ;
    wire \current_shift_inst.control_input_cry_16 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ;
    wire \current_shift_inst.control_input_cry_17 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ;
    wire \current_shift_inst.control_input_cry_18 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ;
    wire \current_shift_inst.control_input_cry_19 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ;
    wire \current_shift_inst.control_input_cry_20 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ;
    wire \current_shift_inst.control_input_cry_21 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ;
    wire \current_shift_inst.control_input_cry_22 ;
    wire \current_shift_inst.control_input_cry_23 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ;
    wire bfn_14_22_0_;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ;
    wire \current_shift_inst.control_input_cry_24 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ;
    wire \current_shift_inst.control_input_cry_25 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ;
    wire \current_shift_inst.control_input_cry_26 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ;
    wire \current_shift_inst.control_input_cry_27 ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ;
    wire \current_shift_inst.control_input_cry_28 ;
    wire \current_shift_inst.control_input_cry_29 ;
    wire \current_shift_inst.control_input_31 ;
    wire \current_shift_inst.control_input_31_cascade_ ;
    wire \current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ;
    wire delay_hc_input_c_g;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ;
    wire \phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ;
    wire bfn_15_7_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_1;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_2;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_3;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_4;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_5;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_6;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_7;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_8;
    wire bfn_15_8_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_9;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_10;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_11;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_12;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_13;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_14;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_16;
    wire bfn_15_9_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_17;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_18;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_19;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_20;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_21;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_22;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_23;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_24;
    wire bfn_15_10_0_;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_25;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_26;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_27;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ;
    wire elapsed_time_ns_1_RNIF13T9_0_3;
    wire \current_shift_inst.timer_s1.counterZ0Z_1 ;
    wire bfn_15_16_0_;
    wire \current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_0 ;
    wire \current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_1 ;
    wire \current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_2 ;
    wire \current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_3 ;
    wire \current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_4 ;
    wire \current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_5 ;
    wire \current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_6 ;
    wire \current_shift_inst.un10_control_input_cry_7 ;
    wire \current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ;
    wire bfn_15_17_0_;
    wire \current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_8 ;
    wire \current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_9 ;
    wire \current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_10 ;
    wire \current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_11 ;
    wire \current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_12 ;
    wire \current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_13 ;
    wire \current_shift_inst.un10_control_input_cry_14 ;
    wire \current_shift_inst.un10_control_input_cry_15 ;
    wire bfn_15_18_0_;
    wire \current_shift_inst.un10_control_input_cry_16 ;
    wire \current_shift_inst.un10_control_input_cry_17 ;
    wire \current_shift_inst.un10_control_input_cry_18 ;
    wire \current_shift_inst.un10_control_input_cry_19 ;
    wire \current_shift_inst.un10_control_input_cry_20 ;
    wire \current_shift_inst.un10_control_input_cry_21 ;
    wire \current_shift_inst.un10_control_input_cry_22 ;
    wire \current_shift_inst.un10_control_input_cry_23 ;
    wire bfn_15_19_0_;
    wire \current_shift_inst.un10_control_input_cry_24 ;
    wire \current_shift_inst.un10_control_input_cry_25 ;
    wire \current_shift_inst.un10_control_input_cry_26 ;
    wire \current_shift_inst.un10_control_input_cry_27 ;
    wire \current_shift_inst.un10_control_input_cry_28 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29 ;
    wire \current_shift_inst.un10_control_input_cry_30 ;
    wire \current_shift_inst.control_input_axb_1 ;
    wire \current_shift_inst.control_input_axb_2 ;
    wire \current_shift_inst.control_input_axb_3 ;
    wire \current_shift_inst.control_input_axb_4 ;
    wire \current_shift_inst.control_input_axb_5 ;
    wire \current_shift_inst.control_input_axb_6 ;
    wire \current_shift_inst.control_input_axb_7 ;
    wire \current_shift_inst.control_input_axb_13 ;
    wire \current_shift_inst.control_input_axb_21 ;
    wire \current_shift_inst.control_input_axb_26 ;
    wire \current_shift_inst.control_input_axb_22 ;
    wire \current_shift_inst.control_input_axb_17 ;
    wire \current_shift_inst.control_input_axb_16 ;
    wire \current_shift_inst.control_input_axb_25 ;
    wire \current_shift_inst.control_input_axb_27 ;
    wire \current_shift_inst.control_input_axb_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ;
    wire \current_shift_inst.control_input_axb_18 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_15;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ;
    wire elapsed_time_ns_1_RNI04EN9_0_31_cascade_;
    wire \phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ;
    wire \phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ;
    wire bfn_16_8_0_;
    wire elapsed_time_ns_1_RNIE03T9_0_2;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ;
    wire \phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ;
    wire bfn_16_9_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ;
    wire bfn_16_10_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ;
    wire bfn_16_11_0_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ;
    wire \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ;
    wire elapsed_time_ns_1_RNI04EN9_0_31;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ;
    wire phase_controller_inst1_stoper_hc_target_ticks_1_i_28;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ;
    wire \current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ;
    wire \current_shift_inst.timer_s1.counterZ0Z_0 ;
    wire \current_shift_inst.un4_control_input_1_axb_1 ;
    wire bfn_16_13_0_;
    wire \current_shift_inst.un4_control_input_1_axb_2 ;
    wire \current_shift_inst.un4_control_input_1_cry_1 ;
    wire \current_shift_inst.un4_control_input_1_axb_3 ;
    wire \current_shift_inst.un4_control_input_1_cry_2 ;
    wire \current_shift_inst.un4_control_input_1_axb_4 ;
    wire \current_shift_inst.un4_control_input_1_cry_3 ;
    wire \current_shift_inst.un4_control_input_1_axb_5 ;
    wire \current_shift_inst.un4_control_input_1_cry_4 ;
    wire \current_shift_inst.un4_control_input_1_axb_6 ;
    wire \current_shift_inst.un4_control_input_1_cry_5 ;
    wire \current_shift_inst.un4_control_input_1_axb_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_6 ;
    wire \current_shift_inst.un4_control_input_1_axb_8 ;
    wire \current_shift_inst.un4_control_input_1_cry_7 ;
    wire \current_shift_inst.un4_control_input_1_cry_8 ;
    wire \current_shift_inst.un4_control_input_1_axb_9 ;
    wire bfn_16_14_0_;
    wire \current_shift_inst.un4_control_input_1_axb_10 ;
    wire \current_shift_inst.un4_control_input_1_cry_9 ;
    wire \current_shift_inst.un4_control_input_1_axb_11 ;
    wire \current_shift_inst.un4_control_input_1_cry_10 ;
    wire \current_shift_inst.un4_control_input_1_axb_12 ;
    wire \current_shift_inst.un4_control_input_1_cry_11 ;
    wire \current_shift_inst.un4_control_input_1_axb_13 ;
    wire \current_shift_inst.un4_control_input_1_cry_12 ;
    wire \current_shift_inst.un4_control_input_1_axb_14 ;
    wire \current_shift_inst.un4_control_input_1_cry_13 ;
    wire \current_shift_inst.un4_control_input_1_axb_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_14 ;
    wire \current_shift_inst.un4_control_input_1_axb_16 ;
    wire \current_shift_inst.un4_control_input_1_cry_15 ;
    wire \current_shift_inst.un4_control_input_1_cry_16 ;
    wire \current_shift_inst.un4_control_input_1_axb_17 ;
    wire bfn_16_15_0_;
    wire \current_shift_inst.un4_control_input_1_cry_17 ;
    wire \current_shift_inst.un4_control_input_1_axb_19 ;
    wire \current_shift_inst.un4_control_input_1_cry_18 ;
    wire \current_shift_inst.un4_control_input_1_axb_20 ;
    wire \current_shift_inst.un4_control_input_1_cry_19 ;
    wire \current_shift_inst.un4_control_input_1_axb_21 ;
    wire \current_shift_inst.un4_control_input_1_cry_20 ;
    wire \current_shift_inst.un4_control_input_1_axb_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_21 ;
    wire \current_shift_inst.un4_control_input_1_axb_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_22 ;
    wire \current_shift_inst.un4_control_input_1_cry_23 ;
    wire \current_shift_inst.un4_control_input_1_cry_24 ;
    wire bfn_16_16_0_;
    wire \current_shift_inst.un4_control_input_1_cry_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_26 ;
    wire \current_shift_inst.un4_control_input_1_axb_28 ;
    wire \current_shift_inst.un4_control_input_1_cry_27 ;
    wire \current_shift_inst.un4_control_input_1_cry_28 ;
    wire \current_shift_inst.un4_control_input1_31 ;
    wire \current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_25 ;
    wire \current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ;
    wire \current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ;
    wire \current_shift_inst.un4_control_input_1_axb_29 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31_rep1 ;
    wire \current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ;
    wire \current_shift_inst.control_input_axb_9 ;
    wire \current_shift_inst.control_input_axb_0 ;
    wire \current_shift_inst.control_input_axb_0_cascade_ ;
    wire \current_shift_inst.N_1379_i ;
    wire \current_shift_inst.control_input_axb_10 ;
    wire \current_shift_inst.control_input_axb_11 ;
    wire \current_shift_inst.control_input_axb_8 ;
    wire \current_shift_inst.control_input_axb_14 ;
    wire \current_shift_inst.control_input_axb_15 ;
    wire \current_shift_inst.control_input_axb_12 ;
    wire \current_shift_inst.control_input_axb_24 ;
    wire \current_shift_inst.control_input_axb_19 ;
    wire \current_shift_inst.elapsed_time_ns_s1_30 ;
    wire \current_shift_inst.un4_control_input1_30 ;
    wire \current_shift_inst.un4_control_input_1_axb_26 ;
    wire \current_shift_inst.control_input_axb_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_29 ;
    wire \current_shift_inst.un4_control_input1_29 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ;
    wire \current_shift_inst.un4_control_input1_25 ;
    wire elapsed_time_ns_1_RNIJ53T9_0_7;
    wire elapsed_time_ns_1_RNIJ53T9_0_7_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ;
    wire elapsed_time_ns_1_RNI25DN9_0_24;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ;
    wire elapsed_time_ns_1_RNIU0DN9_0_20;
    wire elapsed_time_ns_1_RNIU0DN9_0_20_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ;
    wire elapsed_time_ns_1_RNIH33T9_0_5;
    wire elapsed_time_ns_1_RNIH33T9_0_5_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ;
    wire elapsed_time_ns_1_RNITUBN9_0_10;
    wire elapsed_time_ns_1_RNITUBN9_0_10_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ;
    wire elapsed_time_ns_1_RNIK63T9_0_8;
    wire elapsed_time_ns_1_RNIK63T9_0_8_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ;
    wire elapsed_time_ns_1_RNI35CN9_0_16;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ;
    wire elapsed_time_ns_1_RNIL73T9_0_9;
    wire elapsed_time_ns_1_RNIL73T9_0_9_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ;
    wire elapsed_time_ns_1_RNII43T9_0_6;
    wire elapsed_time_ns_1_RNII43T9_0_6_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ;
    wire elapsed_time_ns_1_RNIUVBN9_0_11;
    wire elapsed_time_ns_1_RNIUVBN9_0_11_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ;
    wire elapsed_time_ns_1_RNI24CN9_0_15;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ;
    wire elapsed_time_ns_1_RNIV0CN9_0_12;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ;
    wire bfn_17_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ;
    wire bfn_17_11_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ;
    wire bfn_17_12_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ;
    wire bfn_17_13_0_;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ;
    wire \delay_measurement_inst.delay_hc_timer.N_165_i ;
    wire \current_shift_inst.un4_control_input_1_axb_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_10 ;
    wire \current_shift_inst.un4_control_input1_10 ;
    wire \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ;
    wire \current_shift_inst.timer_s1.N_163_i_g ;
    wire \current_shift_inst.un4_control_input1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_3 ;
    wire \current_shift_inst.elapsed_time_ns_s1_i_1 ;
    wire \current_shift_inst.un4_control_input1_1 ;
    wire \current_shift_inst.un4_control_input1_1_cascade_ ;
    wire \current_shift_inst.elapsed_time_ns_s1_1 ;
    wire \current_shift_inst.elapsed_time_ns_s1_13 ;
    wire \current_shift_inst.un4_control_input1_13 ;
    wire \current_shift_inst.elapsed_time_ns_s1_22 ;
    wire \current_shift_inst.un4_control_input1_22 ;
    wire \current_shift_inst.elapsed_time_ns_s1_5 ;
    wire \current_shift_inst.un4_control_input1_5 ;
    wire \current_shift_inst.elapsed_time_ns_s1_16 ;
    wire \current_shift_inst.un4_control_input1_16 ;
    wire \current_shift_inst.elapsed_time_ns_s1_28 ;
    wire \current_shift_inst.un4_control_input1_28 ;
    wire \current_shift_inst.elapsed_time_ns_s1_27 ;
    wire \current_shift_inst.un4_control_input1_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_26 ;
    wire \current_shift_inst.un4_control_input1_26 ;
    wire \current_shift_inst.un4_control_input1_31_THRU_CO ;
    wire \current_shift_inst.elapsed_time_ns_s1_21 ;
    wire \current_shift_inst.un4_control_input1_21 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0_sf ;
    wire bfn_17_18_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ;
    wire \current_shift_inst.un38_control_input_cry_0_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ;
    wire \current_shift_inst.un38_control_input_cry_1_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ;
    wire \current_shift_inst.un38_control_input_0_s0_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ;
    wire \current_shift_inst.un38_control_input_0_s0_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ;
    wire \current_shift_inst.un38_control_input_0_s0_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s0 ;
    wire \current_shift_inst.un38_control_input_0_s0_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s0 ;
    wire \current_shift_inst.un38_control_input_cry_7_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ;
    wire \current_shift_inst.un38_control_input_0_s0_8 ;
    wire bfn_17_19_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ;
    wire \current_shift_inst.un38_control_input_0_s0_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ;
    wire \current_shift_inst.un38_control_input_0_s0_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ;
    wire \current_shift_inst.un38_control_input_0_s0_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ;
    wire \current_shift_inst.un38_control_input_0_s0_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ;
    wire \current_shift_inst.un38_control_input_0_s0_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ;
    wire \current_shift_inst.un38_control_input_0_s0_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ;
    wire \current_shift_inst.un38_control_input_0_s0_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s0 ;
    wire \current_shift_inst.un38_control_input_cry_15_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ;
    wire \current_shift_inst.un38_control_input_0_s0_16 ;
    wire bfn_17_20_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ;
    wire \current_shift_inst.un38_control_input_0_s0_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ;
    wire \current_shift_inst.un38_control_input_0_s0_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ;
    wire \current_shift_inst.un38_control_input_0_s0_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ;
    wire \current_shift_inst.un38_control_input_0_s0_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ;
    wire \current_shift_inst.un38_control_input_0_s0_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ;
    wire \current_shift_inst.un38_control_input_0_s0_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ;
    wire \current_shift_inst.un38_control_input_0_s0_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s0 ;
    wire \current_shift_inst.un38_control_input_cry_23_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ;
    wire \current_shift_inst.un38_control_input_0_s0_24 ;
    wire bfn_17_21_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ;
    wire \current_shift_inst.un38_control_input_0_s0_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ;
    wire \current_shift_inst.un38_control_input_0_s0_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ;
    wire \current_shift_inst.un38_control_input_0_s0_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s0 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ;
    wire \current_shift_inst.un38_control_input_0_s0_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s0 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ;
    wire \current_shift_inst.un38_control_input_0_s0_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s0 ;
    wire \current_shift_inst.un38_control_input_axb_31_s0 ;
    wire \current_shift_inst.un38_control_input_cry_30_s0 ;
    wire \current_shift_inst.control_input_axb_28 ;
    wire elapsed_time_ns_1_RNI58DN9_0_27;
    wire elapsed_time_ns_1_RNI58DN9_0_27_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ;
    wire elapsed_time_ns_1_RNI46CN9_0_17;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ;
    wire bfn_18_7_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_0 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_1 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_2 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_3 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_4 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_5 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_6 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_7 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ;
    wire bfn_18_8_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_8 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_9 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_10 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_11 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_12 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_13 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_14 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_15 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ;
    wire bfn_18_9_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_16 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_17 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_18 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_19 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_20 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_21 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_22 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_23 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ;
    wire bfn_18_10_0_;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_24 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_25 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_26 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_27 ;
    wire \delay_measurement_inst.delay_hc_timer.counter_cry_28 ;
    wire \delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ;
    wire elapsed_time_ns_1_RNI69DN9_0_28;
    wire elapsed_time_ns_1_RNI69DN9_0_28_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ;
    wire elapsed_time_ns_1_RNIDV2T9_0_1;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ;
    wire elapsed_time_ns_1_RNI57CN9_0_18;
    wire elapsed_time_ns_1_RNI57CN9_0_18_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ;
    wire \delay_measurement_inst.delay_hc_timer.running_i ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ;
    wire \current_shift_inst.elapsed_time_ns_s1_25 ;
    wire \current_shift_inst.un4_control_input_1_axb_24 ;
    wire \current_shift_inst.elapsed_time_ns_s1_7 ;
    wire \current_shift_inst.un4_control_input1_7 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ;
    wire elapsed_time_ns_1_RNI68CN9_0_19;
    wire elapsed_time_ns_1_RNI68CN9_0_19_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ;
    wire elapsed_time_ns_1_RNIV1DN9_0_21;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ;
    wire \delay_measurement_inst.start_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.runningZ0 ;
    wire \delay_measurement_inst.stop_timer_hcZ0 ;
    wire \delay_measurement_inst.delay_hc_timer.N_166_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_17 ;
    wire \current_shift_inst.un4_control_input1_17 ;
    wire \current_shift_inst.timer_s1.N_164_i ;
    wire \current_shift_inst.un4_control_input1_12 ;
    wire \current_shift_inst.elapsed_time_ns_s1_12 ;
    wire \current_shift_inst.timer_s1.running_i ;
    wire \current_shift_inst.un4_control_input1_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_15 ;
    wire \current_shift_inst.elapsed_time_ns_s1_11 ;
    wire \current_shift_inst.un4_control_input1_11 ;
    wire \current_shift_inst.timer_s1.N_163_i ;
    wire \current_shift_inst.elapsed_time_ns_s1_9 ;
    wire \current_shift_inst.un4_control_input1_9 ;
    wire \current_shift_inst.elapsed_time_ns_s1_23 ;
    wire \current_shift_inst.un4_control_input1_23 ;
    wire \current_shift_inst.elapsed_time_ns_s1_24 ;
    wire \current_shift_inst.un4_control_input1_24 ;
    wire \current_shift_inst.un4_control_input1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_18 ;
    wire \current_shift_inst.elapsed_time_ns_s1_19 ;
    wire \current_shift_inst.un4_control_input1_19 ;
    wire \current_shift_inst.un4_control_input1_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_20 ;
    wire \current_shift_inst.elapsed_time_ns_s1_14 ;
    wire \current_shift_inst.un4_control_input1_14 ;
    wire \current_shift_inst.un4_control_input1_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_6 ;
    wire \current_shift_inst.elapsed_time_ns_s1_4 ;
    wire \current_shift_inst.un4_control_input1_4 ;
    wire \current_shift_inst.un4_control_input1_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_2 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ;
    wire \current_shift_inst.un4_control_input1_8 ;
    wire \current_shift_inst.elapsed_time_ns_s1_8 ;
    wire bfn_18_17_0_;
    wire \current_shift_inst.un38_control_input_5_1 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_0_s1 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ;
    wire \current_shift_inst.un38_control_input_cry_1_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ;
    wire \current_shift_inst.un38_control_input_0_s1_3 ;
    wire \current_shift_inst.un38_control_input_cry_2_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ;
    wire \current_shift_inst.un38_control_input_0_s1_4 ;
    wire \current_shift_inst.un38_control_input_cry_3_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ;
    wire \current_shift_inst.un38_control_input_0_s1_5 ;
    wire \current_shift_inst.un38_control_input_cry_4_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ;
    wire \current_shift_inst.un38_control_input_0_s1_6 ;
    wire \current_shift_inst.un38_control_input_cry_5_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ;
    wire \current_shift_inst.un38_control_input_0_s1_7 ;
    wire \current_shift_inst.un38_control_input_cry_6_s1 ;
    wire \current_shift_inst.un38_control_input_cry_7_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ;
    wire \current_shift_inst.un38_control_input_0_s1_8 ;
    wire bfn_18_18_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ;
    wire \current_shift_inst.un38_control_input_0_s1_9 ;
    wire \current_shift_inst.un38_control_input_cry_8_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ;
    wire \current_shift_inst.un38_control_input_0_s1_10 ;
    wire \current_shift_inst.un38_control_input_cry_9_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ;
    wire \current_shift_inst.un38_control_input_0_s1_11 ;
    wire \current_shift_inst.un38_control_input_cry_10_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ;
    wire \current_shift_inst.un38_control_input_0_s1_12 ;
    wire \current_shift_inst.un38_control_input_cry_11_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ;
    wire \current_shift_inst.un38_control_input_0_s1_13 ;
    wire \current_shift_inst.un38_control_input_cry_12_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ;
    wire \current_shift_inst.un38_control_input_0_s1_14 ;
    wire \current_shift_inst.un38_control_input_cry_13_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ;
    wire \current_shift_inst.un38_control_input_0_s1_15 ;
    wire \current_shift_inst.un38_control_input_cry_14_s1 ;
    wire \current_shift_inst.un38_control_input_cry_15_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNISST11_17 ;
    wire \current_shift_inst.un38_control_input_0_s1_16 ;
    wire bfn_18_19_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ;
    wire \current_shift_inst.un38_control_input_0_s1_17 ;
    wire \current_shift_inst.un38_control_input_cry_16_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI25021_19 ;
    wire \current_shift_inst.un38_control_input_0_s1_18 ;
    wire \current_shift_inst.un38_control_input_cry_17_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ;
    wire \current_shift_inst.un38_control_input_0_s1_19 ;
    wire \current_shift_inst.un38_control_input_cry_18_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ;
    wire \current_shift_inst.un38_control_input_0_s1_20 ;
    wire \current_shift_inst.un38_control_input_cry_19_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ;
    wire \current_shift_inst.un38_control_input_0_s1_21 ;
    wire \current_shift_inst.un38_control_input_cry_20_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ;
    wire \current_shift_inst.un38_control_input_0_s1_22 ;
    wire \current_shift_inst.un38_control_input_cry_21_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ;
    wire \current_shift_inst.un38_control_input_0_s1_23 ;
    wire \current_shift_inst.un38_control_input_cry_22_s1 ;
    wire \current_shift_inst.un38_control_input_cry_23_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ;
    wire \current_shift_inst.un38_control_input_0_s1_24 ;
    wire bfn_18_20_0_;
    wire \current_shift_inst.elapsed_time_ns_1_RNISV131_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_25 ;
    wire \current_shift_inst.un38_control_input_cry_24_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ;
    wire \current_shift_inst.un38_control_input_cry_25_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI28431_28 ;
    wire \current_shift_inst.un38_control_input_0_s1_27 ;
    wire \current_shift_inst.un38_control_input_cry_26_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ;
    wire \current_shift_inst.un38_control_input_0_s1_28 ;
    wire \current_shift_inst.un38_control_input_cry_27_s1 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ;
    wire \current_shift_inst.un38_control_input_0_s1_29 ;
    wire \current_shift_inst.un38_control_input_cry_28_s1 ;
    wire \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ;
    wire \current_shift_inst.un38_control_input_0_s1_30 ;
    wire \current_shift_inst.un38_control_input_cry_29_s1 ;
    wire \current_shift_inst.un38_control_input_5_2 ;
    wire \current_shift_inst.elapsed_time_ns_s1_31 ;
    wire \current_shift_inst.un38_control_input_cry_30_s1 ;
    wire \current_shift_inst.un38_control_input_0_s1_31 ;
    wire \current_shift_inst.un38_control_input_0_s0_26 ;
    wire \current_shift_inst.un38_control_input_0_s1_26 ;
    wire \current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ;
    wire \current_shift_inst.control_input_axb_23 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ;
    wire elapsed_time_ns_1_RNI02CN9_0_13;
    wire elapsed_time_ns_1_RNI02CN9_0_13_cascade_;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ;
    wire elapsed_time_ns_1_RNI47DN9_0_26;
    wire \phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ;
    wire elapsed_time_ns_1_RNI14DN9_0_23;
    wire \delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ;
    wire \delay_measurement_inst.delay_hc_timer.delay_hc3 ;
    wire elapsed_time_ns_1_RNI13CN9_0_14;
    wire s1_phy_c;
    wire state_3;
    wire \current_shift_inst.stop_timer_sZ0Z1 ;
    wire \current_shift_inst.start_timer_sZ0Z1 ;
    wire \current_shift_inst.timer_s1.runningZ0 ;
    wire \current_shift_inst.PI_CTRL.prop_term_1_0 ;
    wire \current_shift_inst.PI_CTRL.prop_termZ0Z_0 ;
    wire CONSTANT_ONE_NET;
    wire \current_shift_inst.elapsed_time_ns_s1_i_31 ;
    wire \current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ;
    wire \current_shift_inst.un38_control_input_5_0 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_31 ;
    wire \current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ;
    wire \current_shift_inst.PI_CTRL.N_145 ;
    wire \current_shift_inst.PI_CTRL.N_96_cascade_ ;
    wire \current_shift_inst.PI_CTRL.N_98 ;
    wire \pwm_generator_inst.un3_threshold ;
    wire \pwm_generator_inst.un3_threshold_iZ0 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ;
    wire pwm_duty_input_9;
    wire pwm_duty_input_10;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ;
    wire pwm_duty_input_1;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ;
    wire pwm_duty_input_2;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ;
    wire pwm_duty_input_6;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ;
    wire pwm_duty_input_5;
    wire \current_shift_inst.PI_CTRL.N_91 ;
    wire \current_shift_inst.PI_CTRL.N_27 ;
    wire \current_shift_inst.PI_CTRL.un7_enablelto4 ;
    wire pwm_duty_input_4;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ;
    wire pwm_duty_input_7;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ;
    wire \current_shift_inst.PI_CTRL.N_162 ;
    wire pwm_duty_input_0;
    wire \current_shift_inst.PI_CTRL.un7_enablelto3 ;
    wire \current_shift_inst.PI_CTRL.N_96 ;
    wire \current_shift_inst.PI_CTRL.N_94 ;
    wire pwm_duty_input_3;
    wire \current_shift_inst.PI_CTRL.un8_enablelto31 ;
    wire \current_shift_inst.PI_CTRL.N_160 ;
    wire \current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ;
    wire \current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ;
    wire pwm_duty_input_8;
    wire _gnd_net_;
    wire clk_100mhz_0;
    wire reset_c_g;

    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .TEST_MODE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FILTER_RANGE=3'b001;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVR=4'b0000;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVQ=3'b011;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DIVF=7'b1000010;
    defparam \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \pll_inst.ICE40_MAIN_PROGRAM_100MHZ_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(),
            .REFERENCECLK(N__24919),
            .RESETB(N__35719),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL(clk_100mhz_0));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_2_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__51645),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__51642),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15}),
            .ADDSUBBOT(),
            .A({N__37882,N__37855,N__38182,N__37822,N__37795,N__38209,N__37504,N__37969,N__38008,N__37912,N__37939,N__37276,N__37531,N__37306,N__37333,N__37357}),
            .C({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31}),
            .B({dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,N__51644,dangling_wire_45,N__51643}),
            .OHOLDTOP(),
            .O({dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ,\current_shift_inst.PI_CTRL.integrator_1_0_2_0 }));
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__51622),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__51619),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .ADDSUBBOT(),
            .A({dangling_wire_78,N__51797,N__51800,N__51798,N__51801,N__51799,N__51868,N__52663,N__53020,N__51676,N__53146,N__53062,N__52927,N__51727,N__51751,N__52990}),
            .C({dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94}),
            .B({dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,N__51621,dangling_wire_108,N__51620}),
            .OHOLDTOP(),
            .O({dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,\pwm_generator_inst.un2_threshold_1_19 ,\pwm_generator_inst.un2_threshold_1_18 ,\pwm_generator_inst.un2_threshold_1_17 ,\pwm_generator_inst.un2_threshold_1_16 ,\pwm_generator_inst.un2_threshold_1_15 ,\pwm_generator_inst.O_0_14 ,\pwm_generator_inst.O_0_13 ,\pwm_generator_inst.O_0_12 ,\pwm_generator_inst.O_0_11 ,\pwm_generator_inst.O_0_10 ,\pwm_generator_inst.O_0_9 ,\pwm_generator_inst.O_0_8 ,\pwm_generator_inst.un3_threshold ,\pwm_generator_inst.O_0_6 ,\pwm_generator_inst.O_0_5 ,\pwm_generator_inst.O_0_4 ,\pwm_generator_inst.O_0_3 ,\pwm_generator_inst.O_0_2 ,\pwm_generator_inst.O_0_1 ,\pwm_generator_inst.O_0_0 }));
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un5_threshold_1_mulonly_0_26_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__51360),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__51355),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136}),
            .ADDSUBBOT(),
            .A({dangling_wire_137,N__22822,N__22861,N__22897,N__51922,N__21625,N__21718,N__21673,N__21694,N__21646,N__21760,N__21739,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141}),
            .C({dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157}),
            .B({dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__51356,N__51372,N__51359,N__51371,N__51357,dangling_wire_164,dangling_wire_165,N__51370,N__51358,N__51369}),
            .OHOLDTOP(),
            .O({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,\pwm_generator_inst.un5_threshold_1_26 ,\pwm_generator_inst.un5_threshold_1_25 ,\pwm_generator_inst.un5_threshold_1_24 ,\pwm_generator_inst.un5_threshold_1_23 ,\pwm_generator_inst.un5_threshold_1_22 ,\pwm_generator_inst.un5_threshold_1_21 ,\pwm_generator_inst.un5_threshold_1_20 ,\pwm_generator_inst.un5_threshold_1_19 ,\pwm_generator_inst.un5_threshold_1_18 ,\pwm_generator_inst.un5_threshold_1_17 ,\pwm_generator_inst.un5_threshold_1_16 ,\pwm_generator_inst.un5_threshold_1_15 ,\pwm_generator_inst.O_14 ,\pwm_generator_inst.O_13 ,\pwm_generator_inst.O_12 ,\pwm_generator_inst.O_11 ,\pwm_generator_inst.O_10 ,\pwm_generator_inst.O_9 ,\pwm_generator_inst.O_8 ,\pwm_generator_inst.O_7 ,\pwm_generator_inst.O_6 ,\pwm_generator_inst.O_5 ,\pwm_generator_inst.O_4 ,\pwm_generator_inst.O_3 ,\pwm_generator_inst.O_2 ,\pwm_generator_inst.O_1 ,\pwm_generator_inst.O_0 }));
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un2_threshold_2_mulonly_0_16_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__51171),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__51168),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181,dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186}),
            .ADDSUBBOT(),
            .A({N__51851,N__51859,N__51850,N__51858,N__51849,N__51857,N__51848,N__51856,N__51847,N__51854,N__51846,N__51855,N__51845,N__51853,N__51844,N__51852}),
            .C({dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202}),
            .B({dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213,dangling_wire_214,dangling_wire_215,N__51170,dangling_wire_216,N__51169}),
            .OHOLDTOP(),
            .O({dangling_wire_217,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,\pwm_generator_inst.un2_threshold_2_12 ,\pwm_generator_inst.un2_threshold_2_11 ,\pwm_generator_inst.un2_threshold_2_10 ,\pwm_generator_inst.un2_threshold_2_9 ,\pwm_generator_inst.un2_threshold_2_8 ,\pwm_generator_inst.un2_threshold_2_7 ,\pwm_generator_inst.un2_threshold_2_6 ,\pwm_generator_inst.un2_threshold_2_5 ,\pwm_generator_inst.un2_threshold_2_4 ,\pwm_generator_inst.un2_threshold_2_3 ,\pwm_generator_inst.un2_threshold_2_2 ,\pwm_generator_inst.un2_threshold_2_1 ,\pwm_generator_inst.un2_threshold_2_0 }));
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .A_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .NEG_TRIGGER=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .MODE_8x8=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .D_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .C_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .B_SIGNED=1'b1;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .B_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0 .A_SIGNED=1'b1;
    SB_MAC16 \pwm_generator_inst.un5_threshold_2_1_mulonly_0_26_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__51090),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__51075),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239,dangling_wire_240,dangling_wire_241,dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251}),
            .ADDSUBBOT(),
            .A({dangling_wire_252,N__23131,N__23140,N__23152,N__22927,N__22936,N__22945,N__22954,N__22963,N__22972,N__22981,N__22990,N__22687,N__22717,N__22750,N__22786}),
            .C({dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257,dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268}),
            .B({dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,N__51076,N__51080,N__51086,N__51079,N__51084,dangling_wire_275,dangling_wire_276,N__51078,N__51085,N__51077}),
            .OHOLDTOP(),
            .O({dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,dangling_wire_283,dangling_wire_284,dangling_wire_285,dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,\pwm_generator_inst.un5_threshold_2_1_16 ,\pwm_generator_inst.un5_threshold_2_1_15 ,\pwm_generator_inst.un5_threshold_2_14 ,\pwm_generator_inst.un5_threshold_2_13 ,\pwm_generator_inst.un5_threshold_2_12 ,\pwm_generator_inst.un5_threshold_2_11 ,\pwm_generator_inst.un5_threshold_2_10 ,\pwm_generator_inst.un5_threshold_2_9 ,\pwm_generator_inst.un5_threshold_2_8 ,\pwm_generator_inst.un5_threshold_2_7 ,\pwm_generator_inst.un5_threshold_2_6 ,\pwm_generator_inst.un5_threshold_2_5 ,\pwm_generator_inst.un5_threshold_2_4 ,\pwm_generator_inst.un5_threshold_2_3 ,\pwm_generator_inst.un5_threshold_2_2 ,\pwm_generator_inst.un5_threshold_2_1 ,\pwm_generator_inst.un5_threshold_2_0 }));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOP_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .TOPADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG2=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .PIPELINE_16x16_MULT_REG1=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .NEG_TRIGGER=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .MODE_8x8=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .D_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .C_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_SIGNED=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .B_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOT_8x8_MULT_REG=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTOUTPUT_SELECT=2'b11;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_UPPERINPUT=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_LOWERINPUT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .BOTADDSUB_CARRYSELECT=2'b00;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0 .A_SIGNED=1'b1;
    SB_MAC16 \current_shift_inst.PI_CTRL.integrator_1_0_1_mulonly_0_19_0  (
            .ACCUMCO(),
            .DHOLD(),
            .AHOLD(N__51494),
            .SIGNEXTOUT(),
            .ORSTTOP(),
            .ORSTBOT(),
            .CI(),
            .IRSTTOP(),
            .ACCUMCI(),
            .OLOADBOT(),
            .CHOLD(),
            .IRSTBOT(),
            .OHOLDBOT(),
            .SIGNEXTIN(),
            .ADDSUBTOP(),
            .OLOADTOP(),
            .CE(),
            .BHOLD(N__51577),
            .CLK(GNDG0),
            .CO(),
            .D({dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301,dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,dangling_wire_306,dangling_wire_307}),
            .ADDSUBBOT(),
            .A({dangling_wire_308,N__37387,N__37417,N__37444,N__37051,N__37078,N__37102,N__37129,N__37162,N__37189,N__37216,N__37243,N__36967,N__36991,N__37018,N__50218}),
            .C({dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324}),
            .B({dangling_wire_325,dangling_wire_326,dangling_wire_327,dangling_wire_328,dangling_wire_329,dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,N__51579,dangling_wire_338,N__51578}),
            .OHOLDTOP(),
            .O({dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345,dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,dangling_wire_350,\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ,\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_15 ,\current_shift_inst.PI_CTRL.integrator_1_14 ,\current_shift_inst.PI_CTRL.integrator_1_13 ,\current_shift_inst.PI_CTRL.integrator_1_12 ,\current_shift_inst.PI_CTRL.integrator_1_11 ,\current_shift_inst.PI_CTRL.integrator_1_10 ,\current_shift_inst.PI_CTRL.integrator_1_9 ,\current_shift_inst.PI_CTRL.integrator_1_8 ,\current_shift_inst.PI_CTRL.integrator_1_7 ,\current_shift_inst.PI_CTRL.integrator_1_6 ,\current_shift_inst.PI_CTRL.integrator_1_5 ,\current_shift_inst.PI_CTRL.integrator_1_4 ,\current_shift_inst.PI_CTRL.integrator_1_3 ,\current_shift_inst.PI_CTRL.integrator_1_2 ,\current_shift_inst.PI_CTRL.un1_integrator }));
    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__53309),
            .GLOBALBUFFEROUTPUT(reset_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__53311),
            .DIN(N__53310),
            .DOUT(N__53309),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__53311),
            .PADOUT(N__53310),
            .PADIN(N__53309),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_output_obuf_iopad (
            .OE(N__53300),
            .DIN(N__53299),
            .DOUT(N__53298),
            .PACKAGEPIN(pwm_output));
    defparam pwm_output_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_output_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_output_obuf_preio (
            .PADOEN(N__53300),
            .PADOUT(N__53299),
            .PADIN(N__53298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23797),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp2_ibuf_iopad (
            .OE(N__53291),
            .DIN(N__53290),
            .DOUT(N__53289),
            .PACKAGEPIN(il_min_comp2));
    defparam il_min_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp2_ibuf_preio (
            .PADOEN(N__53291),
            .PADOUT(N__53290),
            .PADIN(N__53289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_phy_obuf_iopad (
            .OE(N__53282),
            .DIN(N__53281),
            .DOUT(N__53280),
            .PACKAGEPIN(s1_phy));
    defparam s1_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_phy_obuf_preio (
            .PADOEN(N__53282),
            .PADOUT(N__53281),
            .PADIN(N__53280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__50368),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s4_phy_obuf_iopad (
            .OE(N__53273),
            .DIN(N__53272),
            .DOUT(N__53271),
            .PACKAGEPIN(s4_phy));
    defparam s4_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s4_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s4_phy_obuf_preio (
            .PADOEN(N__53273),
            .PADOUT(N__53272),
            .PADIN(N__53271),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_min_comp1_ibuf_iopad (
            .OE(N__53264),
            .DIN(N__53263),
            .DOUT(N__53262),
            .PACKAGEPIN(il_min_comp1));
    defparam il_min_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_min_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_min_comp1_ibuf_preio (
            .PADOEN(N__53264),
            .PADOUT(N__53263),
            .PADIN(N__53262),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_min_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_phy_obuf_iopad (
            .OE(N__53255),
            .DIN(N__53254),
            .DOUT(N__53253),
            .PACKAGEPIN(s3_phy));
    defparam s3_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_phy_obuf_preio (
            .PADOEN(N__53255),
            .PADOUT(N__53254),
            .PADIN(N__53253),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__29143),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start_stop_ibuf_iopad (
            .OE(N__53246),
            .DIN(N__53245),
            .DOUT(N__53244),
            .PACKAGEPIN(start_stop));
    defparam start_stop_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam start_stop_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO start_stop_ibuf_preio (
            .PADOEN(N__53246),
            .PADOUT(N__53245),
            .PADIN(N__53244),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(start_stop_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp2_ibuf_iopad (
            .OE(N__53237),
            .DIN(N__53236),
            .DOUT(N__53235),
            .PACKAGEPIN(il_max_comp2));
    defparam il_max_comp2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp2_ibuf_preio (
            .PADOEN(N__53237),
            .PADOUT(N__53236),
            .PADIN(N__53235),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD il_max_comp1_ibuf_iopad (
            .OE(N__53228),
            .DIN(N__53227),
            .DOUT(N__53226),
            .PACKAGEPIN(il_max_comp1));
    defparam il_max_comp1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam il_max_comp1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO il_max_comp1_ibuf_preio (
            .PADOEN(N__53228),
            .PADOUT(N__53227),
            .PADIN(N__53226),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(il_max_comp1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_phy_obuf_iopad (
            .OE(N__53219),
            .DIN(N__53218),
            .DOUT(N__53217),
            .PACKAGEPIN(s2_phy));
    defparam s2_phy_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_phy_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_phy_obuf_preio (
            .PADOEN(N__53219),
            .PADOUT(N__53218),
            .PADIN(N__53217),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__38071),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_hc_input_ibuf_gb_io_iopad (
            .OE(N__53210),
            .DIN(N__53209),
            .DOUT(N__53208),
            .PACKAGEPIN(delay_hc_input));
    defparam delay_hc_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_hc_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_hc_input_ibuf_gb_io_preio (
            .PADOEN(N__53210),
            .PADOUT(N__53209),
            .PADIN(N__53208),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_hc_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD delay_tr_input_ibuf_gb_io_iopad (
            .OE(N__53201),
            .DIN(N__53200),
            .DOUT(N__53199),
            .PACKAGEPIN(delay_tr_input));
    defparam delay_tr_input_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam delay_tr_input_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO delay_tr_input_ibuf_gb_io_preio (
            .PADOEN(N__53201),
            .PADOUT(N__53200),
            .PADIN(N__53199),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(delay_tr_input_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__12303 (
            .O(N__53182),
            .I(N__53179));
    InMux I__12302 (
            .O(N__53179),
            .I(N__53176));
    LocalMux I__12301 (
            .O(N__53176),
            .I(N__53172));
    InMux I__12300 (
            .O(N__53175),
            .I(N__53169));
    Span4Mux_s2_h I__12299 (
            .O(N__53172),
            .I(N__53163));
    LocalMux I__12298 (
            .O(N__53169),
            .I(N__53163));
    InMux I__12297 (
            .O(N__53168),
            .I(N__53160));
    Span4Mux_h I__12296 (
            .O(N__53163),
            .I(N__53155));
    LocalMux I__12295 (
            .O(N__53160),
            .I(N__53155));
    Span4Mux_v I__12294 (
            .O(N__53155),
            .I(N__53152));
    Sp12to4 I__12293 (
            .O(N__53152),
            .I(N__53149));
    Odrv12 I__12292 (
            .O(N__53149),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ));
    InMux I__12291 (
            .O(N__53146),
            .I(N__53143));
    LocalMux I__12290 (
            .O(N__53143),
            .I(pwm_duty_input_5));
    InMux I__12289 (
            .O(N__53140),
            .I(N__53137));
    LocalMux I__12288 (
            .O(N__53137),
            .I(N__53134));
    Odrv4 I__12287 (
            .O(N__53134),
            .I(\current_shift_inst.PI_CTRL.N_91 ));
    CascadeMux I__12286 (
            .O(N__53131),
            .I(N__53128));
    InMux I__12285 (
            .O(N__53128),
            .I(N__53125));
    LocalMux I__12284 (
            .O(N__53125),
            .I(N__53121));
    InMux I__12283 (
            .O(N__53124),
            .I(N__53118));
    Odrv4 I__12282 (
            .O(N__53121),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    LocalMux I__12281 (
            .O(N__53118),
            .I(\current_shift_inst.PI_CTRL.N_27 ));
    CascadeMux I__12280 (
            .O(N__53113),
            .I(N__53108));
    InMux I__12279 (
            .O(N__53112),
            .I(N__53105));
    InMux I__12278 (
            .O(N__53111),
            .I(N__53099));
    InMux I__12277 (
            .O(N__53108),
            .I(N__53099));
    LocalMux I__12276 (
            .O(N__53105),
            .I(N__53096));
    InMux I__12275 (
            .O(N__53104),
            .I(N__53093));
    LocalMux I__12274 (
            .O(N__53099),
            .I(N__53090));
    Span4Mux_v I__12273 (
            .O(N__53096),
            .I(N__53085));
    LocalMux I__12272 (
            .O(N__53093),
            .I(N__53085));
    Span4Mux_h I__12271 (
            .O(N__53090),
            .I(N__53082));
    Span4Mux_h I__12270 (
            .O(N__53085),
            .I(N__53079));
    Span4Mux_h I__12269 (
            .O(N__53082),
            .I(N__53076));
    Span4Mux_h I__12268 (
            .O(N__53079),
            .I(N__53073));
    Span4Mux_h I__12267 (
            .O(N__53076),
            .I(N__53070));
    Span4Mux_h I__12266 (
            .O(N__53073),
            .I(N__53067));
    Odrv4 I__12265 (
            .O(N__53070),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    Odrv4 I__12264 (
            .O(N__53067),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto4 ));
    InMux I__12263 (
            .O(N__53062),
            .I(N__53059));
    LocalMux I__12262 (
            .O(N__53059),
            .I(pwm_duty_input_4));
    InMux I__12261 (
            .O(N__53056),
            .I(N__53053));
    LocalMux I__12260 (
            .O(N__53053),
            .I(N__53048));
    InMux I__12259 (
            .O(N__53052),
            .I(N__53045));
    InMux I__12258 (
            .O(N__53051),
            .I(N__53042));
    Span4Mux_s2_h I__12257 (
            .O(N__53048),
            .I(N__53039));
    LocalMux I__12256 (
            .O(N__53045),
            .I(N__53034));
    LocalMux I__12255 (
            .O(N__53042),
            .I(N__53034));
    Span4Mux_v I__12254 (
            .O(N__53039),
            .I(N__53031));
    Sp12to4 I__12253 (
            .O(N__53034),
            .I(N__53028));
    Sp12to4 I__12252 (
            .O(N__53031),
            .I(N__53023));
    Span12Mux_v I__12251 (
            .O(N__53028),
            .I(N__53023));
    Odrv12 I__12250 (
            .O(N__53023),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ));
    InMux I__12249 (
            .O(N__53020),
            .I(N__53017));
    LocalMux I__12248 (
            .O(N__53017),
            .I(pwm_duty_input_7));
    InMux I__12247 (
            .O(N__53014),
            .I(N__53011));
    LocalMux I__12246 (
            .O(N__53011),
            .I(N__53008));
    Odrv12 I__12245 (
            .O(N__53008),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ));
    InMux I__12244 (
            .O(N__53005),
            .I(N__52998));
    InMux I__12243 (
            .O(N__53004),
            .I(N__52998));
    InMux I__12242 (
            .O(N__53003),
            .I(N__52995));
    LocalMux I__12241 (
            .O(N__52998),
            .I(\current_shift_inst.PI_CTRL.N_162 ));
    LocalMux I__12240 (
            .O(N__52995),
            .I(\current_shift_inst.PI_CTRL.N_162 ));
    InMux I__12239 (
            .O(N__52990),
            .I(N__52987));
    LocalMux I__12238 (
            .O(N__52987),
            .I(pwm_duty_input_0));
    InMux I__12237 (
            .O(N__52984),
            .I(N__52980));
    InMux I__12236 (
            .O(N__52983),
            .I(N__52977));
    LocalMux I__12235 (
            .O(N__52980),
            .I(N__52971));
    LocalMux I__12234 (
            .O(N__52977),
            .I(N__52971));
    InMux I__12233 (
            .O(N__52976),
            .I(N__52968));
    Span4Mux_v I__12232 (
            .O(N__52971),
            .I(N__52965));
    LocalMux I__12231 (
            .O(N__52968),
            .I(N__52962));
    Span4Mux_h I__12230 (
            .O(N__52965),
            .I(N__52957));
    Span4Mux_h I__12229 (
            .O(N__52962),
            .I(N__52957));
    Span4Mux_h I__12228 (
            .O(N__52957),
            .I(N__52954));
    Span4Mux_h I__12227 (
            .O(N__52954),
            .I(N__52951));
    Odrv4 I__12226 (
            .O(N__52951),
            .I(\current_shift_inst.PI_CTRL.un7_enablelto3 ));
    InMux I__12225 (
            .O(N__52948),
            .I(N__52945));
    LocalMux I__12224 (
            .O(N__52945),
            .I(\current_shift_inst.PI_CTRL.N_96 ));
    InMux I__12223 (
            .O(N__52942),
            .I(N__52939));
    LocalMux I__12222 (
            .O(N__52939),
            .I(N__52935));
    InMux I__12221 (
            .O(N__52938),
            .I(N__52932));
    Odrv4 I__12220 (
            .O(N__52935),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    LocalMux I__12219 (
            .O(N__52932),
            .I(\current_shift_inst.PI_CTRL.N_94 ));
    InMux I__12218 (
            .O(N__52927),
            .I(N__52924));
    LocalMux I__12217 (
            .O(N__52924),
            .I(pwm_duty_input_3));
    InMux I__12216 (
            .O(N__52921),
            .I(N__52911));
    InMux I__12215 (
            .O(N__52920),
            .I(N__52911));
    InMux I__12214 (
            .O(N__52919),
            .I(N__52908));
    InMux I__12213 (
            .O(N__52918),
            .I(N__52901));
    InMux I__12212 (
            .O(N__52917),
            .I(N__52901));
    InMux I__12211 (
            .O(N__52916),
            .I(N__52901));
    LocalMux I__12210 (
            .O(N__52911),
            .I(N__52897));
    LocalMux I__12209 (
            .O(N__52908),
            .I(N__52894));
    LocalMux I__12208 (
            .O(N__52901),
            .I(N__52891));
    InMux I__12207 (
            .O(N__52900),
            .I(N__52888));
    Span4Mux_v I__12206 (
            .O(N__52897),
            .I(N__52885));
    Span4Mux_s3_h I__12205 (
            .O(N__52894),
            .I(N__52882));
    Span4Mux_s2_h I__12204 (
            .O(N__52891),
            .I(N__52877));
    LocalMux I__12203 (
            .O(N__52888),
            .I(N__52877));
    Span4Mux_v I__12202 (
            .O(N__52885),
            .I(N__52871));
    Span4Mux_v I__12201 (
            .O(N__52882),
            .I(N__52868));
    Span4Mux_v I__12200 (
            .O(N__52877),
            .I(N__52865));
    InMux I__12199 (
            .O(N__52876),
            .I(N__52858));
    InMux I__12198 (
            .O(N__52875),
            .I(N__52858));
    InMux I__12197 (
            .O(N__52874),
            .I(N__52858));
    Span4Mux_h I__12196 (
            .O(N__52871),
            .I(N__52855));
    Sp12to4 I__12195 (
            .O(N__52868),
            .I(N__52852));
    Span4Mux_v I__12194 (
            .O(N__52865),
            .I(N__52849));
    LocalMux I__12193 (
            .O(N__52858),
            .I(N__52846));
    Sp12to4 I__12192 (
            .O(N__52855),
            .I(N__52837));
    Span12Mux_s7_v I__12191 (
            .O(N__52852),
            .I(N__52837));
    Sp12to4 I__12190 (
            .O(N__52849),
            .I(N__52837));
    Span12Mux_v I__12189 (
            .O(N__52846),
            .I(N__52837));
    Odrv12 I__12188 (
            .O(N__52837),
            .I(\current_shift_inst.PI_CTRL.un8_enablelto31 ));
    InMux I__12187 (
            .O(N__52834),
            .I(N__52824));
    InMux I__12186 (
            .O(N__52833),
            .I(N__52824));
    InMux I__12185 (
            .O(N__52832),
            .I(N__52816));
    InMux I__12184 (
            .O(N__52831),
            .I(N__52816));
    InMux I__12183 (
            .O(N__52830),
            .I(N__52816));
    InMux I__12182 (
            .O(N__52829),
            .I(N__52813));
    LocalMux I__12181 (
            .O(N__52824),
            .I(N__52810));
    InMux I__12180 (
            .O(N__52823),
            .I(N__52807));
    LocalMux I__12179 (
            .O(N__52816),
            .I(N__52802));
    LocalMux I__12178 (
            .O(N__52813),
            .I(N__52802));
    Span4Mux_s2_h I__12177 (
            .O(N__52810),
            .I(N__52797));
    LocalMux I__12176 (
            .O(N__52807),
            .I(N__52797));
    Span4Mux_v I__12175 (
            .O(N__52802),
            .I(N__52794));
    Span4Mux_v I__12174 (
            .O(N__52797),
            .I(N__52791));
    Span4Mux_h I__12173 (
            .O(N__52794),
            .I(N__52788));
    Span4Mux_h I__12172 (
            .O(N__52791),
            .I(N__52785));
    Span4Mux_h I__12171 (
            .O(N__52788),
            .I(N__52782));
    Span4Mux_h I__12170 (
            .O(N__52785),
            .I(N__52779));
    Odrv4 I__12169 (
            .O(N__52782),
            .I(\current_shift_inst.PI_CTRL.N_160 ));
    Odrv4 I__12168 (
            .O(N__52779),
            .I(\current_shift_inst.PI_CTRL.N_160 ));
    CascadeMux I__12167 (
            .O(N__52774),
            .I(N__52771));
    InMux I__12166 (
            .O(N__52771),
            .I(N__52767));
    InMux I__12165 (
            .O(N__52770),
            .I(N__52764));
    LocalMux I__12164 (
            .O(N__52767),
            .I(N__52761));
    LocalMux I__12163 (
            .O(N__52764),
            .I(N__52758));
    Span4Mux_v I__12162 (
            .O(N__52761),
            .I(N__52754));
    Span4Mux_h I__12161 (
            .O(N__52758),
            .I(N__52751));
    InMux I__12160 (
            .O(N__52757),
            .I(N__52748));
    Sp12to4 I__12159 (
            .O(N__52754),
            .I(N__52745));
    Span4Mux_v I__12158 (
            .O(N__52751),
            .I(N__52742));
    LocalMux I__12157 (
            .O(N__52748),
            .I(N__52739));
    Span12Mux_s4_h I__12156 (
            .O(N__52745),
            .I(N__52732));
    Sp12to4 I__12155 (
            .O(N__52742),
            .I(N__52732));
    Span12Mux_v I__12154 (
            .O(N__52739),
            .I(N__52732));
    Odrv12 I__12153 (
            .O(N__52732),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ));
    CascadeMux I__12152 (
            .O(N__52729),
            .I(N__52723));
    CascadeMux I__12151 (
            .O(N__52728),
            .I(N__52719));
    InMux I__12150 (
            .O(N__52727),
            .I(N__52715));
    InMux I__12149 (
            .O(N__52726),
            .I(N__52710));
    InMux I__12148 (
            .O(N__52723),
            .I(N__52710));
    InMux I__12147 (
            .O(N__52722),
            .I(N__52705));
    InMux I__12146 (
            .O(N__52719),
            .I(N__52705));
    CascadeMux I__12145 (
            .O(N__52718),
            .I(N__52702));
    LocalMux I__12144 (
            .O(N__52715),
            .I(N__52697));
    LocalMux I__12143 (
            .O(N__52710),
            .I(N__52692));
    LocalMux I__12142 (
            .O(N__52705),
            .I(N__52692));
    InMux I__12141 (
            .O(N__52702),
            .I(N__52687));
    InMux I__12140 (
            .O(N__52701),
            .I(N__52687));
    InMux I__12139 (
            .O(N__52700),
            .I(N__52684));
    Span4Mux_v I__12138 (
            .O(N__52697),
            .I(N__52675));
    Span4Mux_v I__12137 (
            .O(N__52692),
            .I(N__52675));
    LocalMux I__12136 (
            .O(N__52687),
            .I(N__52675));
    LocalMux I__12135 (
            .O(N__52684),
            .I(N__52675));
    Span4Mux_h I__12134 (
            .O(N__52675),
            .I(N__52672));
    Span4Mux_v I__12133 (
            .O(N__52672),
            .I(N__52669));
    Span4Mux_h I__12132 (
            .O(N__52669),
            .I(N__52666));
    Odrv4 I__12131 (
            .O(N__52666),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ));
    InMux I__12130 (
            .O(N__52663),
            .I(N__52660));
    LocalMux I__12129 (
            .O(N__52660),
            .I(pwm_duty_input_8));
    ClkMux I__12128 (
            .O(N__52657),
            .I(N__52297));
    ClkMux I__12127 (
            .O(N__52656),
            .I(N__52297));
    ClkMux I__12126 (
            .O(N__52655),
            .I(N__52297));
    ClkMux I__12125 (
            .O(N__52654),
            .I(N__52297));
    ClkMux I__12124 (
            .O(N__52653),
            .I(N__52297));
    ClkMux I__12123 (
            .O(N__52652),
            .I(N__52297));
    ClkMux I__12122 (
            .O(N__52651),
            .I(N__52297));
    ClkMux I__12121 (
            .O(N__52650),
            .I(N__52297));
    ClkMux I__12120 (
            .O(N__52649),
            .I(N__52297));
    ClkMux I__12119 (
            .O(N__52648),
            .I(N__52297));
    ClkMux I__12118 (
            .O(N__52647),
            .I(N__52297));
    ClkMux I__12117 (
            .O(N__52646),
            .I(N__52297));
    ClkMux I__12116 (
            .O(N__52645),
            .I(N__52297));
    ClkMux I__12115 (
            .O(N__52644),
            .I(N__52297));
    ClkMux I__12114 (
            .O(N__52643),
            .I(N__52297));
    ClkMux I__12113 (
            .O(N__52642),
            .I(N__52297));
    ClkMux I__12112 (
            .O(N__52641),
            .I(N__52297));
    ClkMux I__12111 (
            .O(N__52640),
            .I(N__52297));
    ClkMux I__12110 (
            .O(N__52639),
            .I(N__52297));
    ClkMux I__12109 (
            .O(N__52638),
            .I(N__52297));
    ClkMux I__12108 (
            .O(N__52637),
            .I(N__52297));
    ClkMux I__12107 (
            .O(N__52636),
            .I(N__52297));
    ClkMux I__12106 (
            .O(N__52635),
            .I(N__52297));
    ClkMux I__12105 (
            .O(N__52634),
            .I(N__52297));
    ClkMux I__12104 (
            .O(N__52633),
            .I(N__52297));
    ClkMux I__12103 (
            .O(N__52632),
            .I(N__52297));
    ClkMux I__12102 (
            .O(N__52631),
            .I(N__52297));
    ClkMux I__12101 (
            .O(N__52630),
            .I(N__52297));
    ClkMux I__12100 (
            .O(N__52629),
            .I(N__52297));
    ClkMux I__12099 (
            .O(N__52628),
            .I(N__52297));
    ClkMux I__12098 (
            .O(N__52627),
            .I(N__52297));
    ClkMux I__12097 (
            .O(N__52626),
            .I(N__52297));
    ClkMux I__12096 (
            .O(N__52625),
            .I(N__52297));
    ClkMux I__12095 (
            .O(N__52624),
            .I(N__52297));
    ClkMux I__12094 (
            .O(N__52623),
            .I(N__52297));
    ClkMux I__12093 (
            .O(N__52622),
            .I(N__52297));
    ClkMux I__12092 (
            .O(N__52621),
            .I(N__52297));
    ClkMux I__12091 (
            .O(N__52620),
            .I(N__52297));
    ClkMux I__12090 (
            .O(N__52619),
            .I(N__52297));
    ClkMux I__12089 (
            .O(N__52618),
            .I(N__52297));
    ClkMux I__12088 (
            .O(N__52617),
            .I(N__52297));
    ClkMux I__12087 (
            .O(N__52616),
            .I(N__52297));
    ClkMux I__12086 (
            .O(N__52615),
            .I(N__52297));
    ClkMux I__12085 (
            .O(N__52614),
            .I(N__52297));
    ClkMux I__12084 (
            .O(N__52613),
            .I(N__52297));
    ClkMux I__12083 (
            .O(N__52612),
            .I(N__52297));
    ClkMux I__12082 (
            .O(N__52611),
            .I(N__52297));
    ClkMux I__12081 (
            .O(N__52610),
            .I(N__52297));
    ClkMux I__12080 (
            .O(N__52609),
            .I(N__52297));
    ClkMux I__12079 (
            .O(N__52608),
            .I(N__52297));
    ClkMux I__12078 (
            .O(N__52607),
            .I(N__52297));
    ClkMux I__12077 (
            .O(N__52606),
            .I(N__52297));
    ClkMux I__12076 (
            .O(N__52605),
            .I(N__52297));
    ClkMux I__12075 (
            .O(N__52604),
            .I(N__52297));
    ClkMux I__12074 (
            .O(N__52603),
            .I(N__52297));
    ClkMux I__12073 (
            .O(N__52602),
            .I(N__52297));
    ClkMux I__12072 (
            .O(N__52601),
            .I(N__52297));
    ClkMux I__12071 (
            .O(N__52600),
            .I(N__52297));
    ClkMux I__12070 (
            .O(N__52599),
            .I(N__52297));
    ClkMux I__12069 (
            .O(N__52598),
            .I(N__52297));
    ClkMux I__12068 (
            .O(N__52597),
            .I(N__52297));
    ClkMux I__12067 (
            .O(N__52596),
            .I(N__52297));
    ClkMux I__12066 (
            .O(N__52595),
            .I(N__52297));
    ClkMux I__12065 (
            .O(N__52594),
            .I(N__52297));
    ClkMux I__12064 (
            .O(N__52593),
            .I(N__52297));
    ClkMux I__12063 (
            .O(N__52592),
            .I(N__52297));
    ClkMux I__12062 (
            .O(N__52591),
            .I(N__52297));
    ClkMux I__12061 (
            .O(N__52590),
            .I(N__52297));
    ClkMux I__12060 (
            .O(N__52589),
            .I(N__52297));
    ClkMux I__12059 (
            .O(N__52588),
            .I(N__52297));
    ClkMux I__12058 (
            .O(N__52587),
            .I(N__52297));
    ClkMux I__12057 (
            .O(N__52586),
            .I(N__52297));
    ClkMux I__12056 (
            .O(N__52585),
            .I(N__52297));
    ClkMux I__12055 (
            .O(N__52584),
            .I(N__52297));
    ClkMux I__12054 (
            .O(N__52583),
            .I(N__52297));
    ClkMux I__12053 (
            .O(N__52582),
            .I(N__52297));
    ClkMux I__12052 (
            .O(N__52581),
            .I(N__52297));
    ClkMux I__12051 (
            .O(N__52580),
            .I(N__52297));
    ClkMux I__12050 (
            .O(N__52579),
            .I(N__52297));
    ClkMux I__12049 (
            .O(N__52578),
            .I(N__52297));
    ClkMux I__12048 (
            .O(N__52577),
            .I(N__52297));
    ClkMux I__12047 (
            .O(N__52576),
            .I(N__52297));
    ClkMux I__12046 (
            .O(N__52575),
            .I(N__52297));
    ClkMux I__12045 (
            .O(N__52574),
            .I(N__52297));
    ClkMux I__12044 (
            .O(N__52573),
            .I(N__52297));
    ClkMux I__12043 (
            .O(N__52572),
            .I(N__52297));
    ClkMux I__12042 (
            .O(N__52571),
            .I(N__52297));
    ClkMux I__12041 (
            .O(N__52570),
            .I(N__52297));
    ClkMux I__12040 (
            .O(N__52569),
            .I(N__52297));
    ClkMux I__12039 (
            .O(N__52568),
            .I(N__52297));
    ClkMux I__12038 (
            .O(N__52567),
            .I(N__52297));
    ClkMux I__12037 (
            .O(N__52566),
            .I(N__52297));
    ClkMux I__12036 (
            .O(N__52565),
            .I(N__52297));
    ClkMux I__12035 (
            .O(N__52564),
            .I(N__52297));
    ClkMux I__12034 (
            .O(N__52563),
            .I(N__52297));
    ClkMux I__12033 (
            .O(N__52562),
            .I(N__52297));
    ClkMux I__12032 (
            .O(N__52561),
            .I(N__52297));
    ClkMux I__12031 (
            .O(N__52560),
            .I(N__52297));
    ClkMux I__12030 (
            .O(N__52559),
            .I(N__52297));
    ClkMux I__12029 (
            .O(N__52558),
            .I(N__52297));
    ClkMux I__12028 (
            .O(N__52557),
            .I(N__52297));
    ClkMux I__12027 (
            .O(N__52556),
            .I(N__52297));
    ClkMux I__12026 (
            .O(N__52555),
            .I(N__52297));
    ClkMux I__12025 (
            .O(N__52554),
            .I(N__52297));
    ClkMux I__12024 (
            .O(N__52553),
            .I(N__52297));
    ClkMux I__12023 (
            .O(N__52552),
            .I(N__52297));
    ClkMux I__12022 (
            .O(N__52551),
            .I(N__52297));
    ClkMux I__12021 (
            .O(N__52550),
            .I(N__52297));
    ClkMux I__12020 (
            .O(N__52549),
            .I(N__52297));
    ClkMux I__12019 (
            .O(N__52548),
            .I(N__52297));
    ClkMux I__12018 (
            .O(N__52547),
            .I(N__52297));
    ClkMux I__12017 (
            .O(N__52546),
            .I(N__52297));
    ClkMux I__12016 (
            .O(N__52545),
            .I(N__52297));
    ClkMux I__12015 (
            .O(N__52544),
            .I(N__52297));
    ClkMux I__12014 (
            .O(N__52543),
            .I(N__52297));
    ClkMux I__12013 (
            .O(N__52542),
            .I(N__52297));
    ClkMux I__12012 (
            .O(N__52541),
            .I(N__52297));
    ClkMux I__12011 (
            .O(N__52540),
            .I(N__52297));
    ClkMux I__12010 (
            .O(N__52539),
            .I(N__52297));
    ClkMux I__12009 (
            .O(N__52538),
            .I(N__52297));
    GlobalMux I__12008 (
            .O(N__52297),
            .I(clk_100mhz_0));
    InMux I__12007 (
            .O(N__52294),
            .I(N__52287));
    InMux I__12006 (
            .O(N__52293),
            .I(N__52284));
    InMux I__12005 (
            .O(N__52292),
            .I(N__52281));
    InMux I__12004 (
            .O(N__52291),
            .I(N__52278));
    InMux I__12003 (
            .O(N__52290),
            .I(N__52275));
    LocalMux I__12002 (
            .O(N__52287),
            .I(N__52272));
    LocalMux I__12001 (
            .O(N__52284),
            .I(N__52226));
    LocalMux I__12000 (
            .O(N__52281),
            .I(N__52203));
    LocalMux I__11999 (
            .O(N__52278),
            .I(N__52200));
    LocalMux I__11998 (
            .O(N__52275),
            .I(N__52184));
    Glb2LocalMux I__11997 (
            .O(N__52272),
            .I(N__51973));
    SRMux I__11996 (
            .O(N__52271),
            .I(N__51973));
    SRMux I__11995 (
            .O(N__52270),
            .I(N__51973));
    SRMux I__11994 (
            .O(N__52269),
            .I(N__51973));
    SRMux I__11993 (
            .O(N__52268),
            .I(N__51973));
    SRMux I__11992 (
            .O(N__52267),
            .I(N__51973));
    SRMux I__11991 (
            .O(N__52266),
            .I(N__51973));
    SRMux I__11990 (
            .O(N__52265),
            .I(N__51973));
    SRMux I__11989 (
            .O(N__52264),
            .I(N__51973));
    SRMux I__11988 (
            .O(N__52263),
            .I(N__51973));
    SRMux I__11987 (
            .O(N__52262),
            .I(N__51973));
    SRMux I__11986 (
            .O(N__52261),
            .I(N__51973));
    SRMux I__11985 (
            .O(N__52260),
            .I(N__51973));
    SRMux I__11984 (
            .O(N__52259),
            .I(N__51973));
    SRMux I__11983 (
            .O(N__52258),
            .I(N__51973));
    SRMux I__11982 (
            .O(N__52257),
            .I(N__51973));
    SRMux I__11981 (
            .O(N__52256),
            .I(N__51973));
    SRMux I__11980 (
            .O(N__52255),
            .I(N__51973));
    SRMux I__11979 (
            .O(N__52254),
            .I(N__51973));
    SRMux I__11978 (
            .O(N__52253),
            .I(N__51973));
    SRMux I__11977 (
            .O(N__52252),
            .I(N__51973));
    SRMux I__11976 (
            .O(N__52251),
            .I(N__51973));
    SRMux I__11975 (
            .O(N__52250),
            .I(N__51973));
    SRMux I__11974 (
            .O(N__52249),
            .I(N__51973));
    SRMux I__11973 (
            .O(N__52248),
            .I(N__51973));
    SRMux I__11972 (
            .O(N__52247),
            .I(N__51973));
    SRMux I__11971 (
            .O(N__52246),
            .I(N__51973));
    SRMux I__11970 (
            .O(N__52245),
            .I(N__51973));
    SRMux I__11969 (
            .O(N__52244),
            .I(N__51973));
    SRMux I__11968 (
            .O(N__52243),
            .I(N__51973));
    SRMux I__11967 (
            .O(N__52242),
            .I(N__51973));
    SRMux I__11966 (
            .O(N__52241),
            .I(N__51973));
    SRMux I__11965 (
            .O(N__52240),
            .I(N__51973));
    SRMux I__11964 (
            .O(N__52239),
            .I(N__51973));
    SRMux I__11963 (
            .O(N__52238),
            .I(N__51973));
    SRMux I__11962 (
            .O(N__52237),
            .I(N__51973));
    SRMux I__11961 (
            .O(N__52236),
            .I(N__51973));
    SRMux I__11960 (
            .O(N__52235),
            .I(N__51973));
    SRMux I__11959 (
            .O(N__52234),
            .I(N__51973));
    SRMux I__11958 (
            .O(N__52233),
            .I(N__51973));
    SRMux I__11957 (
            .O(N__52232),
            .I(N__51973));
    SRMux I__11956 (
            .O(N__52231),
            .I(N__51973));
    SRMux I__11955 (
            .O(N__52230),
            .I(N__51973));
    SRMux I__11954 (
            .O(N__52229),
            .I(N__51973));
    Glb2LocalMux I__11953 (
            .O(N__52226),
            .I(N__51973));
    SRMux I__11952 (
            .O(N__52225),
            .I(N__51973));
    SRMux I__11951 (
            .O(N__52224),
            .I(N__51973));
    SRMux I__11950 (
            .O(N__52223),
            .I(N__51973));
    SRMux I__11949 (
            .O(N__52222),
            .I(N__51973));
    SRMux I__11948 (
            .O(N__52221),
            .I(N__51973));
    SRMux I__11947 (
            .O(N__52220),
            .I(N__51973));
    SRMux I__11946 (
            .O(N__52219),
            .I(N__51973));
    SRMux I__11945 (
            .O(N__52218),
            .I(N__51973));
    SRMux I__11944 (
            .O(N__52217),
            .I(N__51973));
    SRMux I__11943 (
            .O(N__52216),
            .I(N__51973));
    SRMux I__11942 (
            .O(N__52215),
            .I(N__51973));
    SRMux I__11941 (
            .O(N__52214),
            .I(N__51973));
    SRMux I__11940 (
            .O(N__52213),
            .I(N__51973));
    SRMux I__11939 (
            .O(N__52212),
            .I(N__51973));
    SRMux I__11938 (
            .O(N__52211),
            .I(N__51973));
    SRMux I__11937 (
            .O(N__52210),
            .I(N__51973));
    SRMux I__11936 (
            .O(N__52209),
            .I(N__51973));
    SRMux I__11935 (
            .O(N__52208),
            .I(N__51973));
    SRMux I__11934 (
            .O(N__52207),
            .I(N__51973));
    SRMux I__11933 (
            .O(N__52206),
            .I(N__51973));
    Glb2LocalMux I__11932 (
            .O(N__52203),
            .I(N__51973));
    Glb2LocalMux I__11931 (
            .O(N__52200),
            .I(N__51973));
    SRMux I__11930 (
            .O(N__52199),
            .I(N__51973));
    SRMux I__11929 (
            .O(N__52198),
            .I(N__51973));
    SRMux I__11928 (
            .O(N__52197),
            .I(N__51973));
    SRMux I__11927 (
            .O(N__52196),
            .I(N__51973));
    SRMux I__11926 (
            .O(N__52195),
            .I(N__51973));
    SRMux I__11925 (
            .O(N__52194),
            .I(N__51973));
    SRMux I__11924 (
            .O(N__52193),
            .I(N__51973));
    SRMux I__11923 (
            .O(N__52192),
            .I(N__51973));
    SRMux I__11922 (
            .O(N__52191),
            .I(N__51973));
    SRMux I__11921 (
            .O(N__52190),
            .I(N__51973));
    SRMux I__11920 (
            .O(N__52189),
            .I(N__51973));
    SRMux I__11919 (
            .O(N__52188),
            .I(N__51973));
    SRMux I__11918 (
            .O(N__52187),
            .I(N__51973));
    Glb2LocalMux I__11917 (
            .O(N__52184),
            .I(N__51973));
    SRMux I__11916 (
            .O(N__52183),
            .I(N__51973));
    SRMux I__11915 (
            .O(N__52182),
            .I(N__51973));
    SRMux I__11914 (
            .O(N__52181),
            .I(N__51973));
    SRMux I__11913 (
            .O(N__52180),
            .I(N__51973));
    SRMux I__11912 (
            .O(N__52179),
            .I(N__51973));
    SRMux I__11911 (
            .O(N__52178),
            .I(N__51973));
    SRMux I__11910 (
            .O(N__52177),
            .I(N__51973));
    SRMux I__11909 (
            .O(N__52176),
            .I(N__51973));
    SRMux I__11908 (
            .O(N__52175),
            .I(N__51973));
    SRMux I__11907 (
            .O(N__52174),
            .I(N__51973));
    SRMux I__11906 (
            .O(N__52173),
            .I(N__51973));
    SRMux I__11905 (
            .O(N__52172),
            .I(N__51973));
    SRMux I__11904 (
            .O(N__52171),
            .I(N__51973));
    SRMux I__11903 (
            .O(N__52170),
            .I(N__51973));
    SRMux I__11902 (
            .O(N__52169),
            .I(N__51973));
    SRMux I__11901 (
            .O(N__52168),
            .I(N__51973));
    GlobalMux I__11900 (
            .O(N__51973),
            .I(N__51970));
    gio2CtrlBuf I__11899 (
            .O(N__51970),
            .I(reset_c_g));
    InMux I__11898 (
            .O(N__51967),
            .I(N__51964));
    LocalMux I__11897 (
            .O(N__51964),
            .I(\current_shift_inst.PI_CTRL.N_145 ));
    CascadeMux I__11896 (
            .O(N__51961),
            .I(\current_shift_inst.PI_CTRL.N_96_cascade_ ));
    CascadeMux I__11895 (
            .O(N__51958),
            .I(N__51955));
    InMux I__11894 (
            .O(N__51955),
            .I(N__51952));
    LocalMux I__11893 (
            .O(N__51952),
            .I(\current_shift_inst.PI_CTRL.N_98 ));
    InMux I__11892 (
            .O(N__51949),
            .I(N__51946));
    LocalMux I__11891 (
            .O(N__51946),
            .I(N__51942));
    InMux I__11890 (
            .O(N__51945),
            .I(N__51939));
    Span12Mux_s8_v I__11889 (
            .O(N__51942),
            .I(N__51936));
    LocalMux I__11888 (
            .O(N__51939),
            .I(N__51933));
    Span12Mux_h I__11887 (
            .O(N__51936),
            .I(N__51930));
    Sp12to4 I__11886 (
            .O(N__51933),
            .I(N__51925));
    Span12Mux_h I__11885 (
            .O(N__51930),
            .I(N__51925));
    Odrv12 I__11884 (
            .O(N__51925),
            .I(\pwm_generator_inst.un3_threshold ));
    InMux I__11883 (
            .O(N__51922),
            .I(N__51919));
    LocalMux I__11882 (
            .O(N__51919),
            .I(N__51916));
    Span12Mux_v I__11881 (
            .O(N__51916),
            .I(N__51913));
    Span12Mux_h I__11880 (
            .O(N__51913),
            .I(N__51910));
    Span12Mux_h I__11879 (
            .O(N__51910),
            .I(N__51907));
    Odrv12 I__11878 (
            .O(N__51907),
            .I(\pwm_generator_inst.un3_threshold_iZ0 ));
    InMux I__11877 (
            .O(N__51904),
            .I(N__51900));
    InMux I__11876 (
            .O(N__51903),
            .I(N__51897));
    LocalMux I__11875 (
            .O(N__51900),
            .I(N__51894));
    LocalMux I__11874 (
            .O(N__51897),
            .I(N__51891));
    Span4Mux_v I__11873 (
            .O(N__51894),
            .I(N__51887));
    Span4Mux_v I__11872 (
            .O(N__51891),
            .I(N__51884));
    InMux I__11871 (
            .O(N__51890),
            .I(N__51881));
    Sp12to4 I__11870 (
            .O(N__51887),
            .I(N__51874));
    Sp12to4 I__11869 (
            .O(N__51884),
            .I(N__51874));
    LocalMux I__11868 (
            .O(N__51881),
            .I(N__51874));
    Span12Mux_h I__11867 (
            .O(N__51874),
            .I(N__51871));
    Odrv12 I__11866 (
            .O(N__51871),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ));
    InMux I__11865 (
            .O(N__51868),
            .I(N__51865));
    LocalMux I__11864 (
            .O(N__51865),
            .I(N__51862));
    Odrv4 I__11863 (
            .O(N__51862),
            .I(pwm_duty_input_9));
    InMux I__11862 (
            .O(N__51859),
            .I(N__51827));
    InMux I__11861 (
            .O(N__51858),
            .I(N__51827));
    InMux I__11860 (
            .O(N__51857),
            .I(N__51827));
    InMux I__11859 (
            .O(N__51856),
            .I(N__51827));
    InMux I__11858 (
            .O(N__51855),
            .I(N__51827));
    InMux I__11857 (
            .O(N__51854),
            .I(N__51827));
    InMux I__11856 (
            .O(N__51853),
            .I(N__51827));
    InMux I__11855 (
            .O(N__51852),
            .I(N__51827));
    InMux I__11854 (
            .O(N__51851),
            .I(N__51810));
    InMux I__11853 (
            .O(N__51850),
            .I(N__51810));
    InMux I__11852 (
            .O(N__51849),
            .I(N__51810));
    InMux I__11851 (
            .O(N__51848),
            .I(N__51810));
    InMux I__11850 (
            .O(N__51847),
            .I(N__51810));
    InMux I__11849 (
            .O(N__51846),
            .I(N__51810));
    InMux I__11848 (
            .O(N__51845),
            .I(N__51810));
    InMux I__11847 (
            .O(N__51844),
            .I(N__51810));
    LocalMux I__11846 (
            .O(N__51827),
            .I(N__51805));
    LocalMux I__11845 (
            .O(N__51810),
            .I(N__51805));
    Span12Mux_v I__11844 (
            .O(N__51805),
            .I(N__51802));
    Span12Mux_h I__11843 (
            .O(N__51802),
            .I(N__51794));
    InMux I__11842 (
            .O(N__51801),
            .I(N__51789));
    InMux I__11841 (
            .O(N__51800),
            .I(N__51789));
    InMux I__11840 (
            .O(N__51799),
            .I(N__51782));
    InMux I__11839 (
            .O(N__51798),
            .I(N__51782));
    InMux I__11838 (
            .O(N__51797),
            .I(N__51782));
    Span12Mux_h I__11837 (
            .O(N__51794),
            .I(N__51779));
    LocalMux I__11836 (
            .O(N__51789),
            .I(N__51774));
    LocalMux I__11835 (
            .O(N__51782),
            .I(N__51774));
    Odrv12 I__11834 (
            .O(N__51779),
            .I(pwm_duty_input_10));
    Odrv4 I__11833 (
            .O(N__51774),
            .I(pwm_duty_input_10));
    InMux I__11832 (
            .O(N__51769),
            .I(N__51766));
    LocalMux I__11831 (
            .O(N__51766),
            .I(N__51763));
    Span4Mux_h I__11830 (
            .O(N__51763),
            .I(N__51760));
    Span4Mux_v I__11829 (
            .O(N__51760),
            .I(N__51757));
    Sp12to4 I__11828 (
            .O(N__51757),
            .I(N__51754));
    Odrv12 I__11827 (
            .O(N__51754),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ));
    InMux I__11826 (
            .O(N__51751),
            .I(N__51748));
    LocalMux I__11825 (
            .O(N__51748),
            .I(N__51745));
    Odrv4 I__11824 (
            .O(N__51745),
            .I(pwm_duty_input_1));
    InMux I__11823 (
            .O(N__51742),
            .I(N__51739));
    LocalMux I__11822 (
            .O(N__51739),
            .I(N__51736));
    Span12Mux_v I__11821 (
            .O(N__51736),
            .I(N__51733));
    Span12Mux_h I__11820 (
            .O(N__51733),
            .I(N__51730));
    Odrv12 I__11819 (
            .O(N__51730),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ));
    InMux I__11818 (
            .O(N__51727),
            .I(N__51724));
    LocalMux I__11817 (
            .O(N__51724),
            .I(N__51721));
    Span4Mux_v I__11816 (
            .O(N__51721),
            .I(N__51718));
    Odrv4 I__11815 (
            .O(N__51718),
            .I(pwm_duty_input_2));
    CascadeMux I__11814 (
            .O(N__51715),
            .I(N__51712));
    InMux I__11813 (
            .O(N__51712),
            .I(N__51708));
    CascadeMux I__11812 (
            .O(N__51711),
            .I(N__51705));
    LocalMux I__11811 (
            .O(N__51708),
            .I(N__51701));
    InMux I__11810 (
            .O(N__51705),
            .I(N__51698));
    InMux I__11809 (
            .O(N__51704),
            .I(N__51695));
    Span4Mux_v I__11808 (
            .O(N__51701),
            .I(N__51688));
    LocalMux I__11807 (
            .O(N__51698),
            .I(N__51688));
    LocalMux I__11806 (
            .O(N__51695),
            .I(N__51688));
    Span4Mux_h I__11805 (
            .O(N__51688),
            .I(N__51685));
    Span4Mux_h I__11804 (
            .O(N__51685),
            .I(N__51682));
    Span4Mux_h I__11803 (
            .O(N__51682),
            .I(N__51679));
    Odrv4 I__11802 (
            .O(N__51679),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ));
    InMux I__11801 (
            .O(N__51676),
            .I(N__51673));
    LocalMux I__11800 (
            .O(N__51673),
            .I(N__51670));
    Odrv4 I__11799 (
            .O(N__51670),
            .I(pwm_duty_input_6));
    InMux I__11798 (
            .O(N__51667),
            .I(N__51664));
    LocalMux I__11797 (
            .O(N__51664),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ));
    CascadeMux I__11796 (
            .O(N__51661),
            .I(N__51656));
    CascadeMux I__11795 (
            .O(N__51660),
            .I(N__51653));
    CascadeMux I__11794 (
            .O(N__51659),
            .I(N__51650));
    InMux I__11793 (
            .O(N__51656),
            .I(N__51635));
    InMux I__11792 (
            .O(N__51653),
            .I(N__51635));
    InMux I__11791 (
            .O(N__51650),
            .I(N__51635));
    CascadeMux I__11790 (
            .O(N__51649),
            .I(N__51632));
    CascadeMux I__11789 (
            .O(N__51648),
            .I(N__51629));
    CascadeMux I__11788 (
            .O(N__51647),
            .I(N__51626));
    CascadeMux I__11787 (
            .O(N__51646),
            .I(N__51623));
    InMux I__11786 (
            .O(N__51645),
            .I(N__51616));
    InMux I__11785 (
            .O(N__51644),
            .I(N__51611));
    InMux I__11784 (
            .O(N__51643),
            .I(N__51611));
    InMux I__11783 (
            .O(N__51642),
            .I(N__51608));
    LocalMux I__11782 (
            .O(N__51635),
            .I(N__51601));
    InMux I__11781 (
            .O(N__51632),
            .I(N__51592));
    InMux I__11780 (
            .O(N__51629),
            .I(N__51592));
    InMux I__11779 (
            .O(N__51626),
            .I(N__51592));
    InMux I__11778 (
            .O(N__51623),
            .I(N__51592));
    InMux I__11777 (
            .O(N__51622),
            .I(N__51574));
    InMux I__11776 (
            .O(N__51621),
            .I(N__51569));
    InMux I__11775 (
            .O(N__51620),
            .I(N__51569));
    InMux I__11774 (
            .O(N__51619),
            .I(N__51566));
    LocalMux I__11773 (
            .O(N__51616),
            .I(N__51559));
    LocalMux I__11772 (
            .O(N__51611),
            .I(N__51559));
    LocalMux I__11771 (
            .O(N__51608),
            .I(N__51559));
    CascadeMux I__11770 (
            .O(N__51607),
            .I(N__51556));
    CascadeMux I__11769 (
            .O(N__51606),
            .I(N__51553));
    CascadeMux I__11768 (
            .O(N__51605),
            .I(N__51550));
    CascadeMux I__11767 (
            .O(N__51604),
            .I(N__51547));
    Span4Mux_v I__11766 (
            .O(N__51601),
            .I(N__51544));
    LocalMux I__11765 (
            .O(N__51592),
            .I(N__51541));
    CascadeMux I__11764 (
            .O(N__51591),
            .I(N__51538));
    CascadeMux I__11763 (
            .O(N__51590),
            .I(N__51535));
    CascadeMux I__11762 (
            .O(N__51589),
            .I(N__51532));
    CascadeMux I__11761 (
            .O(N__51588),
            .I(N__51529));
    CascadeMux I__11760 (
            .O(N__51587),
            .I(N__51526));
    CascadeMux I__11759 (
            .O(N__51586),
            .I(N__51523));
    CascadeMux I__11758 (
            .O(N__51585),
            .I(N__51520));
    CascadeMux I__11757 (
            .O(N__51584),
            .I(N__51517));
    CascadeMux I__11756 (
            .O(N__51583),
            .I(N__51514));
    CascadeMux I__11755 (
            .O(N__51582),
            .I(N__51511));
    CascadeMux I__11754 (
            .O(N__51581),
            .I(N__51508));
    CascadeMux I__11753 (
            .O(N__51580),
            .I(N__51505));
    InMux I__11752 (
            .O(N__51579),
            .I(N__51489));
    InMux I__11751 (
            .O(N__51578),
            .I(N__51489));
    InMux I__11750 (
            .O(N__51577),
            .I(N__51486));
    LocalMux I__11749 (
            .O(N__51574),
            .I(N__51479));
    LocalMux I__11748 (
            .O(N__51569),
            .I(N__51479));
    LocalMux I__11747 (
            .O(N__51566),
            .I(N__51479));
    Span4Mux_v I__11746 (
            .O(N__51559),
            .I(N__51476));
    InMux I__11745 (
            .O(N__51556),
            .I(N__51454));
    InMux I__11744 (
            .O(N__51553),
            .I(N__51454));
    InMux I__11743 (
            .O(N__51550),
            .I(N__51454));
    InMux I__11742 (
            .O(N__51547),
            .I(N__51454));
    Span4Mux_h I__11741 (
            .O(N__51544),
            .I(N__51449));
    Span4Mux_v I__11740 (
            .O(N__51541),
            .I(N__51449));
    InMux I__11739 (
            .O(N__51538),
            .I(N__51440));
    InMux I__11738 (
            .O(N__51535),
            .I(N__51440));
    InMux I__11737 (
            .O(N__51532),
            .I(N__51440));
    InMux I__11736 (
            .O(N__51529),
            .I(N__51440));
    InMux I__11735 (
            .O(N__51526),
            .I(N__51431));
    InMux I__11734 (
            .O(N__51523),
            .I(N__51431));
    InMux I__11733 (
            .O(N__51520),
            .I(N__51431));
    InMux I__11732 (
            .O(N__51517),
            .I(N__51431));
    InMux I__11731 (
            .O(N__51514),
            .I(N__51422));
    InMux I__11730 (
            .O(N__51511),
            .I(N__51422));
    InMux I__11729 (
            .O(N__51508),
            .I(N__51422));
    InMux I__11728 (
            .O(N__51505),
            .I(N__51422));
    CascadeMux I__11727 (
            .O(N__51504),
            .I(N__51414));
    CascadeMux I__11726 (
            .O(N__51503),
            .I(N__51410));
    CascadeMux I__11725 (
            .O(N__51502),
            .I(N__51406));
    CascadeMux I__11724 (
            .O(N__51501),
            .I(N__51402));
    CascadeMux I__11723 (
            .O(N__51500),
            .I(N__51398));
    CascadeMux I__11722 (
            .O(N__51499),
            .I(N__51394));
    CascadeMux I__11721 (
            .O(N__51498),
            .I(N__51390));
    CascadeMux I__11720 (
            .O(N__51497),
            .I(N__51383));
    CascadeMux I__11719 (
            .O(N__51496),
            .I(N__51380));
    CascadeMux I__11718 (
            .O(N__51495),
            .I(N__51377));
    InMux I__11717 (
            .O(N__51494),
            .I(N__51366));
    LocalMux I__11716 (
            .O(N__51489),
            .I(N__51361));
    LocalMux I__11715 (
            .O(N__51486),
            .I(N__51361));
    Span4Mux_v I__11714 (
            .O(N__51479),
            .I(N__51352));
    Span4Mux_h I__11713 (
            .O(N__51476),
            .I(N__51349));
    InMux I__11712 (
            .O(N__51475),
            .I(N__51346));
    CascadeMux I__11711 (
            .O(N__51474),
            .I(N__51335));
    CascadeMux I__11710 (
            .O(N__51473),
            .I(N__51332));
    CascadeMux I__11709 (
            .O(N__51472),
            .I(N__51329));
    CascadeMux I__11708 (
            .O(N__51471),
            .I(N__51326));
    CascadeMux I__11707 (
            .O(N__51470),
            .I(N__51323));
    CascadeMux I__11706 (
            .O(N__51469),
            .I(N__51320));
    CascadeMux I__11705 (
            .O(N__51468),
            .I(N__51317));
    CascadeMux I__11704 (
            .O(N__51467),
            .I(N__51314));
    CascadeMux I__11703 (
            .O(N__51466),
            .I(N__51311));
    CascadeMux I__11702 (
            .O(N__51465),
            .I(N__51308));
    CascadeMux I__11701 (
            .O(N__51464),
            .I(N__51305));
    CascadeMux I__11700 (
            .O(N__51463),
            .I(N__51302));
    LocalMux I__11699 (
            .O(N__51454),
            .I(N__51286));
    Span4Mux_v I__11698 (
            .O(N__51449),
            .I(N__51277));
    LocalMux I__11697 (
            .O(N__51440),
            .I(N__51277));
    LocalMux I__11696 (
            .O(N__51431),
            .I(N__51277));
    LocalMux I__11695 (
            .O(N__51422),
            .I(N__51277));
    CascadeMux I__11694 (
            .O(N__51421),
            .I(N__51274));
    CascadeMux I__11693 (
            .O(N__51420),
            .I(N__51271));
    CascadeMux I__11692 (
            .O(N__51419),
            .I(N__51268));
    CascadeMux I__11691 (
            .O(N__51418),
            .I(N__51265));
    InMux I__11690 (
            .O(N__51417),
            .I(N__51250));
    InMux I__11689 (
            .O(N__51414),
            .I(N__51250));
    InMux I__11688 (
            .O(N__51413),
            .I(N__51250));
    InMux I__11687 (
            .O(N__51410),
            .I(N__51250));
    InMux I__11686 (
            .O(N__51409),
            .I(N__51250));
    InMux I__11685 (
            .O(N__51406),
            .I(N__51250));
    InMux I__11684 (
            .O(N__51405),
            .I(N__51250));
    InMux I__11683 (
            .O(N__51402),
            .I(N__51233));
    InMux I__11682 (
            .O(N__51401),
            .I(N__51233));
    InMux I__11681 (
            .O(N__51398),
            .I(N__51233));
    InMux I__11680 (
            .O(N__51397),
            .I(N__51233));
    InMux I__11679 (
            .O(N__51394),
            .I(N__51233));
    InMux I__11678 (
            .O(N__51393),
            .I(N__51233));
    InMux I__11677 (
            .O(N__51390),
            .I(N__51233));
    InMux I__11676 (
            .O(N__51389),
            .I(N__51233));
    CascadeMux I__11675 (
            .O(N__51388),
            .I(N__51229));
    CascadeMux I__11674 (
            .O(N__51387),
            .I(N__51225));
    CascadeMux I__11673 (
            .O(N__51386),
            .I(N__51221));
    InMux I__11672 (
            .O(N__51383),
            .I(N__51213));
    InMux I__11671 (
            .O(N__51380),
            .I(N__51213));
    InMux I__11670 (
            .O(N__51377),
            .I(N__51213));
    CascadeMux I__11669 (
            .O(N__51376),
            .I(N__51210));
    CascadeMux I__11668 (
            .O(N__51375),
            .I(N__51207));
    CascadeMux I__11667 (
            .O(N__51374),
            .I(N__51204));
    CascadeMux I__11666 (
            .O(N__51373),
            .I(N__51201));
    InMux I__11665 (
            .O(N__51372),
            .I(N__51192));
    InMux I__11664 (
            .O(N__51371),
            .I(N__51192));
    InMux I__11663 (
            .O(N__51370),
            .I(N__51192));
    InMux I__11662 (
            .O(N__51369),
            .I(N__51192));
    LocalMux I__11661 (
            .O(N__51366),
            .I(N__51189));
    Span4Mux_s1_h I__11660 (
            .O(N__51361),
            .I(N__51186));
    InMux I__11659 (
            .O(N__51360),
            .I(N__51183));
    InMux I__11658 (
            .O(N__51359),
            .I(N__51172));
    InMux I__11657 (
            .O(N__51358),
            .I(N__51172));
    InMux I__11656 (
            .O(N__51357),
            .I(N__51172));
    InMux I__11655 (
            .O(N__51356),
            .I(N__51172));
    InMux I__11654 (
            .O(N__51355),
            .I(N__51172));
    Span4Mux_h I__11653 (
            .O(N__51352),
            .I(N__51161));
    Span4Mux_v I__11652 (
            .O(N__51349),
            .I(N__51161));
    LocalMux I__11651 (
            .O(N__51346),
            .I(N__51161));
    InMux I__11650 (
            .O(N__51345),
            .I(N__51152));
    InMux I__11649 (
            .O(N__51344),
            .I(N__51152));
    InMux I__11648 (
            .O(N__51343),
            .I(N__51152));
    InMux I__11647 (
            .O(N__51342),
            .I(N__51152));
    InMux I__11646 (
            .O(N__51341),
            .I(N__51143));
    InMux I__11645 (
            .O(N__51340),
            .I(N__51143));
    InMux I__11644 (
            .O(N__51339),
            .I(N__51143));
    InMux I__11643 (
            .O(N__51338),
            .I(N__51143));
    InMux I__11642 (
            .O(N__51335),
            .I(N__51133));
    InMux I__11641 (
            .O(N__51332),
            .I(N__51133));
    InMux I__11640 (
            .O(N__51329),
            .I(N__51133));
    InMux I__11639 (
            .O(N__51326),
            .I(N__51133));
    InMux I__11638 (
            .O(N__51323),
            .I(N__51124));
    InMux I__11637 (
            .O(N__51320),
            .I(N__51124));
    InMux I__11636 (
            .O(N__51317),
            .I(N__51124));
    InMux I__11635 (
            .O(N__51314),
            .I(N__51124));
    InMux I__11634 (
            .O(N__51311),
            .I(N__51115));
    InMux I__11633 (
            .O(N__51308),
            .I(N__51115));
    InMux I__11632 (
            .O(N__51305),
            .I(N__51115));
    InMux I__11631 (
            .O(N__51302),
            .I(N__51115));
    CascadeMux I__11630 (
            .O(N__51301),
            .I(N__51112));
    CascadeMux I__11629 (
            .O(N__51300),
            .I(N__51109));
    CascadeMux I__11628 (
            .O(N__51299),
            .I(N__51106));
    CascadeMux I__11627 (
            .O(N__51298),
            .I(N__51103));
    CascadeMux I__11626 (
            .O(N__51297),
            .I(N__51100));
    CascadeMux I__11625 (
            .O(N__51296),
            .I(N__51097));
    CascadeMux I__11624 (
            .O(N__51295),
            .I(N__51094));
    CascadeMux I__11623 (
            .O(N__51294),
            .I(N__51091));
    InMux I__11622 (
            .O(N__51293),
            .I(N__51087));
    InMux I__11621 (
            .O(N__51292),
            .I(N__51081));
    CascadeMux I__11620 (
            .O(N__51291),
            .I(N__51071));
    CascadeMux I__11619 (
            .O(N__51290),
            .I(N__51067));
    CascadeMux I__11618 (
            .O(N__51289),
            .I(N__51063));
    Span4Mux_v I__11617 (
            .O(N__51286),
            .I(N__51055));
    Span4Mux_v I__11616 (
            .O(N__51277),
            .I(N__51055));
    InMux I__11615 (
            .O(N__51274),
            .I(N__51050));
    InMux I__11614 (
            .O(N__51271),
            .I(N__51050));
    InMux I__11613 (
            .O(N__51268),
            .I(N__51045));
    InMux I__11612 (
            .O(N__51265),
            .I(N__51045));
    LocalMux I__11611 (
            .O(N__51250),
            .I(N__51040));
    LocalMux I__11610 (
            .O(N__51233),
            .I(N__51040));
    InMux I__11609 (
            .O(N__51232),
            .I(N__51025));
    InMux I__11608 (
            .O(N__51229),
            .I(N__51025));
    InMux I__11607 (
            .O(N__51228),
            .I(N__51025));
    InMux I__11606 (
            .O(N__51225),
            .I(N__51025));
    InMux I__11605 (
            .O(N__51224),
            .I(N__51025));
    InMux I__11604 (
            .O(N__51221),
            .I(N__51025));
    InMux I__11603 (
            .O(N__51220),
            .I(N__51025));
    LocalMux I__11602 (
            .O(N__51213),
            .I(N__51022));
    InMux I__11601 (
            .O(N__51210),
            .I(N__51013));
    InMux I__11600 (
            .O(N__51207),
            .I(N__51013));
    InMux I__11599 (
            .O(N__51204),
            .I(N__51013));
    InMux I__11598 (
            .O(N__51201),
            .I(N__51013));
    LocalMux I__11597 (
            .O(N__51192),
            .I(N__51010));
    Span4Mux_v I__11596 (
            .O(N__51189),
            .I(N__51001));
    Span4Mux_v I__11595 (
            .O(N__51186),
            .I(N__51001));
    LocalMux I__11594 (
            .O(N__51183),
            .I(N__51001));
    LocalMux I__11593 (
            .O(N__51172),
            .I(N__51001));
    InMux I__11592 (
            .O(N__51171),
            .I(N__50998));
    InMux I__11591 (
            .O(N__51170),
            .I(N__50993));
    InMux I__11590 (
            .O(N__51169),
            .I(N__50993));
    InMux I__11589 (
            .O(N__51168),
            .I(N__50990));
    Span4Mux_h I__11588 (
            .O(N__51161),
            .I(N__50982));
    LocalMux I__11587 (
            .O(N__51152),
            .I(N__50982));
    LocalMux I__11586 (
            .O(N__51143),
            .I(N__50982));
    InMux I__11585 (
            .O(N__51142),
            .I(N__50979));
    LocalMux I__11584 (
            .O(N__51133),
            .I(N__50976));
    LocalMux I__11583 (
            .O(N__51124),
            .I(N__50971));
    LocalMux I__11582 (
            .O(N__51115),
            .I(N__50971));
    InMux I__11581 (
            .O(N__51112),
            .I(N__50962));
    InMux I__11580 (
            .O(N__51109),
            .I(N__50962));
    InMux I__11579 (
            .O(N__51106),
            .I(N__50962));
    InMux I__11578 (
            .O(N__51103),
            .I(N__50962));
    InMux I__11577 (
            .O(N__51100),
            .I(N__50957));
    InMux I__11576 (
            .O(N__51097),
            .I(N__50957));
    InMux I__11575 (
            .O(N__51094),
            .I(N__50952));
    InMux I__11574 (
            .O(N__51091),
            .I(N__50952));
    InMux I__11573 (
            .O(N__51090),
            .I(N__50949));
    LocalMux I__11572 (
            .O(N__51087),
            .I(N__50946));
    InMux I__11571 (
            .O(N__51086),
            .I(N__50939));
    InMux I__11570 (
            .O(N__51085),
            .I(N__50939));
    InMux I__11569 (
            .O(N__51084),
            .I(N__50939));
    LocalMux I__11568 (
            .O(N__51081),
            .I(N__50936));
    InMux I__11567 (
            .O(N__51080),
            .I(N__50927));
    InMux I__11566 (
            .O(N__51079),
            .I(N__50927));
    InMux I__11565 (
            .O(N__51078),
            .I(N__50927));
    InMux I__11564 (
            .O(N__51077),
            .I(N__50927));
    InMux I__11563 (
            .O(N__51076),
            .I(N__50922));
    InMux I__11562 (
            .O(N__51075),
            .I(N__50922));
    InMux I__11561 (
            .O(N__51074),
            .I(N__50907));
    InMux I__11560 (
            .O(N__51071),
            .I(N__50907));
    InMux I__11559 (
            .O(N__51070),
            .I(N__50907));
    InMux I__11558 (
            .O(N__51067),
            .I(N__50907));
    InMux I__11557 (
            .O(N__51066),
            .I(N__50907));
    InMux I__11556 (
            .O(N__51063),
            .I(N__50907));
    InMux I__11555 (
            .O(N__51062),
            .I(N__50907));
    CascadeMux I__11554 (
            .O(N__51061),
            .I(N__50904));
    CascadeMux I__11553 (
            .O(N__51060),
            .I(N__50901));
    Sp12to4 I__11552 (
            .O(N__51055),
            .I(N__50893));
    LocalMux I__11551 (
            .O(N__51050),
            .I(N__50893));
    LocalMux I__11550 (
            .O(N__51045),
            .I(N__50893));
    Span4Mux_v I__11549 (
            .O(N__51040),
            .I(N__50888));
    LocalMux I__11548 (
            .O(N__51025),
            .I(N__50888));
    Span4Mux_h I__11547 (
            .O(N__51022),
            .I(N__50885));
    LocalMux I__11546 (
            .O(N__51013),
            .I(N__50882));
    Span4Mux_v I__11545 (
            .O(N__51010),
            .I(N__50871));
    Span4Mux_v I__11544 (
            .O(N__51001),
            .I(N__50871));
    LocalMux I__11543 (
            .O(N__50998),
            .I(N__50871));
    LocalMux I__11542 (
            .O(N__50993),
            .I(N__50871));
    LocalMux I__11541 (
            .O(N__50990),
            .I(N__50871));
    InMux I__11540 (
            .O(N__50989),
            .I(N__50868));
    Span4Mux_h I__11539 (
            .O(N__50982),
            .I(N__50863));
    LocalMux I__11538 (
            .O(N__50979),
            .I(N__50863));
    Span4Mux_v I__11537 (
            .O(N__50976),
            .I(N__50852));
    Span4Mux_h I__11536 (
            .O(N__50971),
            .I(N__50852));
    LocalMux I__11535 (
            .O(N__50962),
            .I(N__50852));
    LocalMux I__11534 (
            .O(N__50957),
            .I(N__50852));
    LocalMux I__11533 (
            .O(N__50952),
            .I(N__50852));
    LocalMux I__11532 (
            .O(N__50949),
            .I(N__50849));
    Span4Mux_v I__11531 (
            .O(N__50946),
            .I(N__50844));
    LocalMux I__11530 (
            .O(N__50939),
            .I(N__50844));
    Span4Mux_v I__11529 (
            .O(N__50936),
            .I(N__50837));
    LocalMux I__11528 (
            .O(N__50927),
            .I(N__50837));
    LocalMux I__11527 (
            .O(N__50922),
            .I(N__50837));
    LocalMux I__11526 (
            .O(N__50907),
            .I(N__50834));
    InMux I__11525 (
            .O(N__50904),
            .I(N__50827));
    InMux I__11524 (
            .O(N__50901),
            .I(N__50827));
    InMux I__11523 (
            .O(N__50900),
            .I(N__50827));
    Span12Mux_h I__11522 (
            .O(N__50893),
            .I(N__50824));
    Span4Mux_v I__11521 (
            .O(N__50888),
            .I(N__50821));
    Span4Mux_v I__11520 (
            .O(N__50885),
            .I(N__50818));
    Span4Mux_v I__11519 (
            .O(N__50882),
            .I(N__50815));
    Span4Mux_v I__11518 (
            .O(N__50871),
            .I(N__50810));
    LocalMux I__11517 (
            .O(N__50868),
            .I(N__50810));
    Span4Mux_h I__11516 (
            .O(N__50863),
            .I(N__50805));
    Span4Mux_v I__11515 (
            .O(N__50852),
            .I(N__50805));
    Span4Mux_v I__11514 (
            .O(N__50849),
            .I(N__50800));
    Span4Mux_v I__11513 (
            .O(N__50844),
            .I(N__50800));
    Span4Mux_v I__11512 (
            .O(N__50837),
            .I(N__50797));
    Span4Mux_v I__11511 (
            .O(N__50834),
            .I(N__50794));
    LocalMux I__11510 (
            .O(N__50827),
            .I(N__50791));
    Span12Mux_v I__11509 (
            .O(N__50824),
            .I(N__50786));
    Sp12to4 I__11508 (
            .O(N__50821),
            .I(N__50786));
    Span4Mux_v I__11507 (
            .O(N__50818),
            .I(N__50783));
    Span4Mux_h I__11506 (
            .O(N__50815),
            .I(N__50778));
    Span4Mux_h I__11505 (
            .O(N__50810),
            .I(N__50778));
    Span4Mux_v I__11504 (
            .O(N__50805),
            .I(N__50771));
    Span4Mux_h I__11503 (
            .O(N__50800),
            .I(N__50771));
    Span4Mux_h I__11502 (
            .O(N__50797),
            .I(N__50771));
    Span4Mux_v I__11501 (
            .O(N__50794),
            .I(N__50766));
    Span4Mux_v I__11500 (
            .O(N__50791),
            .I(N__50766));
    Odrv12 I__11499 (
            .O(N__50786),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11498 (
            .O(N__50783),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11497 (
            .O(N__50778),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11496 (
            .O(N__50771),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__11495 (
            .O(N__50766),
            .I(CONSTANT_ONE_NET));
    InMux I__11494 (
            .O(N__50755),
            .I(N__50751));
    InMux I__11493 (
            .O(N__50754),
            .I(N__50745));
    LocalMux I__11492 (
            .O(N__50751),
            .I(N__50741));
    InMux I__11491 (
            .O(N__50750),
            .I(N__50736));
    InMux I__11490 (
            .O(N__50749),
            .I(N__50736));
    InMux I__11489 (
            .O(N__50748),
            .I(N__50733));
    LocalMux I__11488 (
            .O(N__50745),
            .I(N__50730));
    InMux I__11487 (
            .O(N__50744),
            .I(N__50727));
    Span4Mux_v I__11486 (
            .O(N__50741),
            .I(N__50722));
    LocalMux I__11485 (
            .O(N__50736),
            .I(N__50722));
    LocalMux I__11484 (
            .O(N__50733),
            .I(N__50719));
    Span4Mux_h I__11483 (
            .O(N__50730),
            .I(N__50716));
    LocalMux I__11482 (
            .O(N__50727),
            .I(N__50713));
    Sp12to4 I__11481 (
            .O(N__50722),
            .I(N__50708));
    Span12Mux_s5_h I__11480 (
            .O(N__50719),
            .I(N__50708));
    Span4Mux_v I__11479 (
            .O(N__50716),
            .I(N__50703));
    Span4Mux_h I__11478 (
            .O(N__50713),
            .I(N__50703));
    Odrv12 I__11477 (
            .O(N__50708),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    Odrv4 I__11476 (
            .O(N__50703),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_31 ));
    InMux I__11475 (
            .O(N__50698),
            .I(N__50695));
    LocalMux I__11474 (
            .O(N__50695),
            .I(N__50691));
    InMux I__11473 (
            .O(N__50694),
            .I(N__50688));
    Span4Mux_v I__11472 (
            .O(N__50691),
            .I(N__50685));
    LocalMux I__11471 (
            .O(N__50688),
            .I(N__50682));
    Odrv4 I__11470 (
            .O(N__50685),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    Odrv4 I__11469 (
            .O(N__50682),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ));
    CascadeMux I__11468 (
            .O(N__50677),
            .I(N__50673));
    CascadeMux I__11467 (
            .O(N__50676),
            .I(N__50670));
    InMux I__11466 (
            .O(N__50673),
            .I(N__50667));
    InMux I__11465 (
            .O(N__50670),
            .I(N__50664));
    LocalMux I__11464 (
            .O(N__50667),
            .I(N__50661));
    LocalMux I__11463 (
            .O(N__50664),
            .I(N__50656));
    Span4Mux_v I__11462 (
            .O(N__50661),
            .I(N__50656));
    Span4Mux_h I__11461 (
            .O(N__50656),
            .I(N__50653));
    Odrv4 I__11460 (
            .O(N__50653),
            .I(\current_shift_inst.un38_control_input_5_0 ));
    CascadeMux I__11459 (
            .O(N__50650),
            .I(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ));
    InMux I__11458 (
            .O(N__50647),
            .I(N__50638));
    InMux I__11457 (
            .O(N__50646),
            .I(N__50638));
    InMux I__11456 (
            .O(N__50645),
            .I(N__50638));
    LocalMux I__11455 (
            .O(N__50638),
            .I(\current_shift_inst.PI_CTRL.N_31 ));
    InMux I__11454 (
            .O(N__50635),
            .I(N__50632));
    LocalMux I__11453 (
            .O(N__50632),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ));
    InMux I__11452 (
            .O(N__50629),
            .I(N__50626));
    LocalMux I__11451 (
            .O(N__50626),
            .I(N__50623));
    Odrv12 I__11450 (
            .O(N__50623),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ));
    InMux I__11449 (
            .O(N__50620),
            .I(N__50616));
    InMux I__11448 (
            .O(N__50619),
            .I(N__50613));
    LocalMux I__11447 (
            .O(N__50616),
            .I(N__50610));
    LocalMux I__11446 (
            .O(N__50613),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    Odrv4 I__11445 (
            .O(N__50610),
            .I(elapsed_time_ns_1_RNI47DN9_0_26));
    InMux I__11444 (
            .O(N__50605),
            .I(N__50602));
    LocalMux I__11443 (
            .O(N__50602),
            .I(N__50599));
    Odrv12 I__11442 (
            .O(N__50599),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ));
    InMux I__11441 (
            .O(N__50596),
            .I(N__50593));
    LocalMux I__11440 (
            .O(N__50593),
            .I(N__50589));
    CascadeMux I__11439 (
            .O(N__50592),
            .I(N__50586));
    Span4Mux_h I__11438 (
            .O(N__50589),
            .I(N__50583));
    InMux I__11437 (
            .O(N__50586),
            .I(N__50580));
    Odrv4 I__11436 (
            .O(N__50583),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    LocalMux I__11435 (
            .O(N__50580),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ));
    InMux I__11434 (
            .O(N__50575),
            .I(N__50571));
    InMux I__11433 (
            .O(N__50574),
            .I(N__50568));
    LocalMux I__11432 (
            .O(N__50571),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    LocalMux I__11431 (
            .O(N__50568),
            .I(elapsed_time_ns_1_RNI14DN9_0_23));
    InMux I__11430 (
            .O(N__50563),
            .I(N__50560));
    LocalMux I__11429 (
            .O(N__50560),
            .I(N__50556));
    InMux I__11428 (
            .O(N__50559),
            .I(N__50553));
    Odrv4 I__11427 (
            .O(N__50556),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    LocalMux I__11426 (
            .O(N__50553),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ));
    InMux I__11425 (
            .O(N__50548),
            .I(N__50541));
    InMux I__11424 (
            .O(N__50547),
            .I(N__50541));
    CascadeMux I__11423 (
            .O(N__50546),
            .I(N__50533));
    LocalMux I__11422 (
            .O(N__50541),
            .I(N__50519));
    InMux I__11421 (
            .O(N__50540),
            .I(N__50510));
    InMux I__11420 (
            .O(N__50539),
            .I(N__50510));
    InMux I__11419 (
            .O(N__50538),
            .I(N__50505));
    InMux I__11418 (
            .O(N__50537),
            .I(N__50505));
    InMux I__11417 (
            .O(N__50536),
            .I(N__50502));
    InMux I__11416 (
            .O(N__50533),
            .I(N__50493));
    InMux I__11415 (
            .O(N__50532),
            .I(N__50493));
    InMux I__11414 (
            .O(N__50531),
            .I(N__50493));
    InMux I__11413 (
            .O(N__50530),
            .I(N__50493));
    InMux I__11412 (
            .O(N__50529),
            .I(N__50490));
    CascadeMux I__11411 (
            .O(N__50528),
            .I(N__50487));
    InMux I__11410 (
            .O(N__50527),
            .I(N__50481));
    InMux I__11409 (
            .O(N__50526),
            .I(N__50474));
    InMux I__11408 (
            .O(N__50525),
            .I(N__50469));
    InMux I__11407 (
            .O(N__50524),
            .I(N__50469));
    InMux I__11406 (
            .O(N__50523),
            .I(N__50464));
    InMux I__11405 (
            .O(N__50522),
            .I(N__50464));
    Span4Mux_h I__11404 (
            .O(N__50519),
            .I(N__50461));
    InMux I__11403 (
            .O(N__50518),
            .I(N__50452));
    InMux I__11402 (
            .O(N__50517),
            .I(N__50452));
    InMux I__11401 (
            .O(N__50516),
            .I(N__50452));
    InMux I__11400 (
            .O(N__50515),
            .I(N__50452));
    LocalMux I__11399 (
            .O(N__50510),
            .I(N__50447));
    LocalMux I__11398 (
            .O(N__50505),
            .I(N__50447));
    LocalMux I__11397 (
            .O(N__50502),
            .I(N__50444));
    LocalMux I__11396 (
            .O(N__50493),
            .I(N__50439));
    LocalMux I__11395 (
            .O(N__50490),
            .I(N__50439));
    InMux I__11394 (
            .O(N__50487),
            .I(N__50430));
    InMux I__11393 (
            .O(N__50486),
            .I(N__50430));
    InMux I__11392 (
            .O(N__50485),
            .I(N__50430));
    InMux I__11391 (
            .O(N__50484),
            .I(N__50430));
    LocalMux I__11390 (
            .O(N__50481),
            .I(N__50427));
    InMux I__11389 (
            .O(N__50480),
            .I(N__50422));
    InMux I__11388 (
            .O(N__50479),
            .I(N__50422));
    InMux I__11387 (
            .O(N__50478),
            .I(N__50417));
    InMux I__11386 (
            .O(N__50477),
            .I(N__50417));
    LocalMux I__11385 (
            .O(N__50474),
            .I(N__50414));
    LocalMux I__11384 (
            .O(N__50469),
            .I(N__50407));
    LocalMux I__11383 (
            .O(N__50464),
            .I(N__50407));
    Span4Mux_v I__11382 (
            .O(N__50461),
            .I(N__50407));
    LocalMux I__11381 (
            .O(N__50452),
            .I(N__50398));
    Span4Mux_v I__11380 (
            .O(N__50447),
            .I(N__50398));
    Span4Mux_v I__11379 (
            .O(N__50444),
            .I(N__50398));
    Span4Mux_h I__11378 (
            .O(N__50439),
            .I(N__50398));
    LocalMux I__11377 (
            .O(N__50430),
            .I(N__50391));
    Span12Mux_s10_v I__11376 (
            .O(N__50427),
            .I(N__50391));
    LocalMux I__11375 (
            .O(N__50422),
            .I(N__50391));
    LocalMux I__11374 (
            .O(N__50417),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11373 (
            .O(N__50414),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11372 (
            .O(N__50407),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv4 I__11371 (
            .O(N__50398),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    Odrv12 I__11370 (
            .O(N__50391),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3 ));
    InMux I__11369 (
            .O(N__50380),
            .I(N__50376));
    InMux I__11368 (
            .O(N__50379),
            .I(N__50373));
    LocalMux I__11367 (
            .O(N__50376),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    LocalMux I__11366 (
            .O(N__50373),
            .I(elapsed_time_ns_1_RNI13CN9_0_14));
    IoInMux I__11365 (
            .O(N__50368),
            .I(N__50365));
    LocalMux I__11364 (
            .O(N__50365),
            .I(N__50362));
    Span12Mux_s4_v I__11363 (
            .O(N__50362),
            .I(N__50359));
    Span12Mux_v I__11362 (
            .O(N__50359),
            .I(N__50354));
    InMux I__11361 (
            .O(N__50358),
            .I(N__50349));
    InMux I__11360 (
            .O(N__50357),
            .I(N__50349));
    Odrv12 I__11359 (
            .O(N__50354),
            .I(s1_phy_c));
    LocalMux I__11358 (
            .O(N__50349),
            .I(s1_phy_c));
    InMux I__11357 (
            .O(N__50344),
            .I(N__50336));
    InMux I__11356 (
            .O(N__50343),
            .I(N__50336));
    InMux I__11355 (
            .O(N__50342),
            .I(N__50333));
    InMux I__11354 (
            .O(N__50341),
            .I(N__50329));
    LocalMux I__11353 (
            .O(N__50336),
            .I(N__50323));
    LocalMux I__11352 (
            .O(N__50333),
            .I(N__50323));
    InMux I__11351 (
            .O(N__50332),
            .I(N__50320));
    LocalMux I__11350 (
            .O(N__50329),
            .I(N__50317));
    InMux I__11349 (
            .O(N__50328),
            .I(N__50314));
    Span12Mux_s6_h I__11348 (
            .O(N__50323),
            .I(N__50311));
    LocalMux I__11347 (
            .O(N__50320),
            .I(state_3));
    Odrv4 I__11346 (
            .O(N__50317),
            .I(state_3));
    LocalMux I__11345 (
            .O(N__50314),
            .I(state_3));
    Odrv12 I__11344 (
            .O(N__50311),
            .I(state_3));
    InMux I__11343 (
            .O(N__50302),
            .I(N__50297));
    CascadeMux I__11342 (
            .O(N__50301),
            .I(N__50293));
    InMux I__11341 (
            .O(N__50300),
            .I(N__50290));
    LocalMux I__11340 (
            .O(N__50297),
            .I(N__50287));
    InMux I__11339 (
            .O(N__50296),
            .I(N__50282));
    InMux I__11338 (
            .O(N__50293),
            .I(N__50282));
    LocalMux I__11337 (
            .O(N__50290),
            .I(N__50279));
    Span4Mux_h I__11336 (
            .O(N__50287),
            .I(N__50276));
    LocalMux I__11335 (
            .O(N__50282),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__11334 (
            .O(N__50279),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    Odrv4 I__11333 (
            .O(N__50276),
            .I(\current_shift_inst.stop_timer_sZ0Z1 ));
    InMux I__11332 (
            .O(N__50269),
            .I(N__50263));
    InMux I__11331 (
            .O(N__50268),
            .I(N__50256));
    InMux I__11330 (
            .O(N__50267),
            .I(N__50256));
    InMux I__11329 (
            .O(N__50266),
            .I(N__50256));
    LocalMux I__11328 (
            .O(N__50263),
            .I(N__50253));
    LocalMux I__11327 (
            .O(N__50256),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    Odrv12 I__11326 (
            .O(N__50253),
            .I(\current_shift_inst.start_timer_sZ0Z1 ));
    InMux I__11325 (
            .O(N__50248),
            .I(N__50245));
    LocalMux I__11324 (
            .O(N__50245),
            .I(N__50240));
    InMux I__11323 (
            .O(N__50244),
            .I(N__50234));
    InMux I__11322 (
            .O(N__50243),
            .I(N__50234));
    Span4Mux_v I__11321 (
            .O(N__50240),
            .I(N__50231));
    InMux I__11320 (
            .O(N__50239),
            .I(N__50228));
    LocalMux I__11319 (
            .O(N__50234),
            .I(N__50223));
    Span4Mux_v I__11318 (
            .O(N__50231),
            .I(N__50223));
    LocalMux I__11317 (
            .O(N__50228),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    Odrv4 I__11316 (
            .O(N__50223),
            .I(\current_shift_inst.timer_s1.runningZ0 ));
    InMux I__11315 (
            .O(N__50218),
            .I(N__50214));
    InMux I__11314 (
            .O(N__50217),
            .I(N__50211));
    LocalMux I__11313 (
            .O(N__50214),
            .I(N__50208));
    LocalMux I__11312 (
            .O(N__50211),
            .I(N__50205));
    Span12Mux_s10_h I__11311 (
            .O(N__50208),
            .I(N__50202));
    Span4Mux_h I__11310 (
            .O(N__50205),
            .I(N__50199));
    Span12Mux_v I__11309 (
            .O(N__50202),
            .I(N__50196));
    Odrv4 I__11308 (
            .O(N__50199),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    Odrv12 I__11307 (
            .O(N__50196),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_0 ));
    CascadeMux I__11306 (
            .O(N__50191),
            .I(N__50188));
    InMux I__11305 (
            .O(N__50188),
            .I(N__50185));
    LocalMux I__11304 (
            .O(N__50185),
            .I(N__50182));
    Odrv4 I__11303 (
            .O(N__50182),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ));
    InMux I__11302 (
            .O(N__50179),
            .I(N__50176));
    LocalMux I__11301 (
            .O(N__50176),
            .I(N__50173));
    Span4Mux_v I__11300 (
            .O(N__50173),
            .I(N__50170));
    Odrv4 I__11299 (
            .O(N__50170),
            .I(\current_shift_inst.un38_control_input_0_s1_28 ));
    InMux I__11298 (
            .O(N__50167),
            .I(\current_shift_inst.un38_control_input_cry_27_s1 ));
    InMux I__11297 (
            .O(N__50164),
            .I(N__50161));
    LocalMux I__11296 (
            .O(N__50161),
            .I(N__50158));
    Odrv4 I__11295 (
            .O(N__50158),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ));
    InMux I__11294 (
            .O(N__50155),
            .I(N__50152));
    LocalMux I__11293 (
            .O(N__50152),
            .I(N__50149));
    Span4Mux_v I__11292 (
            .O(N__50149),
            .I(N__50146));
    Odrv4 I__11291 (
            .O(N__50146),
            .I(\current_shift_inst.un38_control_input_0_s1_29 ));
    InMux I__11290 (
            .O(N__50143),
            .I(\current_shift_inst.un38_control_input_cry_28_s1 ));
    CascadeMux I__11289 (
            .O(N__50140),
            .I(N__50137));
    InMux I__11288 (
            .O(N__50137),
            .I(N__50134));
    LocalMux I__11287 (
            .O(N__50134),
            .I(N__50131));
    Odrv4 I__11286 (
            .O(N__50131),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ));
    InMux I__11285 (
            .O(N__50128),
            .I(N__50125));
    LocalMux I__11284 (
            .O(N__50125),
            .I(N__50122));
    Span4Mux_h I__11283 (
            .O(N__50122),
            .I(N__50119));
    Odrv4 I__11282 (
            .O(N__50119),
            .I(\current_shift_inst.un38_control_input_0_s1_30 ));
    InMux I__11281 (
            .O(N__50116),
            .I(\current_shift_inst.un38_control_input_cry_29_s1 ));
    CascadeMux I__11280 (
            .O(N__50113),
            .I(N__50109));
    CascadeMux I__11279 (
            .O(N__50112),
            .I(N__50106));
    InMux I__11278 (
            .O(N__50109),
            .I(N__50101));
    InMux I__11277 (
            .O(N__50106),
            .I(N__50097));
    CascadeMux I__11276 (
            .O(N__50105),
            .I(N__50093));
    CascadeMux I__11275 (
            .O(N__50104),
            .I(N__50070));
    LocalMux I__11274 (
            .O(N__50101),
            .I(N__50063));
    CascadeMux I__11273 (
            .O(N__50100),
            .I(N__50058));
    LocalMux I__11272 (
            .O(N__50097),
            .I(N__50043));
    InMux I__11271 (
            .O(N__50096),
            .I(N__50038));
    InMux I__11270 (
            .O(N__50093),
            .I(N__50038));
    CascadeMux I__11269 (
            .O(N__50092),
            .I(N__50034));
    CascadeMux I__11268 (
            .O(N__50091),
            .I(N__50029));
    CascadeMux I__11267 (
            .O(N__50090),
            .I(N__50026));
    CascadeMux I__11266 (
            .O(N__50089),
            .I(N__50023));
    CascadeMux I__11265 (
            .O(N__50088),
            .I(N__50020));
    CascadeMux I__11264 (
            .O(N__50087),
            .I(N__50015));
    CascadeMux I__11263 (
            .O(N__50086),
            .I(N__50008));
    CascadeMux I__11262 (
            .O(N__50085),
            .I(N__49994));
    InMux I__11261 (
            .O(N__50084),
            .I(N__49979));
    InMux I__11260 (
            .O(N__50083),
            .I(N__49979));
    InMux I__11259 (
            .O(N__50082),
            .I(N__49979));
    InMux I__11258 (
            .O(N__50081),
            .I(N__49979));
    InMux I__11257 (
            .O(N__50080),
            .I(N__49979));
    InMux I__11256 (
            .O(N__50079),
            .I(N__49979));
    InMux I__11255 (
            .O(N__50078),
            .I(N__49979));
    InMux I__11254 (
            .O(N__50077),
            .I(N__49974));
    InMux I__11253 (
            .O(N__50076),
            .I(N__49974));
    InMux I__11252 (
            .O(N__50075),
            .I(N__49965));
    InMux I__11251 (
            .O(N__50074),
            .I(N__49965));
    InMux I__11250 (
            .O(N__50073),
            .I(N__49965));
    InMux I__11249 (
            .O(N__50070),
            .I(N__49965));
    CascadeMux I__11248 (
            .O(N__50069),
            .I(N__49960));
    CascadeMux I__11247 (
            .O(N__50068),
            .I(N__49956));
    CascadeMux I__11246 (
            .O(N__50067),
            .I(N__49952));
    InMux I__11245 (
            .O(N__50066),
            .I(N__49944));
    Span4Mux_v I__11244 (
            .O(N__50063),
            .I(N__49941));
    InMux I__11243 (
            .O(N__50062),
            .I(N__49930));
    InMux I__11242 (
            .O(N__50061),
            .I(N__49930));
    InMux I__11241 (
            .O(N__50058),
            .I(N__49930));
    InMux I__11240 (
            .O(N__50057),
            .I(N__49930));
    InMux I__11239 (
            .O(N__50056),
            .I(N__49930));
    InMux I__11238 (
            .O(N__50055),
            .I(N__49923));
    InMux I__11237 (
            .O(N__50054),
            .I(N__49923));
    InMux I__11236 (
            .O(N__50053),
            .I(N__49923));
    CascadeMux I__11235 (
            .O(N__50052),
            .I(N__49919));
    CascadeMux I__11234 (
            .O(N__50051),
            .I(N__49915));
    CascadeMux I__11233 (
            .O(N__50050),
            .I(N__49911));
    CascadeMux I__11232 (
            .O(N__50049),
            .I(N__49907));
    CascadeMux I__11231 (
            .O(N__50048),
            .I(N__49903));
    CascadeMux I__11230 (
            .O(N__50047),
            .I(N__49899));
    CascadeMux I__11229 (
            .O(N__50046),
            .I(N__49895));
    Span4Mux_v I__11228 (
            .O(N__50043),
            .I(N__49878));
    LocalMux I__11227 (
            .O(N__50038),
            .I(N__49874));
    InMux I__11226 (
            .O(N__50037),
            .I(N__49861));
    InMux I__11225 (
            .O(N__50034),
            .I(N__49861));
    InMux I__11224 (
            .O(N__50033),
            .I(N__49861));
    InMux I__11223 (
            .O(N__50032),
            .I(N__49861));
    InMux I__11222 (
            .O(N__50029),
            .I(N__49861));
    InMux I__11221 (
            .O(N__50026),
            .I(N__49861));
    InMux I__11220 (
            .O(N__50023),
            .I(N__49850));
    InMux I__11219 (
            .O(N__50020),
            .I(N__49850));
    InMux I__11218 (
            .O(N__50019),
            .I(N__49850));
    InMux I__11217 (
            .O(N__50018),
            .I(N__49850));
    InMux I__11216 (
            .O(N__50015),
            .I(N__49850));
    InMux I__11215 (
            .O(N__50014),
            .I(N__49833));
    InMux I__11214 (
            .O(N__50013),
            .I(N__49833));
    InMux I__11213 (
            .O(N__50012),
            .I(N__49833));
    InMux I__11212 (
            .O(N__50011),
            .I(N__49833));
    InMux I__11211 (
            .O(N__50008),
            .I(N__49833));
    InMux I__11210 (
            .O(N__50007),
            .I(N__49833));
    InMux I__11209 (
            .O(N__50006),
            .I(N__49833));
    InMux I__11208 (
            .O(N__50005),
            .I(N__49833));
    CascadeMux I__11207 (
            .O(N__50004),
            .I(N__49830));
    CascadeMux I__11206 (
            .O(N__50003),
            .I(N__49826));
    CascadeMux I__11205 (
            .O(N__50002),
            .I(N__49821));
    CascadeMux I__11204 (
            .O(N__50001),
            .I(N__49818));
    CascadeMux I__11203 (
            .O(N__50000),
            .I(N__49814));
    InMux I__11202 (
            .O(N__49999),
            .I(N__49805));
    InMux I__11201 (
            .O(N__49998),
            .I(N__49805));
    InMux I__11200 (
            .O(N__49997),
            .I(N__49805));
    InMux I__11199 (
            .O(N__49994),
            .I(N__49805));
    LocalMux I__11198 (
            .O(N__49979),
            .I(N__49800));
    LocalMux I__11197 (
            .O(N__49974),
            .I(N__49800));
    LocalMux I__11196 (
            .O(N__49965),
            .I(N__49797));
    InMux I__11195 (
            .O(N__49964),
            .I(N__49780));
    InMux I__11194 (
            .O(N__49963),
            .I(N__49780));
    InMux I__11193 (
            .O(N__49960),
            .I(N__49780));
    InMux I__11192 (
            .O(N__49959),
            .I(N__49780));
    InMux I__11191 (
            .O(N__49956),
            .I(N__49780));
    InMux I__11190 (
            .O(N__49955),
            .I(N__49780));
    InMux I__11189 (
            .O(N__49952),
            .I(N__49780));
    InMux I__11188 (
            .O(N__49951),
            .I(N__49780));
    CascadeMux I__11187 (
            .O(N__49950),
            .I(N__49776));
    CascadeMux I__11186 (
            .O(N__49949),
            .I(N__49772));
    CascadeMux I__11185 (
            .O(N__49948),
            .I(N__49768));
    CascadeMux I__11184 (
            .O(N__49947),
            .I(N__49764));
    LocalMux I__11183 (
            .O(N__49944),
            .I(N__49761));
    Span4Mux_h I__11182 (
            .O(N__49941),
            .I(N__49754));
    LocalMux I__11181 (
            .O(N__49930),
            .I(N__49754));
    LocalMux I__11180 (
            .O(N__49923),
            .I(N__49754));
    InMux I__11179 (
            .O(N__49922),
            .I(N__49739));
    InMux I__11178 (
            .O(N__49919),
            .I(N__49739));
    InMux I__11177 (
            .O(N__49918),
            .I(N__49739));
    InMux I__11176 (
            .O(N__49915),
            .I(N__49739));
    InMux I__11175 (
            .O(N__49914),
            .I(N__49739));
    InMux I__11174 (
            .O(N__49911),
            .I(N__49739));
    InMux I__11173 (
            .O(N__49910),
            .I(N__49739));
    InMux I__11172 (
            .O(N__49907),
            .I(N__49722));
    InMux I__11171 (
            .O(N__49906),
            .I(N__49722));
    InMux I__11170 (
            .O(N__49903),
            .I(N__49722));
    InMux I__11169 (
            .O(N__49902),
            .I(N__49722));
    InMux I__11168 (
            .O(N__49899),
            .I(N__49722));
    InMux I__11167 (
            .O(N__49898),
            .I(N__49722));
    InMux I__11166 (
            .O(N__49895),
            .I(N__49722));
    InMux I__11165 (
            .O(N__49894),
            .I(N__49722));
    CascadeMux I__11164 (
            .O(N__49893),
            .I(N__49719));
    CascadeMux I__11163 (
            .O(N__49892),
            .I(N__49715));
    CascadeMux I__11162 (
            .O(N__49891),
            .I(N__49711));
    CascadeMux I__11161 (
            .O(N__49890),
            .I(N__49707));
    CascadeMux I__11160 (
            .O(N__49889),
            .I(N__49703));
    CascadeMux I__11159 (
            .O(N__49888),
            .I(N__49699));
    CascadeMux I__11158 (
            .O(N__49887),
            .I(N__49695));
    CascadeMux I__11157 (
            .O(N__49886),
            .I(N__49691));
    CascadeMux I__11156 (
            .O(N__49885),
            .I(N__49685));
    CascadeMux I__11155 (
            .O(N__49884),
            .I(N__49681));
    CascadeMux I__11154 (
            .O(N__49883),
            .I(N__49676));
    CascadeMux I__11153 (
            .O(N__49882),
            .I(N__49672));
    CascadeMux I__11152 (
            .O(N__49881),
            .I(N__49668));
    Span4Mux_v I__11151 (
            .O(N__49878),
            .I(N__49665));
    InMux I__11150 (
            .O(N__49877),
            .I(N__49662));
    Span4Mux_v I__11149 (
            .O(N__49874),
            .I(N__49653));
    LocalMux I__11148 (
            .O(N__49861),
            .I(N__49653));
    LocalMux I__11147 (
            .O(N__49850),
            .I(N__49653));
    LocalMux I__11146 (
            .O(N__49833),
            .I(N__49653));
    InMux I__11145 (
            .O(N__49830),
            .I(N__49650));
    InMux I__11144 (
            .O(N__49829),
            .I(N__49633));
    InMux I__11143 (
            .O(N__49826),
            .I(N__49633));
    InMux I__11142 (
            .O(N__49825),
            .I(N__49633));
    InMux I__11141 (
            .O(N__49824),
            .I(N__49633));
    InMux I__11140 (
            .O(N__49821),
            .I(N__49633));
    InMux I__11139 (
            .O(N__49818),
            .I(N__49633));
    InMux I__11138 (
            .O(N__49817),
            .I(N__49633));
    InMux I__11137 (
            .O(N__49814),
            .I(N__49633));
    LocalMux I__11136 (
            .O(N__49805),
            .I(N__49628));
    Span4Mux_v I__11135 (
            .O(N__49800),
            .I(N__49628));
    Span4Mux_v I__11134 (
            .O(N__49797),
            .I(N__49623));
    LocalMux I__11133 (
            .O(N__49780),
            .I(N__49623));
    InMux I__11132 (
            .O(N__49779),
            .I(N__49606));
    InMux I__11131 (
            .O(N__49776),
            .I(N__49606));
    InMux I__11130 (
            .O(N__49775),
            .I(N__49606));
    InMux I__11129 (
            .O(N__49772),
            .I(N__49606));
    InMux I__11128 (
            .O(N__49771),
            .I(N__49606));
    InMux I__11127 (
            .O(N__49768),
            .I(N__49606));
    InMux I__11126 (
            .O(N__49767),
            .I(N__49606));
    InMux I__11125 (
            .O(N__49764),
            .I(N__49606));
    Sp12to4 I__11124 (
            .O(N__49761),
            .I(N__49597));
    Sp12to4 I__11123 (
            .O(N__49754),
            .I(N__49597));
    LocalMux I__11122 (
            .O(N__49739),
            .I(N__49597));
    LocalMux I__11121 (
            .O(N__49722),
            .I(N__49597));
    InMux I__11120 (
            .O(N__49719),
            .I(N__49580));
    InMux I__11119 (
            .O(N__49718),
            .I(N__49580));
    InMux I__11118 (
            .O(N__49715),
            .I(N__49580));
    InMux I__11117 (
            .O(N__49714),
            .I(N__49580));
    InMux I__11116 (
            .O(N__49711),
            .I(N__49580));
    InMux I__11115 (
            .O(N__49710),
            .I(N__49580));
    InMux I__11114 (
            .O(N__49707),
            .I(N__49580));
    InMux I__11113 (
            .O(N__49706),
            .I(N__49580));
    InMux I__11112 (
            .O(N__49703),
            .I(N__49563));
    InMux I__11111 (
            .O(N__49702),
            .I(N__49563));
    InMux I__11110 (
            .O(N__49699),
            .I(N__49563));
    InMux I__11109 (
            .O(N__49698),
            .I(N__49563));
    InMux I__11108 (
            .O(N__49695),
            .I(N__49563));
    InMux I__11107 (
            .O(N__49694),
            .I(N__49563));
    InMux I__11106 (
            .O(N__49691),
            .I(N__49563));
    InMux I__11105 (
            .O(N__49690),
            .I(N__49563));
    InMux I__11104 (
            .O(N__49689),
            .I(N__49560));
    InMux I__11103 (
            .O(N__49688),
            .I(N__49549));
    InMux I__11102 (
            .O(N__49685),
            .I(N__49549));
    InMux I__11101 (
            .O(N__49684),
            .I(N__49549));
    InMux I__11100 (
            .O(N__49681),
            .I(N__49549));
    InMux I__11099 (
            .O(N__49680),
            .I(N__49549));
    InMux I__11098 (
            .O(N__49679),
            .I(N__49536));
    InMux I__11097 (
            .O(N__49676),
            .I(N__49536));
    InMux I__11096 (
            .O(N__49675),
            .I(N__49536));
    InMux I__11095 (
            .O(N__49672),
            .I(N__49536));
    InMux I__11094 (
            .O(N__49671),
            .I(N__49536));
    InMux I__11093 (
            .O(N__49668),
            .I(N__49536));
    Odrv4 I__11092 (
            .O(N__49665),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11091 (
            .O(N__49662),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11090 (
            .O(N__49653),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11089 (
            .O(N__49650),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11088 (
            .O(N__49633),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11087 (
            .O(N__49628),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv4 I__11086 (
            .O(N__49623),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11085 (
            .O(N__49606),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    Odrv12 I__11084 (
            .O(N__49597),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11083 (
            .O(N__49580),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11082 (
            .O(N__49563),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11081 (
            .O(N__49560),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11080 (
            .O(N__49549),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    LocalMux I__11079 (
            .O(N__49536),
            .I(\current_shift_inst.un38_control_input_5_2 ));
    InMux I__11078 (
            .O(N__49507),
            .I(N__49483));
    InMux I__11077 (
            .O(N__49506),
            .I(N__49483));
    InMux I__11076 (
            .O(N__49505),
            .I(N__49483));
    InMux I__11075 (
            .O(N__49504),
            .I(N__49483));
    InMux I__11074 (
            .O(N__49503),
            .I(N__49483));
    InMux I__11073 (
            .O(N__49502),
            .I(N__49480));
    InMux I__11072 (
            .O(N__49501),
            .I(N__49473));
    InMux I__11071 (
            .O(N__49500),
            .I(N__49473));
    InMux I__11070 (
            .O(N__49499),
            .I(N__49473));
    InMux I__11069 (
            .O(N__49498),
            .I(N__49460));
    InMux I__11068 (
            .O(N__49497),
            .I(N__49460));
    InMux I__11067 (
            .O(N__49496),
            .I(N__49457));
    InMux I__11066 (
            .O(N__49495),
            .I(N__49454));
    InMux I__11065 (
            .O(N__49494),
            .I(N__49449));
    LocalMux I__11064 (
            .O(N__49483),
            .I(N__49439));
    LocalMux I__11063 (
            .O(N__49480),
            .I(N__49439));
    LocalMux I__11062 (
            .O(N__49473),
            .I(N__49439));
    InMux I__11061 (
            .O(N__49472),
            .I(N__49422));
    InMux I__11060 (
            .O(N__49471),
            .I(N__49422));
    InMux I__11059 (
            .O(N__49470),
            .I(N__49422));
    InMux I__11058 (
            .O(N__49469),
            .I(N__49422));
    InMux I__11057 (
            .O(N__49468),
            .I(N__49422));
    InMux I__11056 (
            .O(N__49467),
            .I(N__49422));
    InMux I__11055 (
            .O(N__49466),
            .I(N__49422));
    InMux I__11054 (
            .O(N__49465),
            .I(N__49422));
    LocalMux I__11053 (
            .O(N__49460),
            .I(N__49419));
    LocalMux I__11052 (
            .O(N__49457),
            .I(N__49416));
    LocalMux I__11051 (
            .O(N__49454),
            .I(N__49405));
    InMux I__11050 (
            .O(N__49453),
            .I(N__49400));
    InMux I__11049 (
            .O(N__49452),
            .I(N__49400));
    LocalMux I__11048 (
            .O(N__49449),
            .I(N__49397));
    InMux I__11047 (
            .O(N__49448),
            .I(N__49390));
    InMux I__11046 (
            .O(N__49447),
            .I(N__49390));
    InMux I__11045 (
            .O(N__49446),
            .I(N__49390));
    Span4Mux_v I__11044 (
            .O(N__49439),
            .I(N__49381));
    LocalMux I__11043 (
            .O(N__49422),
            .I(N__49381));
    Span4Mux_v I__11042 (
            .O(N__49419),
            .I(N__49381));
    Span4Mux_h I__11041 (
            .O(N__49416),
            .I(N__49381));
    InMux I__11040 (
            .O(N__49415),
            .I(N__49355));
    InMux I__11039 (
            .O(N__49414),
            .I(N__49355));
    InMux I__11038 (
            .O(N__49413),
            .I(N__49334));
    InMux I__11037 (
            .O(N__49412),
            .I(N__49334));
    InMux I__11036 (
            .O(N__49411),
            .I(N__49334));
    InMux I__11035 (
            .O(N__49410),
            .I(N__49334));
    InMux I__11034 (
            .O(N__49409),
            .I(N__49334));
    CascadeMux I__11033 (
            .O(N__49408),
            .I(N__49328));
    Span4Mux_h I__11032 (
            .O(N__49405),
            .I(N__49321));
    LocalMux I__11031 (
            .O(N__49400),
            .I(N__49321));
    Span4Mux_v I__11030 (
            .O(N__49397),
            .I(N__49316));
    LocalMux I__11029 (
            .O(N__49390),
            .I(N__49316));
    Span4Mux_v I__11028 (
            .O(N__49381),
            .I(N__49313));
    InMux I__11027 (
            .O(N__49380),
            .I(N__49304));
    InMux I__11026 (
            .O(N__49379),
            .I(N__49304));
    InMux I__11025 (
            .O(N__49378),
            .I(N__49304));
    InMux I__11024 (
            .O(N__49377),
            .I(N__49304));
    InMux I__11023 (
            .O(N__49376),
            .I(N__49291));
    InMux I__11022 (
            .O(N__49375),
            .I(N__49291));
    InMux I__11021 (
            .O(N__49374),
            .I(N__49291));
    InMux I__11020 (
            .O(N__49373),
            .I(N__49291));
    InMux I__11019 (
            .O(N__49372),
            .I(N__49291));
    InMux I__11018 (
            .O(N__49371),
            .I(N__49291));
    InMux I__11017 (
            .O(N__49370),
            .I(N__49274));
    InMux I__11016 (
            .O(N__49369),
            .I(N__49274));
    InMux I__11015 (
            .O(N__49368),
            .I(N__49274));
    InMux I__11014 (
            .O(N__49367),
            .I(N__49274));
    InMux I__11013 (
            .O(N__49366),
            .I(N__49274));
    InMux I__11012 (
            .O(N__49365),
            .I(N__49274));
    InMux I__11011 (
            .O(N__49364),
            .I(N__49274));
    InMux I__11010 (
            .O(N__49363),
            .I(N__49274));
    InMux I__11009 (
            .O(N__49362),
            .I(N__49267));
    InMux I__11008 (
            .O(N__49361),
            .I(N__49267));
    InMux I__11007 (
            .O(N__49360),
            .I(N__49267));
    LocalMux I__11006 (
            .O(N__49355),
            .I(N__49264));
    InMux I__11005 (
            .O(N__49354),
            .I(N__49249));
    InMux I__11004 (
            .O(N__49353),
            .I(N__49249));
    InMux I__11003 (
            .O(N__49352),
            .I(N__49249));
    InMux I__11002 (
            .O(N__49351),
            .I(N__49249));
    InMux I__11001 (
            .O(N__49350),
            .I(N__49249));
    InMux I__11000 (
            .O(N__49349),
            .I(N__49249));
    InMux I__10999 (
            .O(N__49348),
            .I(N__49249));
    InMux I__10998 (
            .O(N__49347),
            .I(N__49242));
    InMux I__10997 (
            .O(N__49346),
            .I(N__49242));
    InMux I__10996 (
            .O(N__49345),
            .I(N__49242));
    LocalMux I__10995 (
            .O(N__49334),
            .I(N__49239));
    InMux I__10994 (
            .O(N__49333),
            .I(N__49226));
    InMux I__10993 (
            .O(N__49332),
            .I(N__49226));
    InMux I__10992 (
            .O(N__49331),
            .I(N__49226));
    InMux I__10991 (
            .O(N__49328),
            .I(N__49226));
    InMux I__10990 (
            .O(N__49327),
            .I(N__49226));
    InMux I__10989 (
            .O(N__49326),
            .I(N__49226));
    Span4Mux_v I__10988 (
            .O(N__49321),
            .I(N__49221));
    Span4Mux_h I__10987 (
            .O(N__49316),
            .I(N__49221));
    Odrv4 I__10986 (
            .O(N__49313),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10985 (
            .O(N__49304),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10984 (
            .O(N__49291),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10983 (
            .O(N__49274),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10982 (
            .O(N__49267),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10981 (
            .O(N__49264),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10980 (
            .O(N__49249),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10979 (
            .O(N__49242),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10978 (
            .O(N__49239),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    LocalMux I__10977 (
            .O(N__49226),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    Odrv4 I__10976 (
            .O(N__49221),
            .I(\current_shift_inst.elapsed_time_ns_s1_31 ));
    InMux I__10975 (
            .O(N__49198),
            .I(\current_shift_inst.un38_control_input_cry_30_s1 ));
    InMux I__10974 (
            .O(N__49195),
            .I(N__49192));
    LocalMux I__10973 (
            .O(N__49192),
            .I(\current_shift_inst.un38_control_input_0_s1_31 ));
    InMux I__10972 (
            .O(N__49189),
            .I(N__49186));
    LocalMux I__10971 (
            .O(N__49186),
            .I(\current_shift_inst.un38_control_input_0_s0_26 ));
    InMux I__10970 (
            .O(N__49183),
            .I(N__49180));
    LocalMux I__10969 (
            .O(N__49180),
            .I(\current_shift_inst.un38_control_input_0_s1_26 ));
    CascadeMux I__10968 (
            .O(N__49177),
            .I(N__49174));
    InMux I__10967 (
            .O(N__49174),
            .I(N__49170));
    InMux I__10966 (
            .O(N__49173),
            .I(N__49167));
    LocalMux I__10965 (
            .O(N__49170),
            .I(N__49150));
    LocalMux I__10964 (
            .O(N__49167),
            .I(N__49150));
    InMux I__10963 (
            .O(N__49166),
            .I(N__49145));
    InMux I__10962 (
            .O(N__49165),
            .I(N__49145));
    InMux I__10961 (
            .O(N__49164),
            .I(N__49142));
    InMux I__10960 (
            .O(N__49163),
            .I(N__49137));
    InMux I__10959 (
            .O(N__49162),
            .I(N__49137));
    InMux I__10958 (
            .O(N__49161),
            .I(N__49122));
    InMux I__10957 (
            .O(N__49160),
            .I(N__49122));
    InMux I__10956 (
            .O(N__49159),
            .I(N__49122));
    InMux I__10955 (
            .O(N__49158),
            .I(N__49122));
    InMux I__10954 (
            .O(N__49157),
            .I(N__49122));
    InMux I__10953 (
            .O(N__49156),
            .I(N__49122));
    InMux I__10952 (
            .O(N__49155),
            .I(N__49122));
    Span4Mux_h I__10951 (
            .O(N__49150),
            .I(N__49101));
    LocalMux I__10950 (
            .O(N__49145),
            .I(N__49098));
    LocalMux I__10949 (
            .O(N__49142),
            .I(N__49091));
    LocalMux I__10948 (
            .O(N__49137),
            .I(N__49091));
    LocalMux I__10947 (
            .O(N__49122),
            .I(N__49091));
    InMux I__10946 (
            .O(N__49121),
            .I(N__49080));
    InMux I__10945 (
            .O(N__49120),
            .I(N__49080));
    InMux I__10944 (
            .O(N__49119),
            .I(N__49080));
    InMux I__10943 (
            .O(N__49118),
            .I(N__49080));
    InMux I__10942 (
            .O(N__49117),
            .I(N__49080));
    InMux I__10941 (
            .O(N__49116),
            .I(N__49063));
    InMux I__10940 (
            .O(N__49115),
            .I(N__49063));
    InMux I__10939 (
            .O(N__49114),
            .I(N__49063));
    InMux I__10938 (
            .O(N__49113),
            .I(N__49063));
    InMux I__10937 (
            .O(N__49112),
            .I(N__49063));
    InMux I__10936 (
            .O(N__49111),
            .I(N__49063));
    InMux I__10935 (
            .O(N__49110),
            .I(N__49063));
    InMux I__10934 (
            .O(N__49109),
            .I(N__49063));
    InMux I__10933 (
            .O(N__49108),
            .I(N__49052));
    InMux I__10932 (
            .O(N__49107),
            .I(N__49052));
    InMux I__10931 (
            .O(N__49106),
            .I(N__49052));
    InMux I__10930 (
            .O(N__49105),
            .I(N__49052));
    InMux I__10929 (
            .O(N__49104),
            .I(N__49052));
    Odrv4 I__10928 (
            .O(N__49101),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10927 (
            .O(N__49098),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    Odrv4 I__10926 (
            .O(N__49091),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10925 (
            .O(N__49080),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10924 (
            .O(N__49063),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    LocalMux I__10923 (
            .O(N__49052),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ));
    InMux I__10922 (
            .O(N__49039),
            .I(N__49036));
    LocalMux I__10921 (
            .O(N__49036),
            .I(N__49033));
    Odrv12 I__10920 (
            .O(N__49033),
            .I(\current_shift_inst.control_input_axb_23 ));
    InMux I__10919 (
            .O(N__49030),
            .I(N__49027));
    LocalMux I__10918 (
            .O(N__49027),
            .I(N__49024));
    Span4Mux_v I__10917 (
            .O(N__49024),
            .I(N__49020));
    InMux I__10916 (
            .O(N__49023),
            .I(N__49017));
    Odrv4 I__10915 (
            .O(N__49020),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    LocalMux I__10914 (
            .O(N__49017),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ));
    InMux I__10913 (
            .O(N__49012),
            .I(N__49009));
    LocalMux I__10912 (
            .O(N__49009),
            .I(elapsed_time_ns_1_RNI02CN9_0_13));
    CascadeMux I__10911 (
            .O(N__49006),
            .I(elapsed_time_ns_1_RNI02CN9_0_13_cascade_));
    InMux I__10910 (
            .O(N__49003),
            .I(N__49000));
    LocalMux I__10909 (
            .O(N__49000),
            .I(N__48997));
    Odrv12 I__10908 (
            .O(N__48997),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ));
    InMux I__10907 (
            .O(N__48994),
            .I(N__48991));
    LocalMux I__10906 (
            .O(N__48991),
            .I(N__48988));
    Span12Mux_s9_v I__10905 (
            .O(N__48988),
            .I(N__48985));
    Odrv12 I__10904 (
            .O(N__48985),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ));
    InMux I__10903 (
            .O(N__48982),
            .I(N__48979));
    LocalMux I__10902 (
            .O(N__48979),
            .I(N__48976));
    Span4Mux_h I__10901 (
            .O(N__48976),
            .I(N__48973));
    Odrv4 I__10900 (
            .O(N__48973),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ));
    InMux I__10899 (
            .O(N__48970),
            .I(N__48967));
    LocalMux I__10898 (
            .O(N__48967),
            .I(N__48964));
    Span4Mux_h I__10897 (
            .O(N__48964),
            .I(N__48961));
    Odrv4 I__10896 (
            .O(N__48961),
            .I(\current_shift_inst.un38_control_input_0_s1_20 ));
    InMux I__10895 (
            .O(N__48958),
            .I(\current_shift_inst.un38_control_input_cry_19_s1 ));
    CascadeMux I__10894 (
            .O(N__48955),
            .I(N__48952));
    InMux I__10893 (
            .O(N__48952),
            .I(N__48949));
    LocalMux I__10892 (
            .O(N__48949),
            .I(N__48946));
    Odrv4 I__10891 (
            .O(N__48946),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ));
    InMux I__10890 (
            .O(N__48943),
            .I(N__48940));
    LocalMux I__10889 (
            .O(N__48940),
            .I(N__48937));
    Span4Mux_h I__10888 (
            .O(N__48937),
            .I(N__48934));
    Odrv4 I__10887 (
            .O(N__48934),
            .I(\current_shift_inst.un38_control_input_0_s1_21 ));
    InMux I__10886 (
            .O(N__48931),
            .I(\current_shift_inst.un38_control_input_cry_20_s1 ));
    InMux I__10885 (
            .O(N__48928),
            .I(N__48925));
    LocalMux I__10884 (
            .O(N__48925),
            .I(N__48922));
    Odrv12 I__10883 (
            .O(N__48922),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ));
    InMux I__10882 (
            .O(N__48919),
            .I(N__48916));
    LocalMux I__10881 (
            .O(N__48916),
            .I(N__48913));
    Span4Mux_h I__10880 (
            .O(N__48913),
            .I(N__48910));
    Odrv4 I__10879 (
            .O(N__48910),
            .I(\current_shift_inst.un38_control_input_0_s1_22 ));
    InMux I__10878 (
            .O(N__48907),
            .I(\current_shift_inst.un38_control_input_cry_21_s1 ));
    CascadeMux I__10877 (
            .O(N__48904),
            .I(N__48901));
    InMux I__10876 (
            .O(N__48901),
            .I(N__48898));
    LocalMux I__10875 (
            .O(N__48898),
            .I(N__48895));
    Odrv12 I__10874 (
            .O(N__48895),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ));
    InMux I__10873 (
            .O(N__48892),
            .I(N__48889));
    LocalMux I__10872 (
            .O(N__48889),
            .I(N__48886));
    Span4Mux_h I__10871 (
            .O(N__48886),
            .I(N__48883));
    Odrv4 I__10870 (
            .O(N__48883),
            .I(\current_shift_inst.un38_control_input_0_s1_23 ));
    InMux I__10869 (
            .O(N__48880),
            .I(\current_shift_inst.un38_control_input_cry_22_s1 ));
    CascadeMux I__10868 (
            .O(N__48877),
            .I(N__48874));
    InMux I__10867 (
            .O(N__48874),
            .I(N__48871));
    LocalMux I__10866 (
            .O(N__48871),
            .I(N__48868));
    Odrv4 I__10865 (
            .O(N__48868),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ));
    InMux I__10864 (
            .O(N__48865),
            .I(N__48862));
    LocalMux I__10863 (
            .O(N__48862),
            .I(N__48859));
    Span4Mux_h I__10862 (
            .O(N__48859),
            .I(N__48856));
    Odrv4 I__10861 (
            .O(N__48856),
            .I(\current_shift_inst.un38_control_input_0_s1_24 ));
    InMux I__10860 (
            .O(N__48853),
            .I(bfn_18_20_0_));
    InMux I__10859 (
            .O(N__48850),
            .I(N__48847));
    LocalMux I__10858 (
            .O(N__48847),
            .I(N__48844));
    Odrv4 I__10857 (
            .O(N__48844),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ));
    InMux I__10856 (
            .O(N__48841),
            .I(N__48838));
    LocalMux I__10855 (
            .O(N__48838),
            .I(N__48835));
    Span4Mux_h I__10854 (
            .O(N__48835),
            .I(N__48832));
    Odrv4 I__10853 (
            .O(N__48832),
            .I(\current_shift_inst.un38_control_input_0_s1_25 ));
    InMux I__10852 (
            .O(N__48829),
            .I(\current_shift_inst.un38_control_input_cry_24_s1 ));
    CascadeMux I__10851 (
            .O(N__48826),
            .I(N__48823));
    InMux I__10850 (
            .O(N__48823),
            .I(N__48820));
    LocalMux I__10849 (
            .O(N__48820),
            .I(N__48817));
    Odrv4 I__10848 (
            .O(N__48817),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ));
    InMux I__10847 (
            .O(N__48814),
            .I(\current_shift_inst.un38_control_input_cry_25_s1 ));
    InMux I__10846 (
            .O(N__48811),
            .I(N__48808));
    LocalMux I__10845 (
            .O(N__48808),
            .I(N__48805));
    Span4Mux_v I__10844 (
            .O(N__48805),
            .I(N__48802));
    Odrv4 I__10843 (
            .O(N__48802),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ));
    InMux I__10842 (
            .O(N__48799),
            .I(N__48796));
    LocalMux I__10841 (
            .O(N__48796),
            .I(N__48793));
    Odrv12 I__10840 (
            .O(N__48793),
            .I(\current_shift_inst.un38_control_input_0_s1_27 ));
    InMux I__10839 (
            .O(N__48790),
            .I(\current_shift_inst.un38_control_input_cry_26_s1 ));
    CascadeMux I__10838 (
            .O(N__48787),
            .I(N__48784));
    InMux I__10837 (
            .O(N__48784),
            .I(N__48781));
    LocalMux I__10836 (
            .O(N__48781),
            .I(N__48778));
    Span4Mux_v I__10835 (
            .O(N__48778),
            .I(N__48775));
    Odrv4 I__10834 (
            .O(N__48775),
            .I(\current_shift_inst.un38_control_input_0_s1_12 ));
    InMux I__10833 (
            .O(N__48772),
            .I(\current_shift_inst.un38_control_input_cry_11_s1 ));
    InMux I__10832 (
            .O(N__48769),
            .I(N__48766));
    LocalMux I__10831 (
            .O(N__48766),
            .I(N__48763));
    Odrv4 I__10830 (
            .O(N__48763),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ));
    InMux I__10829 (
            .O(N__48760),
            .I(N__48757));
    LocalMux I__10828 (
            .O(N__48757),
            .I(N__48754));
    Span4Mux_v I__10827 (
            .O(N__48754),
            .I(N__48751));
    Odrv4 I__10826 (
            .O(N__48751),
            .I(\current_shift_inst.un38_control_input_0_s1_13 ));
    InMux I__10825 (
            .O(N__48748),
            .I(\current_shift_inst.un38_control_input_cry_12_s1 ));
    CascadeMux I__10824 (
            .O(N__48745),
            .I(N__48742));
    InMux I__10823 (
            .O(N__48742),
            .I(N__48739));
    LocalMux I__10822 (
            .O(N__48739),
            .I(N__48736));
    Span4Mux_v I__10821 (
            .O(N__48736),
            .I(N__48733));
    Odrv4 I__10820 (
            .O(N__48733),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ));
    InMux I__10819 (
            .O(N__48730),
            .I(N__48727));
    LocalMux I__10818 (
            .O(N__48727),
            .I(N__48724));
    Span4Mux_h I__10817 (
            .O(N__48724),
            .I(N__48721));
    Odrv4 I__10816 (
            .O(N__48721),
            .I(\current_shift_inst.un38_control_input_0_s1_14 ));
    InMux I__10815 (
            .O(N__48718),
            .I(\current_shift_inst.un38_control_input_cry_13_s1 ));
    InMux I__10814 (
            .O(N__48715),
            .I(N__48712));
    LocalMux I__10813 (
            .O(N__48712),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ));
    InMux I__10812 (
            .O(N__48709),
            .I(N__48706));
    LocalMux I__10811 (
            .O(N__48706),
            .I(N__48703));
    Span4Mux_h I__10810 (
            .O(N__48703),
            .I(N__48700));
    Odrv4 I__10809 (
            .O(N__48700),
            .I(\current_shift_inst.un38_control_input_0_s1_15 ));
    InMux I__10808 (
            .O(N__48697),
            .I(\current_shift_inst.un38_control_input_cry_14_s1 ));
    InMux I__10807 (
            .O(N__48694),
            .I(N__48691));
    LocalMux I__10806 (
            .O(N__48691),
            .I(N__48688));
    Odrv12 I__10805 (
            .O(N__48688),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ));
    InMux I__10804 (
            .O(N__48685),
            .I(N__48682));
    LocalMux I__10803 (
            .O(N__48682),
            .I(N__48679));
    Span4Mux_h I__10802 (
            .O(N__48679),
            .I(N__48676));
    Odrv4 I__10801 (
            .O(N__48676),
            .I(\current_shift_inst.un38_control_input_0_s1_16 ));
    InMux I__10800 (
            .O(N__48673),
            .I(bfn_18_19_0_));
    CascadeMux I__10799 (
            .O(N__48670),
            .I(N__48667));
    InMux I__10798 (
            .O(N__48667),
            .I(N__48664));
    LocalMux I__10797 (
            .O(N__48664),
            .I(N__48661));
    Odrv12 I__10796 (
            .O(N__48661),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ));
    InMux I__10795 (
            .O(N__48658),
            .I(N__48655));
    LocalMux I__10794 (
            .O(N__48655),
            .I(N__48652));
    Span4Mux_h I__10793 (
            .O(N__48652),
            .I(N__48649));
    Odrv4 I__10792 (
            .O(N__48649),
            .I(\current_shift_inst.un38_control_input_0_s1_17 ));
    InMux I__10791 (
            .O(N__48646),
            .I(\current_shift_inst.un38_control_input_cry_16_s1 ));
    InMux I__10790 (
            .O(N__48643),
            .I(N__48640));
    LocalMux I__10789 (
            .O(N__48640),
            .I(N__48637));
    Odrv12 I__10788 (
            .O(N__48637),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ));
    InMux I__10787 (
            .O(N__48634),
            .I(N__48631));
    LocalMux I__10786 (
            .O(N__48631),
            .I(N__48628));
    Span4Mux_h I__10785 (
            .O(N__48628),
            .I(N__48625));
    Odrv4 I__10784 (
            .O(N__48625),
            .I(\current_shift_inst.un38_control_input_0_s1_18 ));
    InMux I__10783 (
            .O(N__48622),
            .I(\current_shift_inst.un38_control_input_cry_17_s1 ));
    CascadeMux I__10782 (
            .O(N__48619),
            .I(N__48616));
    InMux I__10781 (
            .O(N__48616),
            .I(N__48613));
    LocalMux I__10780 (
            .O(N__48613),
            .I(N__48610));
    Span4Mux_v I__10779 (
            .O(N__48610),
            .I(N__48607));
    Odrv4 I__10778 (
            .O(N__48607),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ));
    InMux I__10777 (
            .O(N__48604),
            .I(N__48601));
    LocalMux I__10776 (
            .O(N__48601),
            .I(N__48598));
    Span4Mux_v I__10775 (
            .O(N__48598),
            .I(N__48595));
    Odrv4 I__10774 (
            .O(N__48595),
            .I(\current_shift_inst.un38_control_input_0_s1_19 ));
    InMux I__10773 (
            .O(N__48592),
            .I(\current_shift_inst.un38_control_input_cry_18_s1 ));
    CascadeMux I__10772 (
            .O(N__48589),
            .I(N__48586));
    InMux I__10771 (
            .O(N__48586),
            .I(N__48583));
    LocalMux I__10770 (
            .O(N__48583),
            .I(N__48580));
    Odrv12 I__10769 (
            .O(N__48580),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ));
    InMux I__10768 (
            .O(N__48577),
            .I(N__48574));
    LocalMux I__10767 (
            .O(N__48574),
            .I(N__48571));
    Span4Mux_h I__10766 (
            .O(N__48571),
            .I(N__48568));
    Odrv4 I__10765 (
            .O(N__48568),
            .I(\current_shift_inst.un38_control_input_0_s1_5 ));
    InMux I__10764 (
            .O(N__48565),
            .I(\current_shift_inst.un38_control_input_cry_4_s1 ));
    InMux I__10763 (
            .O(N__48562),
            .I(N__48559));
    LocalMux I__10762 (
            .O(N__48559),
            .I(N__48556));
    Odrv12 I__10761 (
            .O(N__48556),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ));
    InMux I__10760 (
            .O(N__48553),
            .I(N__48550));
    LocalMux I__10759 (
            .O(N__48550),
            .I(N__48547));
    Span4Mux_v I__10758 (
            .O(N__48547),
            .I(N__48544));
    Odrv4 I__10757 (
            .O(N__48544),
            .I(\current_shift_inst.un38_control_input_0_s1_6 ));
    InMux I__10756 (
            .O(N__48541),
            .I(\current_shift_inst.un38_control_input_cry_5_s1 ));
    CascadeMux I__10755 (
            .O(N__48538),
            .I(N__48535));
    InMux I__10754 (
            .O(N__48535),
            .I(N__48532));
    LocalMux I__10753 (
            .O(N__48532),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ));
    InMux I__10752 (
            .O(N__48529),
            .I(N__48526));
    LocalMux I__10751 (
            .O(N__48526),
            .I(N__48523));
    Span4Mux_h I__10750 (
            .O(N__48523),
            .I(N__48520));
    Odrv4 I__10749 (
            .O(N__48520),
            .I(\current_shift_inst.un38_control_input_0_s1_7 ));
    InMux I__10748 (
            .O(N__48517),
            .I(\current_shift_inst.un38_control_input_cry_6_s1 ));
    CascadeMux I__10747 (
            .O(N__48514),
            .I(N__48511));
    InMux I__10746 (
            .O(N__48511),
            .I(N__48508));
    LocalMux I__10745 (
            .O(N__48508),
            .I(N__48505));
    Span4Mux_v I__10744 (
            .O(N__48505),
            .I(N__48502));
    Odrv4 I__10743 (
            .O(N__48502),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ));
    InMux I__10742 (
            .O(N__48499),
            .I(N__48496));
    LocalMux I__10741 (
            .O(N__48496),
            .I(N__48493));
    Span4Mux_h I__10740 (
            .O(N__48493),
            .I(N__48490));
    Odrv4 I__10739 (
            .O(N__48490),
            .I(\current_shift_inst.un38_control_input_0_s1_8 ));
    InMux I__10738 (
            .O(N__48487),
            .I(bfn_18_18_0_));
    InMux I__10737 (
            .O(N__48484),
            .I(N__48481));
    LocalMux I__10736 (
            .O(N__48481),
            .I(N__48478));
    Span4Mux_v I__10735 (
            .O(N__48478),
            .I(N__48475));
    Odrv4 I__10734 (
            .O(N__48475),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ));
    InMux I__10733 (
            .O(N__48472),
            .I(N__48469));
    LocalMux I__10732 (
            .O(N__48469),
            .I(N__48466));
    Span4Mux_h I__10731 (
            .O(N__48466),
            .I(N__48463));
    Odrv4 I__10730 (
            .O(N__48463),
            .I(\current_shift_inst.un38_control_input_0_s1_9 ));
    InMux I__10729 (
            .O(N__48460),
            .I(\current_shift_inst.un38_control_input_cry_8_s1 ));
    CascadeMux I__10728 (
            .O(N__48457),
            .I(N__48454));
    InMux I__10727 (
            .O(N__48454),
            .I(N__48451));
    LocalMux I__10726 (
            .O(N__48451),
            .I(N__48448));
    Odrv12 I__10725 (
            .O(N__48448),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ));
    InMux I__10724 (
            .O(N__48445),
            .I(N__48442));
    LocalMux I__10723 (
            .O(N__48442),
            .I(N__48439));
    Span4Mux_v I__10722 (
            .O(N__48439),
            .I(N__48436));
    Odrv4 I__10721 (
            .O(N__48436),
            .I(\current_shift_inst.un38_control_input_0_s1_10 ));
    InMux I__10720 (
            .O(N__48433),
            .I(\current_shift_inst.un38_control_input_cry_9_s1 ));
    InMux I__10719 (
            .O(N__48430),
            .I(N__48427));
    LocalMux I__10718 (
            .O(N__48427),
            .I(N__48424));
    Odrv12 I__10717 (
            .O(N__48424),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ));
    InMux I__10716 (
            .O(N__48421),
            .I(N__48418));
    LocalMux I__10715 (
            .O(N__48418),
            .I(N__48415));
    Span4Mux_v I__10714 (
            .O(N__48415),
            .I(N__48412));
    Odrv4 I__10713 (
            .O(N__48412),
            .I(\current_shift_inst.un38_control_input_0_s1_11 ));
    InMux I__10712 (
            .O(N__48409),
            .I(\current_shift_inst.un38_control_input_cry_10_s1 ));
    CascadeMux I__10711 (
            .O(N__48406),
            .I(N__48403));
    InMux I__10710 (
            .O(N__48403),
            .I(N__48400));
    LocalMux I__10709 (
            .O(N__48400),
            .I(N__48397));
    Odrv4 I__10708 (
            .O(N__48397),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ));
    InMux I__10707 (
            .O(N__48394),
            .I(N__48390));
    InMux I__10706 (
            .O(N__48393),
            .I(N__48387));
    LocalMux I__10705 (
            .O(N__48390),
            .I(N__48381));
    LocalMux I__10704 (
            .O(N__48387),
            .I(N__48381));
    InMux I__10703 (
            .O(N__48386),
            .I(N__48378));
    Span4Mux_v I__10702 (
            .O(N__48381),
            .I(N__48373));
    LocalMux I__10701 (
            .O(N__48378),
            .I(N__48373));
    Span4Mux_h I__10700 (
            .O(N__48373),
            .I(N__48369));
    InMux I__10699 (
            .O(N__48372),
            .I(N__48366));
    Odrv4 I__10698 (
            .O(N__48369),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    LocalMux I__10697 (
            .O(N__48366),
            .I(\current_shift_inst.elapsed_time_ns_s1_4 ));
    InMux I__10696 (
            .O(N__48361),
            .I(N__48357));
    CascadeMux I__10695 (
            .O(N__48360),
            .I(N__48354));
    LocalMux I__10694 (
            .O(N__48357),
            .I(N__48351));
    InMux I__10693 (
            .O(N__48354),
            .I(N__48347));
    Span4Mux_h I__10692 (
            .O(N__48351),
            .I(N__48344));
    InMux I__10691 (
            .O(N__48350),
            .I(N__48341));
    LocalMux I__10690 (
            .O(N__48347),
            .I(\current_shift_inst.un4_control_input1_4 ));
    Odrv4 I__10689 (
            .O(N__48344),
            .I(\current_shift_inst.un4_control_input1_4 ));
    LocalMux I__10688 (
            .O(N__48341),
            .I(\current_shift_inst.un4_control_input1_4 ));
    InMux I__10687 (
            .O(N__48334),
            .I(N__48331));
    LocalMux I__10686 (
            .O(N__48331),
            .I(N__48328));
    Span4Mux_v I__10685 (
            .O(N__48328),
            .I(N__48323));
    InMux I__10684 (
            .O(N__48327),
            .I(N__48318));
    InMux I__10683 (
            .O(N__48326),
            .I(N__48318));
    Odrv4 I__10682 (
            .O(N__48323),
            .I(\current_shift_inst.un4_control_input1_2 ));
    LocalMux I__10681 (
            .O(N__48318),
            .I(\current_shift_inst.un4_control_input1_2 ));
    CascadeMux I__10680 (
            .O(N__48313),
            .I(N__48310));
    InMux I__10679 (
            .O(N__48310),
            .I(N__48307));
    LocalMux I__10678 (
            .O(N__48307),
            .I(N__48304));
    Span4Mux_v I__10677 (
            .O(N__48304),
            .I(N__48298));
    InMux I__10676 (
            .O(N__48303),
            .I(N__48291));
    InMux I__10675 (
            .O(N__48302),
            .I(N__48291));
    InMux I__10674 (
            .O(N__48301),
            .I(N__48291));
    Odrv4 I__10673 (
            .O(N__48298),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    LocalMux I__10672 (
            .O(N__48291),
            .I(\current_shift_inst.elapsed_time_ns_s1_2 ));
    CascadeMux I__10671 (
            .O(N__48286),
            .I(N__48283));
    InMux I__10670 (
            .O(N__48283),
            .I(N__48280));
    LocalMux I__10669 (
            .O(N__48280),
            .I(N__48277));
    Odrv4 I__10668 (
            .O(N__48277),
            .I(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ));
    InMux I__10667 (
            .O(N__48274),
            .I(N__48268));
    InMux I__10666 (
            .O(N__48273),
            .I(N__48268));
    LocalMux I__10665 (
            .O(N__48268),
            .I(N__48265));
    Span4Mux_h I__10664 (
            .O(N__48265),
            .I(N__48261));
    InMux I__10663 (
            .O(N__48264),
            .I(N__48258));
    Odrv4 I__10662 (
            .O(N__48261),
            .I(\current_shift_inst.un4_control_input1_8 ));
    LocalMux I__10661 (
            .O(N__48258),
            .I(\current_shift_inst.un4_control_input1_8 ));
    CascadeMux I__10660 (
            .O(N__48253),
            .I(N__48250));
    InMux I__10659 (
            .O(N__48250),
            .I(N__48244));
    InMux I__10658 (
            .O(N__48249),
            .I(N__48244));
    LocalMux I__10657 (
            .O(N__48244),
            .I(N__48239));
    InMux I__10656 (
            .O(N__48243),
            .I(N__48234));
    InMux I__10655 (
            .O(N__48242),
            .I(N__48234));
    Span4Mux_v I__10654 (
            .O(N__48239),
            .I(N__48231));
    LocalMux I__10653 (
            .O(N__48234),
            .I(N__48228));
    Odrv4 I__10652 (
            .O(N__48231),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    Odrv4 I__10651 (
            .O(N__48228),
            .I(\current_shift_inst.elapsed_time_ns_s1_8 ));
    CascadeMux I__10650 (
            .O(N__48223),
            .I(N__48220));
    InMux I__10649 (
            .O(N__48220),
            .I(N__48217));
    LocalMux I__10648 (
            .O(N__48217),
            .I(N__48214));
    Span4Mux_v I__10647 (
            .O(N__48214),
            .I(N__48210));
    InMux I__10646 (
            .O(N__48213),
            .I(N__48207));
    Span4Mux_v I__10645 (
            .O(N__48210),
            .I(N__48202));
    LocalMux I__10644 (
            .O(N__48207),
            .I(N__48199));
    InMux I__10643 (
            .O(N__48206),
            .I(N__48196));
    InMux I__10642 (
            .O(N__48205),
            .I(N__48193));
    Odrv4 I__10641 (
            .O(N__48202),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    Odrv4 I__10640 (
            .O(N__48199),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__10639 (
            .O(N__48196),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    LocalMux I__10638 (
            .O(N__48193),
            .I(\current_shift_inst.un38_control_input_5_1 ));
    CascadeMux I__10637 (
            .O(N__48184),
            .I(N__48181));
    InMux I__10636 (
            .O(N__48181),
            .I(N__48178));
    LocalMux I__10635 (
            .O(N__48178),
            .I(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ));
    InMux I__10634 (
            .O(N__48175),
            .I(N__48172));
    LocalMux I__10633 (
            .O(N__48172),
            .I(N__48169));
    Odrv4 I__10632 (
            .O(N__48169),
            .I(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ));
    CascadeMux I__10631 (
            .O(N__48166),
            .I(N__48163));
    InMux I__10630 (
            .O(N__48163),
            .I(N__48160));
    LocalMux I__10629 (
            .O(N__48160),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ));
    InMux I__10628 (
            .O(N__48157),
            .I(N__48154));
    LocalMux I__10627 (
            .O(N__48154),
            .I(N__48151));
    Span4Mux_v I__10626 (
            .O(N__48151),
            .I(N__48148));
    Odrv4 I__10625 (
            .O(N__48148),
            .I(\current_shift_inst.un38_control_input_0_s1_3 ));
    InMux I__10624 (
            .O(N__48145),
            .I(\current_shift_inst.un38_control_input_cry_2_s1 ));
    InMux I__10623 (
            .O(N__48142),
            .I(N__48139));
    LocalMux I__10622 (
            .O(N__48139),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ));
    InMux I__10621 (
            .O(N__48136),
            .I(N__48133));
    LocalMux I__10620 (
            .O(N__48133),
            .I(N__48130));
    Span4Mux_h I__10619 (
            .O(N__48130),
            .I(N__48127));
    Odrv4 I__10618 (
            .O(N__48127),
            .I(\current_shift_inst.un38_control_input_0_s1_4 ));
    InMux I__10617 (
            .O(N__48124),
            .I(\current_shift_inst.un38_control_input_cry_3_s1 ));
    InMux I__10616 (
            .O(N__48121),
            .I(N__48118));
    LocalMux I__10615 (
            .O(N__48118),
            .I(N__48112));
    InMux I__10614 (
            .O(N__48117),
            .I(N__48109));
    InMux I__10613 (
            .O(N__48116),
            .I(N__48104));
    InMux I__10612 (
            .O(N__48115),
            .I(N__48104));
    Odrv12 I__10611 (
            .O(N__48112),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__10610 (
            .O(N__48109),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    LocalMux I__10609 (
            .O(N__48104),
            .I(\current_shift_inst.elapsed_time_ns_s1_9 ));
    InMux I__10608 (
            .O(N__48097),
            .I(N__48093));
    InMux I__10607 (
            .O(N__48096),
            .I(N__48090));
    LocalMux I__10606 (
            .O(N__48093),
            .I(N__48087));
    LocalMux I__10605 (
            .O(N__48090),
            .I(N__48084));
    Span4Mux_h I__10604 (
            .O(N__48087),
            .I(N__48078));
    Span4Mux_h I__10603 (
            .O(N__48084),
            .I(N__48078));
    InMux I__10602 (
            .O(N__48083),
            .I(N__48075));
    Odrv4 I__10601 (
            .O(N__48078),
            .I(\current_shift_inst.un4_control_input1_9 ));
    LocalMux I__10600 (
            .O(N__48075),
            .I(\current_shift_inst.un4_control_input1_9 ));
    CascadeMux I__10599 (
            .O(N__48070),
            .I(N__48067));
    InMux I__10598 (
            .O(N__48067),
            .I(N__48063));
    InMux I__10597 (
            .O(N__48066),
            .I(N__48060));
    LocalMux I__10596 (
            .O(N__48063),
            .I(N__48054));
    LocalMux I__10595 (
            .O(N__48060),
            .I(N__48054));
    InMux I__10594 (
            .O(N__48059),
            .I(N__48051));
    Span4Mux_v I__10593 (
            .O(N__48054),
            .I(N__48045));
    LocalMux I__10592 (
            .O(N__48051),
            .I(N__48045));
    InMux I__10591 (
            .O(N__48050),
            .I(N__48042));
    Odrv4 I__10590 (
            .O(N__48045),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    LocalMux I__10589 (
            .O(N__48042),
            .I(\current_shift_inst.elapsed_time_ns_s1_23 ));
    CascadeMux I__10588 (
            .O(N__48037),
            .I(N__48034));
    InMux I__10587 (
            .O(N__48034),
            .I(N__48029));
    InMux I__10586 (
            .O(N__48033),
            .I(N__48026));
    InMux I__10585 (
            .O(N__48032),
            .I(N__48023));
    LocalMux I__10584 (
            .O(N__48029),
            .I(N__48020));
    LocalMux I__10583 (
            .O(N__48026),
            .I(N__48017));
    LocalMux I__10582 (
            .O(N__48023),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv12 I__10581 (
            .O(N__48020),
            .I(\current_shift_inst.un4_control_input1_23 ));
    Odrv4 I__10580 (
            .O(N__48017),
            .I(\current_shift_inst.un4_control_input1_23 ));
    CascadeMux I__10579 (
            .O(N__48010),
            .I(N__48007));
    InMux I__10578 (
            .O(N__48007),
            .I(N__48002));
    InMux I__10577 (
            .O(N__48006),
            .I(N__47999));
    InMux I__10576 (
            .O(N__48005),
            .I(N__47996));
    LocalMux I__10575 (
            .O(N__48002),
            .I(N__47993));
    LocalMux I__10574 (
            .O(N__47999),
            .I(N__47990));
    LocalMux I__10573 (
            .O(N__47996),
            .I(N__47987));
    Span4Mux_h I__10572 (
            .O(N__47993),
            .I(N__47983));
    Span4Mux_h I__10571 (
            .O(N__47990),
            .I(N__47980));
    Span4Mux_v I__10570 (
            .O(N__47987),
            .I(N__47977));
    InMux I__10569 (
            .O(N__47986),
            .I(N__47974));
    Odrv4 I__10568 (
            .O(N__47983),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10567 (
            .O(N__47980),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    Odrv4 I__10566 (
            .O(N__47977),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    LocalMux I__10565 (
            .O(N__47974),
            .I(\current_shift_inst.elapsed_time_ns_s1_24 ));
    InMux I__10564 (
            .O(N__47965),
            .I(N__47961));
    InMux I__10563 (
            .O(N__47964),
            .I(N__47957));
    LocalMux I__10562 (
            .O(N__47961),
            .I(N__47954));
    InMux I__10561 (
            .O(N__47960),
            .I(N__47951));
    LocalMux I__10560 (
            .O(N__47957),
            .I(N__47948));
    Span4Mux_v I__10559 (
            .O(N__47954),
            .I(N__47945));
    LocalMux I__10558 (
            .O(N__47951),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__10557 (
            .O(N__47948),
            .I(\current_shift_inst.un4_control_input1_24 ));
    Odrv4 I__10556 (
            .O(N__47945),
            .I(\current_shift_inst.un4_control_input1_24 ));
    InMux I__10555 (
            .O(N__47938),
            .I(N__47935));
    LocalMux I__10554 (
            .O(N__47935),
            .I(N__47931));
    InMux I__10553 (
            .O(N__47934),
            .I(N__47927));
    Span4Mux_v I__10552 (
            .O(N__47931),
            .I(N__47924));
    InMux I__10551 (
            .O(N__47930),
            .I(N__47921));
    LocalMux I__10550 (
            .O(N__47927),
            .I(\current_shift_inst.un4_control_input1_18 ));
    Odrv4 I__10549 (
            .O(N__47924),
            .I(\current_shift_inst.un4_control_input1_18 ));
    LocalMux I__10548 (
            .O(N__47921),
            .I(\current_shift_inst.un4_control_input1_18 ));
    CascadeMux I__10547 (
            .O(N__47914),
            .I(N__47911));
    InMux I__10546 (
            .O(N__47911),
            .I(N__47907));
    CascadeMux I__10545 (
            .O(N__47910),
            .I(N__47904));
    LocalMux I__10544 (
            .O(N__47907),
            .I(N__47901));
    InMux I__10543 (
            .O(N__47904),
            .I(N__47898));
    Span4Mux_h I__10542 (
            .O(N__47901),
            .I(N__47894));
    LocalMux I__10541 (
            .O(N__47898),
            .I(N__47891));
    InMux I__10540 (
            .O(N__47897),
            .I(N__47888));
    Span4Mux_h I__10539 (
            .O(N__47894),
            .I(N__47884));
    Span4Mux_h I__10538 (
            .O(N__47891),
            .I(N__47879));
    LocalMux I__10537 (
            .O(N__47888),
            .I(N__47879));
    InMux I__10536 (
            .O(N__47887),
            .I(N__47876));
    Odrv4 I__10535 (
            .O(N__47884),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    Odrv4 I__10534 (
            .O(N__47879),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    LocalMux I__10533 (
            .O(N__47876),
            .I(\current_shift_inst.elapsed_time_ns_s1_18 ));
    InMux I__10532 (
            .O(N__47869),
            .I(N__47862));
    InMux I__10531 (
            .O(N__47868),
            .I(N__47862));
    InMux I__10530 (
            .O(N__47867),
            .I(N__47859));
    LocalMux I__10529 (
            .O(N__47862),
            .I(N__47855));
    LocalMux I__10528 (
            .O(N__47859),
            .I(N__47852));
    InMux I__10527 (
            .O(N__47858),
            .I(N__47849));
    Span4Mux_v I__10526 (
            .O(N__47855),
            .I(N__47846));
    Span4Mux_v I__10525 (
            .O(N__47852),
            .I(N__47841));
    LocalMux I__10524 (
            .O(N__47849),
            .I(N__47841));
    Span4Mux_v I__10523 (
            .O(N__47846),
            .I(N__47838));
    Span4Mux_h I__10522 (
            .O(N__47841),
            .I(N__47835));
    Odrv4 I__10521 (
            .O(N__47838),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    Odrv4 I__10520 (
            .O(N__47835),
            .I(\current_shift_inst.elapsed_time_ns_s1_19 ));
    CascadeMux I__10519 (
            .O(N__47830),
            .I(N__47826));
    InMux I__10518 (
            .O(N__47829),
            .I(N__47822));
    InMux I__10517 (
            .O(N__47826),
            .I(N__47817));
    InMux I__10516 (
            .O(N__47825),
            .I(N__47817));
    LocalMux I__10515 (
            .O(N__47822),
            .I(N__47814));
    LocalMux I__10514 (
            .O(N__47817),
            .I(N__47811));
    Odrv4 I__10513 (
            .O(N__47814),
            .I(\current_shift_inst.un4_control_input1_19 ));
    Odrv4 I__10512 (
            .O(N__47811),
            .I(\current_shift_inst.un4_control_input1_19 ));
    InMux I__10511 (
            .O(N__47806),
            .I(N__47803));
    LocalMux I__10510 (
            .O(N__47803),
            .I(N__47798));
    InMux I__10509 (
            .O(N__47802),
            .I(N__47795));
    InMux I__10508 (
            .O(N__47801),
            .I(N__47792));
    Span12Mux_s9_h I__10507 (
            .O(N__47798),
            .I(N__47789));
    LocalMux I__10506 (
            .O(N__47795),
            .I(N__47786));
    LocalMux I__10505 (
            .O(N__47792),
            .I(N__47783));
    Odrv12 I__10504 (
            .O(N__47789),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv12 I__10503 (
            .O(N__47786),
            .I(\current_shift_inst.un4_control_input1_20 ));
    Odrv4 I__10502 (
            .O(N__47783),
            .I(\current_shift_inst.un4_control_input1_20 ));
    CascadeMux I__10501 (
            .O(N__47776),
            .I(N__47772));
    CascadeMux I__10500 (
            .O(N__47775),
            .I(N__47769));
    InMux I__10499 (
            .O(N__47772),
            .I(N__47765));
    InMux I__10498 (
            .O(N__47769),
            .I(N__47762));
    InMux I__10497 (
            .O(N__47768),
            .I(N__47759));
    LocalMux I__10496 (
            .O(N__47765),
            .I(N__47755));
    LocalMux I__10495 (
            .O(N__47762),
            .I(N__47750));
    LocalMux I__10494 (
            .O(N__47759),
            .I(N__47750));
    InMux I__10493 (
            .O(N__47758),
            .I(N__47747));
    Span4Mux_h I__10492 (
            .O(N__47755),
            .I(N__47744));
    Span4Mux_h I__10491 (
            .O(N__47750),
            .I(N__47741));
    LocalMux I__10490 (
            .O(N__47747),
            .I(N__47738));
    Odrv4 I__10489 (
            .O(N__47744),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10488 (
            .O(N__47741),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    Odrv4 I__10487 (
            .O(N__47738),
            .I(\current_shift_inst.elapsed_time_ns_s1_20 ));
    CascadeMux I__10486 (
            .O(N__47731),
            .I(N__47728));
    InMux I__10485 (
            .O(N__47728),
            .I(N__47724));
    InMux I__10484 (
            .O(N__47727),
            .I(N__47721));
    LocalMux I__10483 (
            .O(N__47724),
            .I(N__47716));
    LocalMux I__10482 (
            .O(N__47721),
            .I(N__47713));
    InMux I__10481 (
            .O(N__47720),
            .I(N__47710));
    InMux I__10480 (
            .O(N__47719),
            .I(N__47707));
    Odrv4 I__10479 (
            .O(N__47716),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    Odrv12 I__10478 (
            .O(N__47713),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__10477 (
            .O(N__47710),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    LocalMux I__10476 (
            .O(N__47707),
            .I(\current_shift_inst.elapsed_time_ns_s1_14 ));
    InMux I__10475 (
            .O(N__47698),
            .I(N__47695));
    LocalMux I__10474 (
            .O(N__47695),
            .I(N__47691));
    InMux I__10473 (
            .O(N__47694),
            .I(N__47688));
    Span4Mux_h I__10472 (
            .O(N__47691),
            .I(N__47684));
    LocalMux I__10471 (
            .O(N__47688),
            .I(N__47681));
    InMux I__10470 (
            .O(N__47687),
            .I(N__47678));
    Odrv4 I__10469 (
            .O(N__47684),
            .I(\current_shift_inst.un4_control_input1_14 ));
    Odrv4 I__10468 (
            .O(N__47681),
            .I(\current_shift_inst.un4_control_input1_14 ));
    LocalMux I__10467 (
            .O(N__47678),
            .I(\current_shift_inst.un4_control_input1_14 ));
    CascadeMux I__10466 (
            .O(N__47671),
            .I(N__47668));
    InMux I__10465 (
            .O(N__47668),
            .I(N__47665));
    LocalMux I__10464 (
            .O(N__47665),
            .I(N__47661));
    InMux I__10463 (
            .O(N__47664),
            .I(N__47657));
    Span4Mux_h I__10462 (
            .O(N__47661),
            .I(N__47654));
    InMux I__10461 (
            .O(N__47660),
            .I(N__47651));
    LocalMux I__10460 (
            .O(N__47657),
            .I(\current_shift_inst.un4_control_input1_6 ));
    Odrv4 I__10459 (
            .O(N__47654),
            .I(\current_shift_inst.un4_control_input1_6 ));
    LocalMux I__10458 (
            .O(N__47651),
            .I(\current_shift_inst.un4_control_input1_6 ));
    CascadeMux I__10457 (
            .O(N__47644),
            .I(N__47641));
    InMux I__10456 (
            .O(N__47641),
            .I(N__47637));
    InMux I__10455 (
            .O(N__47640),
            .I(N__47634));
    LocalMux I__10454 (
            .O(N__47637),
            .I(N__47630));
    LocalMux I__10453 (
            .O(N__47634),
            .I(N__47627));
    InMux I__10452 (
            .O(N__47633),
            .I(N__47624));
    Span4Mux_h I__10451 (
            .O(N__47630),
            .I(N__47620));
    Span4Mux_h I__10450 (
            .O(N__47627),
            .I(N__47615));
    LocalMux I__10449 (
            .O(N__47624),
            .I(N__47615));
    InMux I__10448 (
            .O(N__47623),
            .I(N__47612));
    Odrv4 I__10447 (
            .O(N__47620),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    Odrv4 I__10446 (
            .O(N__47615),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    LocalMux I__10445 (
            .O(N__47612),
            .I(\current_shift_inst.elapsed_time_ns_s1_6 ));
    InMux I__10444 (
            .O(N__47605),
            .I(N__47601));
    InMux I__10443 (
            .O(N__47604),
            .I(N__47598));
    LocalMux I__10442 (
            .O(N__47601),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    LocalMux I__10441 (
            .O(N__47598),
            .I(elapsed_time_ns_1_RNIV1DN9_0_21));
    InMux I__10440 (
            .O(N__47593),
            .I(N__47590));
    LocalMux I__10439 (
            .O(N__47590),
            .I(N__47587));
    Span4Mux_h I__10438 (
            .O(N__47587),
            .I(N__47584));
    Odrv4 I__10437 (
            .O(N__47584),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ));
    InMux I__10436 (
            .O(N__47581),
            .I(N__47577));
    InMux I__10435 (
            .O(N__47580),
            .I(N__47574));
    LocalMux I__10434 (
            .O(N__47577),
            .I(N__47571));
    LocalMux I__10433 (
            .O(N__47574),
            .I(N__47568));
    Span4Mux_v I__10432 (
            .O(N__47571),
            .I(N__47565));
    Span4Mux_v I__10431 (
            .O(N__47568),
            .I(N__47560));
    Span4Mux_h I__10430 (
            .O(N__47565),
            .I(N__47557));
    InMux I__10429 (
            .O(N__47564),
            .I(N__47552));
    InMux I__10428 (
            .O(N__47563),
            .I(N__47552));
    Span4Mux_v I__10427 (
            .O(N__47560),
            .I(N__47549));
    Span4Mux_v I__10426 (
            .O(N__47557),
            .I(N__47546));
    LocalMux I__10425 (
            .O(N__47552),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__10424 (
            .O(N__47549),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    Odrv4 I__10423 (
            .O(N__47546),
            .I(\delay_measurement_inst.start_timer_hcZ0 ));
    InMux I__10422 (
            .O(N__47539),
            .I(N__47536));
    LocalMux I__10421 (
            .O(N__47536),
            .I(N__47531));
    InMux I__10420 (
            .O(N__47535),
            .I(N__47528));
    CascadeMux I__10419 (
            .O(N__47534),
            .I(N__47525));
    Span4Mux_v I__10418 (
            .O(N__47531),
            .I(N__47519));
    LocalMux I__10417 (
            .O(N__47528),
            .I(N__47519));
    InMux I__10416 (
            .O(N__47525),
            .I(N__47514));
    InMux I__10415 (
            .O(N__47524),
            .I(N__47514));
    Span4Mux_h I__10414 (
            .O(N__47519),
            .I(N__47511));
    LocalMux I__10413 (
            .O(N__47514),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    Odrv4 I__10412 (
            .O(N__47511),
            .I(\delay_measurement_inst.delay_hc_timer.runningZ0 ));
    InMux I__10411 (
            .O(N__47506),
            .I(N__47503));
    LocalMux I__10410 (
            .O(N__47503),
            .I(N__47498));
    InMux I__10409 (
            .O(N__47502),
            .I(N__47493));
    InMux I__10408 (
            .O(N__47501),
            .I(N__47493));
    Span4Mux_v I__10407 (
            .O(N__47498),
            .I(N__47490));
    LocalMux I__10406 (
            .O(N__47493),
            .I(N__47487));
    Span4Mux_h I__10405 (
            .O(N__47490),
            .I(N__47484));
    Span4Mux_v I__10404 (
            .O(N__47487),
            .I(N__47481));
    Span4Mux_v I__10403 (
            .O(N__47484),
            .I(N__47478));
    Span4Mux_v I__10402 (
            .O(N__47481),
            .I(N__47475));
    Odrv4 I__10401 (
            .O(N__47478),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    Odrv4 I__10400 (
            .O(N__47475),
            .I(\delay_measurement_inst.stop_timer_hcZ0 ));
    CEMux I__10399 (
            .O(N__47470),
            .I(N__47464));
    CEMux I__10398 (
            .O(N__47469),
            .I(N__47461));
    CEMux I__10397 (
            .O(N__47468),
            .I(N__47458));
    CEMux I__10396 (
            .O(N__47467),
            .I(N__47455));
    LocalMux I__10395 (
            .O(N__47464),
            .I(N__47452));
    LocalMux I__10394 (
            .O(N__47461),
            .I(N__47447));
    LocalMux I__10393 (
            .O(N__47458),
            .I(N__47447));
    LocalMux I__10392 (
            .O(N__47455),
            .I(N__47444));
    Span4Mux_v I__10391 (
            .O(N__47452),
            .I(N__47437));
    Span4Mux_v I__10390 (
            .O(N__47447),
            .I(N__47437));
    Span4Mux_h I__10389 (
            .O(N__47444),
            .I(N__47437));
    Odrv4 I__10388 (
            .O(N__47437),
            .I(\delay_measurement_inst.delay_hc_timer.N_166_i ));
    InMux I__10387 (
            .O(N__47434),
            .I(N__47430));
    InMux I__10386 (
            .O(N__47433),
            .I(N__47427));
    LocalMux I__10385 (
            .O(N__47430),
            .I(N__47421));
    LocalMux I__10384 (
            .O(N__47427),
            .I(N__47421));
    InMux I__10383 (
            .O(N__47426),
            .I(N__47418));
    Span4Mux_v I__10382 (
            .O(N__47421),
            .I(N__47413));
    LocalMux I__10381 (
            .O(N__47418),
            .I(N__47413));
    Span4Mux_h I__10380 (
            .O(N__47413),
            .I(N__47409));
    InMux I__10379 (
            .O(N__47412),
            .I(N__47406));
    Odrv4 I__10378 (
            .O(N__47409),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    LocalMux I__10377 (
            .O(N__47406),
            .I(\current_shift_inst.elapsed_time_ns_s1_17 ));
    CascadeMux I__10376 (
            .O(N__47401),
            .I(N__47397));
    CascadeMux I__10375 (
            .O(N__47400),
            .I(N__47394));
    InMux I__10374 (
            .O(N__47397),
            .I(N__47390));
    InMux I__10373 (
            .O(N__47394),
            .I(N__47387));
    InMux I__10372 (
            .O(N__47393),
            .I(N__47384));
    LocalMux I__10371 (
            .O(N__47390),
            .I(N__47379));
    LocalMux I__10370 (
            .O(N__47387),
            .I(N__47379));
    LocalMux I__10369 (
            .O(N__47384),
            .I(N__47376));
    Odrv4 I__10368 (
            .O(N__47379),
            .I(\current_shift_inst.un4_control_input1_17 ));
    Odrv4 I__10367 (
            .O(N__47376),
            .I(\current_shift_inst.un4_control_input1_17 ));
    CEMux I__10366 (
            .O(N__47371),
            .I(N__47368));
    LocalMux I__10365 (
            .O(N__47368),
            .I(N__47364));
    CEMux I__10364 (
            .O(N__47367),
            .I(N__47361));
    Span4Mux_v I__10363 (
            .O(N__47364),
            .I(N__47357));
    LocalMux I__10362 (
            .O(N__47361),
            .I(N__47354));
    CEMux I__10361 (
            .O(N__47360),
            .I(N__47350));
    Span4Mux_h I__10360 (
            .O(N__47357),
            .I(N__47345));
    Span4Mux_h I__10359 (
            .O(N__47354),
            .I(N__47345));
    CEMux I__10358 (
            .O(N__47353),
            .I(N__47342));
    LocalMux I__10357 (
            .O(N__47350),
            .I(N__47339));
    Span4Mux_h I__10356 (
            .O(N__47345),
            .I(N__47336));
    LocalMux I__10355 (
            .O(N__47342),
            .I(N__47333));
    Span4Mux_h I__10354 (
            .O(N__47339),
            .I(N__47330));
    Span4Mux_h I__10353 (
            .O(N__47336),
            .I(N__47327));
    Odrv12 I__10352 (
            .O(N__47333),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    Odrv4 I__10351 (
            .O(N__47330),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    Odrv4 I__10350 (
            .O(N__47327),
            .I(\current_shift_inst.timer_s1.N_164_i ));
    InMux I__10349 (
            .O(N__47320),
            .I(N__47316));
    InMux I__10348 (
            .O(N__47319),
            .I(N__47312));
    LocalMux I__10347 (
            .O(N__47316),
            .I(N__47309));
    InMux I__10346 (
            .O(N__47315),
            .I(N__47306));
    LocalMux I__10345 (
            .O(N__47312),
            .I(\current_shift_inst.un4_control_input1_12 ));
    Odrv12 I__10344 (
            .O(N__47309),
            .I(\current_shift_inst.un4_control_input1_12 ));
    LocalMux I__10343 (
            .O(N__47306),
            .I(\current_shift_inst.un4_control_input1_12 ));
    CascadeMux I__10342 (
            .O(N__47299),
            .I(N__47295));
    CascadeMux I__10341 (
            .O(N__47298),
            .I(N__47292));
    InMux I__10340 (
            .O(N__47295),
            .I(N__47289));
    InMux I__10339 (
            .O(N__47292),
            .I(N__47286));
    LocalMux I__10338 (
            .O(N__47289),
            .I(N__47282));
    LocalMux I__10337 (
            .O(N__47286),
            .I(N__47279));
    InMux I__10336 (
            .O(N__47285),
            .I(N__47276));
    Span4Mux_h I__10335 (
            .O(N__47282),
            .I(N__47270));
    Span4Mux_h I__10334 (
            .O(N__47279),
            .I(N__47270));
    LocalMux I__10333 (
            .O(N__47276),
            .I(N__47267));
    InMux I__10332 (
            .O(N__47275),
            .I(N__47264));
    Odrv4 I__10331 (
            .O(N__47270),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    Odrv4 I__10330 (
            .O(N__47267),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    LocalMux I__10329 (
            .O(N__47264),
            .I(\current_shift_inst.elapsed_time_ns_s1_12 ));
    InMux I__10328 (
            .O(N__47257),
            .I(N__47219));
    InMux I__10327 (
            .O(N__47256),
            .I(N__47219));
    InMux I__10326 (
            .O(N__47255),
            .I(N__47219));
    InMux I__10325 (
            .O(N__47254),
            .I(N__47219));
    InMux I__10324 (
            .O(N__47253),
            .I(N__47210));
    InMux I__10323 (
            .O(N__47252),
            .I(N__47210));
    InMux I__10322 (
            .O(N__47251),
            .I(N__47210));
    InMux I__10321 (
            .O(N__47250),
            .I(N__47210));
    InMux I__10320 (
            .O(N__47249),
            .I(N__47201));
    InMux I__10319 (
            .O(N__47248),
            .I(N__47201));
    InMux I__10318 (
            .O(N__47247),
            .I(N__47201));
    InMux I__10317 (
            .O(N__47246),
            .I(N__47201));
    InMux I__10316 (
            .O(N__47245),
            .I(N__47192));
    InMux I__10315 (
            .O(N__47244),
            .I(N__47192));
    InMux I__10314 (
            .O(N__47243),
            .I(N__47192));
    InMux I__10313 (
            .O(N__47242),
            .I(N__47192));
    InMux I__10312 (
            .O(N__47241),
            .I(N__47183));
    InMux I__10311 (
            .O(N__47240),
            .I(N__47183));
    InMux I__10310 (
            .O(N__47239),
            .I(N__47183));
    InMux I__10309 (
            .O(N__47238),
            .I(N__47183));
    InMux I__10308 (
            .O(N__47237),
            .I(N__47174));
    InMux I__10307 (
            .O(N__47236),
            .I(N__47174));
    InMux I__10306 (
            .O(N__47235),
            .I(N__47174));
    InMux I__10305 (
            .O(N__47234),
            .I(N__47174));
    InMux I__10304 (
            .O(N__47233),
            .I(N__47169));
    InMux I__10303 (
            .O(N__47232),
            .I(N__47169));
    InMux I__10302 (
            .O(N__47231),
            .I(N__47160));
    InMux I__10301 (
            .O(N__47230),
            .I(N__47160));
    InMux I__10300 (
            .O(N__47229),
            .I(N__47160));
    InMux I__10299 (
            .O(N__47228),
            .I(N__47160));
    LocalMux I__10298 (
            .O(N__47219),
            .I(N__47157));
    LocalMux I__10297 (
            .O(N__47210),
            .I(N__47146));
    LocalMux I__10296 (
            .O(N__47201),
            .I(N__47146));
    LocalMux I__10295 (
            .O(N__47192),
            .I(N__47146));
    LocalMux I__10294 (
            .O(N__47183),
            .I(N__47146));
    LocalMux I__10293 (
            .O(N__47174),
            .I(N__47146));
    LocalMux I__10292 (
            .O(N__47169),
            .I(N__47137));
    LocalMux I__10291 (
            .O(N__47160),
            .I(N__47137));
    Span4Mux_v I__10290 (
            .O(N__47157),
            .I(N__47137));
    Span4Mux_v I__10289 (
            .O(N__47146),
            .I(N__47137));
    Span4Mux_h I__10288 (
            .O(N__47137),
            .I(N__47134));
    Odrv4 I__10287 (
            .O(N__47134),
            .I(\current_shift_inst.timer_s1.running_i ));
    InMux I__10286 (
            .O(N__47131),
            .I(N__47128));
    LocalMux I__10285 (
            .O(N__47128),
            .I(N__47124));
    InMux I__10284 (
            .O(N__47127),
            .I(N__47120));
    Span4Mux_h I__10283 (
            .O(N__47124),
            .I(N__47117));
    InMux I__10282 (
            .O(N__47123),
            .I(N__47114));
    LocalMux I__10281 (
            .O(N__47120),
            .I(\current_shift_inst.un4_control_input1_15 ));
    Odrv4 I__10280 (
            .O(N__47117),
            .I(\current_shift_inst.un4_control_input1_15 ));
    LocalMux I__10279 (
            .O(N__47114),
            .I(\current_shift_inst.un4_control_input1_15 ));
    CascadeMux I__10278 (
            .O(N__47107),
            .I(N__47103));
    CascadeMux I__10277 (
            .O(N__47106),
            .I(N__47100));
    InMux I__10276 (
            .O(N__47103),
            .I(N__47097));
    InMux I__10275 (
            .O(N__47100),
            .I(N__47094));
    LocalMux I__10274 (
            .O(N__47097),
            .I(N__47089));
    LocalMux I__10273 (
            .O(N__47094),
            .I(N__47089));
    Span4Mux_h I__10272 (
            .O(N__47089),
            .I(N__47084));
    InMux I__10271 (
            .O(N__47088),
            .I(N__47079));
    InMux I__10270 (
            .O(N__47087),
            .I(N__47079));
    Odrv4 I__10269 (
            .O(N__47084),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    LocalMux I__10268 (
            .O(N__47079),
            .I(\current_shift_inst.elapsed_time_ns_s1_15 ));
    CascadeMux I__10267 (
            .O(N__47074),
            .I(N__47071));
    InMux I__10266 (
            .O(N__47071),
            .I(N__47067));
    InMux I__10265 (
            .O(N__47070),
            .I(N__47064));
    LocalMux I__10264 (
            .O(N__47067),
            .I(N__47058));
    LocalMux I__10263 (
            .O(N__47064),
            .I(N__47058));
    InMux I__10262 (
            .O(N__47063),
            .I(N__47055));
    Span4Mux_h I__10261 (
            .O(N__47058),
            .I(N__47051));
    LocalMux I__10260 (
            .O(N__47055),
            .I(N__47048));
    InMux I__10259 (
            .O(N__47054),
            .I(N__47045));
    Odrv4 I__10258 (
            .O(N__47051),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    Odrv4 I__10257 (
            .O(N__47048),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    LocalMux I__10256 (
            .O(N__47045),
            .I(\current_shift_inst.elapsed_time_ns_s1_11 ));
    InMux I__10255 (
            .O(N__47038),
            .I(N__47033));
    InMux I__10254 (
            .O(N__47037),
            .I(N__47030));
    InMux I__10253 (
            .O(N__47036),
            .I(N__47027));
    LocalMux I__10252 (
            .O(N__47033),
            .I(N__47022));
    LocalMux I__10251 (
            .O(N__47030),
            .I(N__47022));
    LocalMux I__10250 (
            .O(N__47027),
            .I(\current_shift_inst.un4_control_input1_11 ));
    Odrv4 I__10249 (
            .O(N__47022),
            .I(\current_shift_inst.un4_control_input1_11 ));
    IoInMux I__10248 (
            .O(N__47017),
            .I(N__47014));
    LocalMux I__10247 (
            .O(N__47014),
            .I(N__47011));
    Span4Mux_s3_v I__10246 (
            .O(N__47011),
            .I(N__47008));
    Sp12to4 I__10245 (
            .O(N__47008),
            .I(N__47005));
    Span12Mux_s11_h I__10244 (
            .O(N__47005),
            .I(N__47002));
    Span12Mux_v I__10243 (
            .O(N__47002),
            .I(N__46999));
    Odrv12 I__10242 (
            .O(N__46999),
            .I(\current_shift_inst.timer_s1.N_163_i ));
    InMux I__10241 (
            .O(N__46996),
            .I(N__46993));
    LocalMux I__10240 (
            .O(N__46993),
            .I(N__46990));
    Span4Mux_v I__10239 (
            .O(N__46990),
            .I(N__46986));
    InMux I__10238 (
            .O(N__46989),
            .I(N__46983));
    Odrv4 I__10237 (
            .O(N__46986),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    LocalMux I__10236 (
            .O(N__46983),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ));
    InMux I__10235 (
            .O(N__46978),
            .I(N__46975));
    LocalMux I__10234 (
            .O(N__46975),
            .I(N__46972));
    Span4Mux_v I__10233 (
            .O(N__46972),
            .I(N__46968));
    InMux I__10232 (
            .O(N__46971),
            .I(N__46965));
    Odrv4 I__10231 (
            .O(N__46968),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    LocalMux I__10230 (
            .O(N__46965),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ));
    InMux I__10229 (
            .O(N__46960),
            .I(N__46957));
    LocalMux I__10228 (
            .O(N__46957),
            .I(N__46954));
    Span4Mux_v I__10227 (
            .O(N__46954),
            .I(N__46950));
    InMux I__10226 (
            .O(N__46953),
            .I(N__46947));
    Odrv4 I__10225 (
            .O(N__46950),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    LocalMux I__10224 (
            .O(N__46947),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ));
    InMux I__10223 (
            .O(N__46942),
            .I(N__46939));
    LocalMux I__10222 (
            .O(N__46939),
            .I(N__46935));
    InMux I__10221 (
            .O(N__46938),
            .I(N__46932));
    Odrv12 I__10220 (
            .O(N__46935),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    LocalMux I__10219 (
            .O(N__46932),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ));
    InMux I__10218 (
            .O(N__46927),
            .I(N__46924));
    LocalMux I__10217 (
            .O(N__46924),
            .I(N__46921));
    Span4Mux_h I__10216 (
            .O(N__46921),
            .I(N__46917));
    InMux I__10215 (
            .O(N__46920),
            .I(N__46914));
    Odrv4 I__10214 (
            .O(N__46917),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    LocalMux I__10213 (
            .O(N__46914),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ));
    CascadeMux I__10212 (
            .O(N__46909),
            .I(N__46905));
    InMux I__10211 (
            .O(N__46908),
            .I(N__46902));
    InMux I__10210 (
            .O(N__46905),
            .I(N__46899));
    LocalMux I__10209 (
            .O(N__46902),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    LocalMux I__10208 (
            .O(N__46899),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ));
    InMux I__10207 (
            .O(N__46894),
            .I(N__46891));
    LocalMux I__10206 (
            .O(N__46891),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ));
    InMux I__10205 (
            .O(N__46888),
            .I(N__46885));
    LocalMux I__10204 (
            .O(N__46885),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ));
    CascadeMux I__10203 (
            .O(N__46882),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ));
    InMux I__10202 (
            .O(N__46879),
            .I(N__46876));
    LocalMux I__10201 (
            .O(N__46876),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ));
    InMux I__10200 (
            .O(N__46873),
            .I(N__46870));
    LocalMux I__10199 (
            .O(N__46870),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ));
    CascadeMux I__10198 (
            .O(N__46867),
            .I(N__46864));
    InMux I__10197 (
            .O(N__46864),
            .I(N__46858));
    CascadeMux I__10196 (
            .O(N__46863),
            .I(N__46855));
    InMux I__10195 (
            .O(N__46862),
            .I(N__46852));
    InMux I__10194 (
            .O(N__46861),
            .I(N__46849));
    LocalMux I__10193 (
            .O(N__46858),
            .I(N__46846));
    InMux I__10192 (
            .O(N__46855),
            .I(N__46843));
    LocalMux I__10191 (
            .O(N__46852),
            .I(N__46840));
    LocalMux I__10190 (
            .O(N__46849),
            .I(N__46837));
    Span4Mux_v I__10189 (
            .O(N__46846),
            .I(N__46832));
    LocalMux I__10188 (
            .O(N__46843),
            .I(N__46832));
    Span4Mux_h I__10187 (
            .O(N__46840),
            .I(N__46829));
    Span4Mux_h I__10186 (
            .O(N__46837),
            .I(N__46826));
    Span4Mux_v I__10185 (
            .O(N__46832),
            .I(N__46821));
    Span4Mux_v I__10184 (
            .O(N__46829),
            .I(N__46821));
    Odrv4 I__10183 (
            .O(N__46826),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    Odrv4 I__10182 (
            .O(N__46821),
            .I(\current_shift_inst.elapsed_time_ns_s1_25 ));
    InMux I__10181 (
            .O(N__46816),
            .I(N__46813));
    LocalMux I__10180 (
            .O(N__46813),
            .I(N__46810));
    Span4Mux_h I__10179 (
            .O(N__46810),
            .I(N__46807));
    Odrv4 I__10178 (
            .O(N__46807),
            .I(\current_shift_inst.un4_control_input_1_axb_24 ));
    CascadeMux I__10177 (
            .O(N__46804),
            .I(N__46800));
    InMux I__10176 (
            .O(N__46803),
            .I(N__46795));
    InMux I__10175 (
            .O(N__46800),
            .I(N__46795));
    LocalMux I__10174 (
            .O(N__46795),
            .I(N__46791));
    InMux I__10173 (
            .O(N__46794),
            .I(N__46788));
    Span4Mux_h I__10172 (
            .O(N__46791),
            .I(N__46784));
    LocalMux I__10171 (
            .O(N__46788),
            .I(N__46781));
    InMux I__10170 (
            .O(N__46787),
            .I(N__46778));
    Odrv4 I__10169 (
            .O(N__46784),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    Odrv4 I__10168 (
            .O(N__46781),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    LocalMux I__10167 (
            .O(N__46778),
            .I(\current_shift_inst.elapsed_time_ns_s1_7 ));
    InMux I__10166 (
            .O(N__46771),
            .I(N__46765));
    InMux I__10165 (
            .O(N__46770),
            .I(N__46765));
    LocalMux I__10164 (
            .O(N__46765),
            .I(N__46761));
    InMux I__10163 (
            .O(N__46764),
            .I(N__46758));
    Odrv4 I__10162 (
            .O(N__46761),
            .I(\current_shift_inst.un4_control_input1_7 ));
    LocalMux I__10161 (
            .O(N__46758),
            .I(\current_shift_inst.un4_control_input1_7 ));
    CascadeMux I__10160 (
            .O(N__46753),
            .I(N__46750));
    InMux I__10159 (
            .O(N__46750),
            .I(N__46747));
    LocalMux I__10158 (
            .O(N__46747),
            .I(N__46744));
    Span4Mux_v I__10157 (
            .O(N__46744),
            .I(N__46741));
    Odrv4 I__10156 (
            .O(N__46741),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ));
    InMux I__10155 (
            .O(N__46738),
            .I(N__46734));
    InMux I__10154 (
            .O(N__46737),
            .I(N__46731));
    LocalMux I__10153 (
            .O(N__46734),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    LocalMux I__10152 (
            .O(N__46731),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ));
    InMux I__10151 (
            .O(N__46726),
            .I(N__46723));
    LocalMux I__10150 (
            .O(N__46723),
            .I(elapsed_time_ns_1_RNI68CN9_0_19));
    CascadeMux I__10149 (
            .O(N__46720),
            .I(elapsed_time_ns_1_RNI68CN9_0_19_cascade_));
    InMux I__10148 (
            .O(N__46717),
            .I(N__46714));
    LocalMux I__10147 (
            .O(N__46714),
            .I(N__46711));
    Span4Mux_v I__10146 (
            .O(N__46711),
            .I(N__46708));
    Odrv4 I__10145 (
            .O(N__46708),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ));
    CascadeMux I__10144 (
            .O(N__46705),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ));
    InMux I__10143 (
            .O(N__46702),
            .I(N__46699));
    LocalMux I__10142 (
            .O(N__46699),
            .I(N__46695));
    InMux I__10141 (
            .O(N__46698),
            .I(N__46692));
    Span4Mux_v I__10140 (
            .O(N__46695),
            .I(N__46689));
    LocalMux I__10139 (
            .O(N__46692),
            .I(N__46686));
    Odrv4 I__10138 (
            .O(N__46689),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    Odrv4 I__10137 (
            .O(N__46686),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ));
    CascadeMux I__10136 (
            .O(N__46681),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22_cascade_ ));
    InMux I__10135 (
            .O(N__46678),
            .I(N__46675));
    LocalMux I__10134 (
            .O(N__46675),
            .I(N__46672));
    Span4Mux_h I__10133 (
            .O(N__46672),
            .I(N__46669));
    Odrv4 I__10132 (
            .O(N__46669),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ));
    CascadeMux I__10131 (
            .O(N__46666),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ));
    InMux I__10130 (
            .O(N__46663),
            .I(N__46660));
    LocalMux I__10129 (
            .O(N__46660),
            .I(N__46656));
    InMux I__10128 (
            .O(N__46659),
            .I(N__46653));
    Odrv4 I__10127 (
            .O(N__46656),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    LocalMux I__10126 (
            .O(N__46653),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ));
    InMux I__10125 (
            .O(N__46648),
            .I(N__46644));
    InMux I__10124 (
            .O(N__46647),
            .I(N__46641));
    LocalMux I__10123 (
            .O(N__46644),
            .I(N__46638));
    LocalMux I__10122 (
            .O(N__46641),
            .I(N__46635));
    Span4Mux_h I__10121 (
            .O(N__46638),
            .I(N__46632));
    Odrv4 I__10120 (
            .O(N__46635),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    Odrv4 I__10119 (
            .O(N__46632),
            .I(elapsed_time_ns_1_RNIDV2T9_0_1));
    InMux I__10118 (
            .O(N__46627),
            .I(N__46624));
    LocalMux I__10117 (
            .O(N__46624),
            .I(N__46620));
    InMux I__10116 (
            .O(N__46623),
            .I(N__46617));
    Odrv4 I__10115 (
            .O(N__46620),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    LocalMux I__10114 (
            .O(N__46617),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ));
    InMux I__10113 (
            .O(N__46612),
            .I(N__46608));
    InMux I__10112 (
            .O(N__46611),
            .I(N__46605));
    LocalMux I__10111 (
            .O(N__46608),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    LocalMux I__10110 (
            .O(N__46605),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ));
    InMux I__10109 (
            .O(N__46600),
            .I(N__46596));
    CascadeMux I__10108 (
            .O(N__46599),
            .I(N__46593));
    LocalMux I__10107 (
            .O(N__46596),
            .I(N__46590));
    InMux I__10106 (
            .O(N__46593),
            .I(N__46587));
    Span4Mux_v I__10105 (
            .O(N__46590),
            .I(N__46584));
    LocalMux I__10104 (
            .O(N__46587),
            .I(N__46581));
    Odrv4 I__10103 (
            .O(N__46584),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    Odrv4 I__10102 (
            .O(N__46581),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ));
    InMux I__10101 (
            .O(N__46576),
            .I(N__46573));
    LocalMux I__10100 (
            .O(N__46573),
            .I(N__46570));
    Span4Mux_h I__10099 (
            .O(N__46570),
            .I(N__46566));
    InMux I__10098 (
            .O(N__46569),
            .I(N__46563));
    Odrv4 I__10097 (
            .O(N__46566),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    LocalMux I__10096 (
            .O(N__46563),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ));
    InMux I__10095 (
            .O(N__46558),
            .I(N__46554));
    InMux I__10094 (
            .O(N__46557),
            .I(N__46551));
    LocalMux I__10093 (
            .O(N__46554),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    LocalMux I__10092 (
            .O(N__46551),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ));
    InMux I__10091 (
            .O(N__46546),
            .I(N__46543));
    LocalMux I__10090 (
            .O(N__46543),
            .I(elapsed_time_ns_1_RNI57CN9_0_18));
    CascadeMux I__10089 (
            .O(N__46540),
            .I(elapsed_time_ns_1_RNI57CN9_0_18_cascade_));
    InMux I__10088 (
            .O(N__46537),
            .I(N__46534));
    LocalMux I__10087 (
            .O(N__46534),
            .I(N__46531));
    Span4Mux_v I__10086 (
            .O(N__46531),
            .I(N__46528));
    Odrv4 I__10085 (
            .O(N__46528),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ));
    InMux I__10084 (
            .O(N__46525),
            .I(N__46509));
    InMux I__10083 (
            .O(N__46524),
            .I(N__46509));
    InMux I__10082 (
            .O(N__46523),
            .I(N__46509));
    InMux I__10081 (
            .O(N__46522),
            .I(N__46509));
    InMux I__10080 (
            .O(N__46521),
            .I(N__46490));
    InMux I__10079 (
            .O(N__46520),
            .I(N__46490));
    InMux I__10078 (
            .O(N__46519),
            .I(N__46490));
    InMux I__10077 (
            .O(N__46518),
            .I(N__46490));
    LocalMux I__10076 (
            .O(N__46509),
            .I(N__46487));
    InMux I__10075 (
            .O(N__46508),
            .I(N__46478));
    InMux I__10074 (
            .O(N__46507),
            .I(N__46478));
    InMux I__10073 (
            .O(N__46506),
            .I(N__46478));
    InMux I__10072 (
            .O(N__46505),
            .I(N__46478));
    InMux I__10071 (
            .O(N__46504),
            .I(N__46469));
    InMux I__10070 (
            .O(N__46503),
            .I(N__46469));
    InMux I__10069 (
            .O(N__46502),
            .I(N__46469));
    InMux I__10068 (
            .O(N__46501),
            .I(N__46469));
    InMux I__10067 (
            .O(N__46500),
            .I(N__46452));
    InMux I__10066 (
            .O(N__46499),
            .I(N__46452));
    LocalMux I__10065 (
            .O(N__46490),
            .I(N__46443));
    Span4Mux_h I__10064 (
            .O(N__46487),
            .I(N__46443));
    LocalMux I__10063 (
            .O(N__46478),
            .I(N__46443));
    LocalMux I__10062 (
            .O(N__46469),
            .I(N__46443));
    InMux I__10061 (
            .O(N__46468),
            .I(N__46434));
    InMux I__10060 (
            .O(N__46467),
            .I(N__46434));
    InMux I__10059 (
            .O(N__46466),
            .I(N__46434));
    InMux I__10058 (
            .O(N__46465),
            .I(N__46434));
    InMux I__10057 (
            .O(N__46464),
            .I(N__46425));
    InMux I__10056 (
            .O(N__46463),
            .I(N__46425));
    InMux I__10055 (
            .O(N__46462),
            .I(N__46425));
    InMux I__10054 (
            .O(N__46461),
            .I(N__46425));
    InMux I__10053 (
            .O(N__46460),
            .I(N__46416));
    InMux I__10052 (
            .O(N__46459),
            .I(N__46416));
    InMux I__10051 (
            .O(N__46458),
            .I(N__46416));
    InMux I__10050 (
            .O(N__46457),
            .I(N__46416));
    LocalMux I__10049 (
            .O(N__46452),
            .I(N__46413));
    Span4Mux_v I__10048 (
            .O(N__46443),
            .I(N__46410));
    LocalMux I__10047 (
            .O(N__46434),
            .I(N__46403));
    LocalMux I__10046 (
            .O(N__46425),
            .I(N__46403));
    LocalMux I__10045 (
            .O(N__46416),
            .I(N__46403));
    Odrv4 I__10044 (
            .O(N__46413),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv4 I__10043 (
            .O(N__46410),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    Odrv12 I__10042 (
            .O(N__46403),
            .I(\delay_measurement_inst.delay_hc_timer.running_i ));
    CascadeMux I__10041 (
            .O(N__46396),
            .I(N__46393));
    InMux I__10040 (
            .O(N__46393),
            .I(N__46389));
    InMux I__10039 (
            .O(N__46392),
            .I(N__46386));
    LocalMux I__10038 (
            .O(N__46389),
            .I(N__46380));
    LocalMux I__10037 (
            .O(N__46386),
            .I(N__46380));
    InMux I__10036 (
            .O(N__46385),
            .I(N__46377));
    Span4Mux_h I__10035 (
            .O(N__46380),
            .I(N__46374));
    LocalMux I__10034 (
            .O(N__46377),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    Odrv4 I__10033 (
            .O(N__46374),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ));
    InMux I__10032 (
            .O(N__46369),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ));
    CascadeMux I__10031 (
            .O(N__46366),
            .I(N__46363));
    InMux I__10030 (
            .O(N__46363),
            .I(N__46359));
    InMux I__10029 (
            .O(N__46362),
            .I(N__46356));
    LocalMux I__10028 (
            .O(N__46359),
            .I(N__46350));
    LocalMux I__10027 (
            .O(N__46356),
            .I(N__46350));
    InMux I__10026 (
            .O(N__46355),
            .I(N__46347));
    Span4Mux_h I__10025 (
            .O(N__46350),
            .I(N__46344));
    LocalMux I__10024 (
            .O(N__46347),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    Odrv4 I__10023 (
            .O(N__46344),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ));
    InMux I__10022 (
            .O(N__46339),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ));
    InMux I__10021 (
            .O(N__46336),
            .I(N__46333));
    LocalMux I__10020 (
            .O(N__46333),
            .I(N__46329));
    InMux I__10019 (
            .O(N__46332),
            .I(N__46326));
    Span4Mux_h I__10018 (
            .O(N__46329),
            .I(N__46323));
    LocalMux I__10017 (
            .O(N__46326),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    Odrv4 I__10016 (
            .O(N__46323),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ));
    InMux I__10015 (
            .O(N__46318),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ));
    InMux I__10014 (
            .O(N__46315),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ));
    InMux I__10013 (
            .O(N__46312),
            .I(N__46308));
    InMux I__10012 (
            .O(N__46311),
            .I(N__46305));
    LocalMux I__10011 (
            .O(N__46308),
            .I(N__46302));
    LocalMux I__10010 (
            .O(N__46305),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    Odrv4 I__10009 (
            .O(N__46302),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ));
    InMux I__10008 (
            .O(N__46297),
            .I(N__46294));
    LocalMux I__10007 (
            .O(N__46294),
            .I(N__46291));
    Span4Mux_v I__10006 (
            .O(N__46291),
            .I(N__46287));
    InMux I__10005 (
            .O(N__46290),
            .I(N__46284));
    Odrv4 I__10004 (
            .O(N__46287),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    LocalMux I__10003 (
            .O(N__46284),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ));
    InMux I__10002 (
            .O(N__46279),
            .I(N__46276));
    LocalMux I__10001 (
            .O(N__46276),
            .I(N__46272));
    InMux I__10000 (
            .O(N__46275),
            .I(N__46269));
    Odrv4 I__9999 (
            .O(N__46272),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    LocalMux I__9998 (
            .O(N__46269),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ));
    InMux I__9997 (
            .O(N__46264),
            .I(N__46260));
    CascadeMux I__9996 (
            .O(N__46263),
            .I(N__46257));
    LocalMux I__9995 (
            .O(N__46260),
            .I(N__46254));
    InMux I__9994 (
            .O(N__46257),
            .I(N__46251));
    Odrv4 I__9993 (
            .O(N__46254),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    LocalMux I__9992 (
            .O(N__46251),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ));
    InMux I__9991 (
            .O(N__46246),
            .I(N__46243));
    LocalMux I__9990 (
            .O(N__46243),
            .I(elapsed_time_ns_1_RNI69DN9_0_28));
    CascadeMux I__9989 (
            .O(N__46240),
            .I(elapsed_time_ns_1_RNI69DN9_0_28_cascade_));
    InMux I__9988 (
            .O(N__46237),
            .I(N__46234));
    LocalMux I__9987 (
            .O(N__46234),
            .I(N__46231));
    Odrv12 I__9986 (
            .O(N__46231),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ));
    InMux I__9985 (
            .O(N__46228),
            .I(N__46225));
    LocalMux I__9984 (
            .O(N__46225),
            .I(N__46221));
    InMux I__9983 (
            .O(N__46224),
            .I(N__46218));
    Odrv4 I__9982 (
            .O(N__46221),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    LocalMux I__9981 (
            .O(N__46218),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ));
    InMux I__9980 (
            .O(N__46213),
            .I(N__46210));
    LocalMux I__9979 (
            .O(N__46210),
            .I(N__46206));
    InMux I__9978 (
            .O(N__46209),
            .I(N__46203));
    Odrv4 I__9977 (
            .O(N__46206),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    LocalMux I__9976 (
            .O(N__46203),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ));
    InMux I__9975 (
            .O(N__46198),
            .I(N__46194));
    CascadeMux I__9974 (
            .O(N__46197),
            .I(N__46191));
    LocalMux I__9973 (
            .O(N__46194),
            .I(N__46188));
    InMux I__9972 (
            .O(N__46191),
            .I(N__46185));
    Odrv4 I__9971 (
            .O(N__46188),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    LocalMux I__9970 (
            .O(N__46185),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ));
    InMux I__9969 (
            .O(N__46180),
            .I(N__46177));
    LocalMux I__9968 (
            .O(N__46177),
            .I(N__46173));
    InMux I__9967 (
            .O(N__46176),
            .I(N__46170));
    Odrv4 I__9966 (
            .O(N__46173),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    LocalMux I__9965 (
            .O(N__46170),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ));
    InMux I__9964 (
            .O(N__46165),
            .I(N__46159));
    InMux I__9963 (
            .O(N__46164),
            .I(N__46159));
    LocalMux I__9962 (
            .O(N__46159),
            .I(N__46155));
    InMux I__9961 (
            .O(N__46158),
            .I(N__46152));
    Span4Mux_h I__9960 (
            .O(N__46155),
            .I(N__46149));
    LocalMux I__9959 (
            .O(N__46152),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    Odrv4 I__9958 (
            .O(N__46149),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ));
    InMux I__9957 (
            .O(N__46144),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ));
    InMux I__9956 (
            .O(N__46141),
            .I(N__46134));
    InMux I__9955 (
            .O(N__46140),
            .I(N__46134));
    InMux I__9954 (
            .O(N__46139),
            .I(N__46131));
    LocalMux I__9953 (
            .O(N__46134),
            .I(N__46128));
    LocalMux I__9952 (
            .O(N__46131),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    Odrv4 I__9951 (
            .O(N__46128),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ));
    InMux I__9950 (
            .O(N__46123),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ));
    CascadeMux I__9949 (
            .O(N__46120),
            .I(N__46116));
    CascadeMux I__9948 (
            .O(N__46119),
            .I(N__46113));
    InMux I__9947 (
            .O(N__46116),
            .I(N__46107));
    InMux I__9946 (
            .O(N__46113),
            .I(N__46107));
    InMux I__9945 (
            .O(N__46112),
            .I(N__46104));
    LocalMux I__9944 (
            .O(N__46107),
            .I(N__46101));
    LocalMux I__9943 (
            .O(N__46104),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    Odrv4 I__9942 (
            .O(N__46101),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ));
    InMux I__9941 (
            .O(N__46096),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ));
    CascadeMux I__9940 (
            .O(N__46093),
            .I(N__46090));
    InMux I__9939 (
            .O(N__46090),
            .I(N__46086));
    InMux I__9938 (
            .O(N__46089),
            .I(N__46082));
    LocalMux I__9937 (
            .O(N__46086),
            .I(N__46079));
    InMux I__9936 (
            .O(N__46085),
            .I(N__46076));
    LocalMux I__9935 (
            .O(N__46082),
            .I(N__46071));
    Span4Mux_h I__9934 (
            .O(N__46079),
            .I(N__46071));
    LocalMux I__9933 (
            .O(N__46076),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    Odrv4 I__9932 (
            .O(N__46071),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ));
    InMux I__9931 (
            .O(N__46066),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ));
    InMux I__9930 (
            .O(N__46063),
            .I(N__46056));
    InMux I__9929 (
            .O(N__46062),
            .I(N__46056));
    InMux I__9928 (
            .O(N__46061),
            .I(N__46053));
    LocalMux I__9927 (
            .O(N__46056),
            .I(N__46050));
    LocalMux I__9926 (
            .O(N__46053),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    Odrv4 I__9925 (
            .O(N__46050),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ));
    InMux I__9924 (
            .O(N__46045),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ));
    CascadeMux I__9923 (
            .O(N__46042),
            .I(N__46038));
    CascadeMux I__9922 (
            .O(N__46041),
            .I(N__46035));
    InMux I__9921 (
            .O(N__46038),
            .I(N__46029));
    InMux I__9920 (
            .O(N__46035),
            .I(N__46029));
    InMux I__9919 (
            .O(N__46034),
            .I(N__46026));
    LocalMux I__9918 (
            .O(N__46029),
            .I(N__46023));
    LocalMux I__9917 (
            .O(N__46026),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    Odrv4 I__9916 (
            .O(N__46023),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ));
    InMux I__9915 (
            .O(N__46018),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ));
    CascadeMux I__9914 (
            .O(N__46015),
            .I(N__46012));
    InMux I__9913 (
            .O(N__46012),
            .I(N__46007));
    CascadeMux I__9912 (
            .O(N__46011),
            .I(N__46004));
    InMux I__9911 (
            .O(N__46010),
            .I(N__46001));
    LocalMux I__9910 (
            .O(N__46007),
            .I(N__45998));
    InMux I__9909 (
            .O(N__46004),
            .I(N__45995));
    LocalMux I__9908 (
            .O(N__46001),
            .I(N__45990));
    Span4Mux_v I__9907 (
            .O(N__45998),
            .I(N__45990));
    LocalMux I__9906 (
            .O(N__45995),
            .I(N__45987));
    Odrv4 I__9905 (
            .O(N__45990),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    Odrv4 I__9904 (
            .O(N__45987),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ));
    InMux I__9903 (
            .O(N__45982),
            .I(bfn_18_10_0_));
    CascadeMux I__9902 (
            .O(N__45979),
            .I(N__45976));
    InMux I__9901 (
            .O(N__45976),
            .I(N__45973));
    LocalMux I__9900 (
            .O(N__45973),
            .I(N__45968));
    InMux I__9899 (
            .O(N__45972),
            .I(N__45965));
    InMux I__9898 (
            .O(N__45971),
            .I(N__45962));
    Span4Mux_v I__9897 (
            .O(N__45968),
            .I(N__45959));
    LocalMux I__9896 (
            .O(N__45965),
            .I(N__45956));
    LocalMux I__9895 (
            .O(N__45962),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__9894 (
            .O(N__45959),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    Odrv4 I__9893 (
            .O(N__45956),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ));
    InMux I__9892 (
            .O(N__45949),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ));
    CascadeMux I__9891 (
            .O(N__45946),
            .I(N__45943));
    InMux I__9890 (
            .O(N__45943),
            .I(N__45938));
    InMux I__9889 (
            .O(N__45942),
            .I(N__45935));
    InMux I__9888 (
            .O(N__45941),
            .I(N__45932));
    LocalMux I__9887 (
            .O(N__45938),
            .I(N__45929));
    LocalMux I__9886 (
            .O(N__45935),
            .I(N__45926));
    LocalMux I__9885 (
            .O(N__45932),
            .I(N__45921));
    Span4Mux_v I__9884 (
            .O(N__45929),
            .I(N__45921));
    Span4Mux_h I__9883 (
            .O(N__45926),
            .I(N__45918));
    Odrv4 I__9882 (
            .O(N__45921),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    Odrv4 I__9881 (
            .O(N__45918),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ));
    InMux I__9880 (
            .O(N__45913),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ));
    CascadeMux I__9879 (
            .O(N__45910),
            .I(N__45906));
    CascadeMux I__9878 (
            .O(N__45909),
            .I(N__45903));
    InMux I__9877 (
            .O(N__45906),
            .I(N__45897));
    InMux I__9876 (
            .O(N__45903),
            .I(N__45897));
    InMux I__9875 (
            .O(N__45902),
            .I(N__45894));
    LocalMux I__9874 (
            .O(N__45897),
            .I(N__45891));
    LocalMux I__9873 (
            .O(N__45894),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    Odrv4 I__9872 (
            .O(N__45891),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ));
    InMux I__9871 (
            .O(N__45886),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ));
    InMux I__9870 (
            .O(N__45883),
            .I(N__45877));
    InMux I__9869 (
            .O(N__45882),
            .I(N__45877));
    LocalMux I__9868 (
            .O(N__45877),
            .I(N__45873));
    InMux I__9867 (
            .O(N__45876),
            .I(N__45870));
    Span4Mux_h I__9866 (
            .O(N__45873),
            .I(N__45867));
    LocalMux I__9865 (
            .O(N__45870),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    Odrv4 I__9864 (
            .O(N__45867),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ));
    InMux I__9863 (
            .O(N__45862),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ));
    CascadeMux I__9862 (
            .O(N__45859),
            .I(N__45856));
    InMux I__9861 (
            .O(N__45856),
            .I(N__45852));
    InMux I__9860 (
            .O(N__45855),
            .I(N__45849));
    LocalMux I__9859 (
            .O(N__45852),
            .I(N__45843));
    LocalMux I__9858 (
            .O(N__45849),
            .I(N__45843));
    InMux I__9857 (
            .O(N__45848),
            .I(N__45840));
    Span4Mux_h I__9856 (
            .O(N__45843),
            .I(N__45837));
    LocalMux I__9855 (
            .O(N__45840),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    Odrv4 I__9854 (
            .O(N__45837),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ));
    InMux I__9853 (
            .O(N__45832),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ));
    CascadeMux I__9852 (
            .O(N__45829),
            .I(N__45826));
    InMux I__9851 (
            .O(N__45826),
            .I(N__45822));
    InMux I__9850 (
            .O(N__45825),
            .I(N__45818));
    LocalMux I__9849 (
            .O(N__45822),
            .I(N__45815));
    InMux I__9848 (
            .O(N__45821),
            .I(N__45812));
    LocalMux I__9847 (
            .O(N__45818),
            .I(N__45807));
    Span4Mux_h I__9846 (
            .O(N__45815),
            .I(N__45807));
    LocalMux I__9845 (
            .O(N__45812),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    Odrv4 I__9844 (
            .O(N__45807),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ));
    InMux I__9843 (
            .O(N__45802),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ));
    InMux I__9842 (
            .O(N__45799),
            .I(N__45792));
    InMux I__9841 (
            .O(N__45798),
            .I(N__45792));
    InMux I__9840 (
            .O(N__45797),
            .I(N__45789));
    LocalMux I__9839 (
            .O(N__45792),
            .I(N__45786));
    LocalMux I__9838 (
            .O(N__45789),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    Odrv4 I__9837 (
            .O(N__45786),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ));
    InMux I__9836 (
            .O(N__45781),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ));
    CascadeMux I__9835 (
            .O(N__45778),
            .I(N__45774));
    CascadeMux I__9834 (
            .O(N__45777),
            .I(N__45771));
    InMux I__9833 (
            .O(N__45774),
            .I(N__45765));
    InMux I__9832 (
            .O(N__45771),
            .I(N__45765));
    InMux I__9831 (
            .O(N__45770),
            .I(N__45762));
    LocalMux I__9830 (
            .O(N__45765),
            .I(N__45759));
    LocalMux I__9829 (
            .O(N__45762),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    Odrv4 I__9828 (
            .O(N__45759),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ));
    InMux I__9827 (
            .O(N__45754),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ));
    CascadeMux I__9826 (
            .O(N__45751),
            .I(N__45748));
    InMux I__9825 (
            .O(N__45748),
            .I(N__45744));
    CascadeMux I__9824 (
            .O(N__45747),
            .I(N__45741));
    LocalMux I__9823 (
            .O(N__45744),
            .I(N__45737));
    InMux I__9822 (
            .O(N__45741),
            .I(N__45734));
    InMux I__9821 (
            .O(N__45740),
            .I(N__45731));
    Span4Mux_v I__9820 (
            .O(N__45737),
            .I(N__45726));
    LocalMux I__9819 (
            .O(N__45734),
            .I(N__45726));
    LocalMux I__9818 (
            .O(N__45731),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    Odrv4 I__9817 (
            .O(N__45726),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ));
    InMux I__9816 (
            .O(N__45721),
            .I(bfn_18_9_0_));
    CascadeMux I__9815 (
            .O(N__45718),
            .I(N__45715));
    InMux I__9814 (
            .O(N__45715),
            .I(N__45712));
    LocalMux I__9813 (
            .O(N__45712),
            .I(N__45707));
    InMux I__9812 (
            .O(N__45711),
            .I(N__45704));
    InMux I__9811 (
            .O(N__45710),
            .I(N__45701));
    Span4Mux_v I__9810 (
            .O(N__45707),
            .I(N__45698));
    LocalMux I__9809 (
            .O(N__45704),
            .I(N__45695));
    LocalMux I__9808 (
            .O(N__45701),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__9807 (
            .O(N__45698),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    Odrv4 I__9806 (
            .O(N__45695),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ));
    InMux I__9805 (
            .O(N__45688),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ));
    InMux I__9804 (
            .O(N__45685),
            .I(N__45681));
    CascadeMux I__9803 (
            .O(N__45684),
            .I(N__45678));
    LocalMux I__9802 (
            .O(N__45681),
            .I(N__45674));
    InMux I__9801 (
            .O(N__45678),
            .I(N__45671));
    InMux I__9800 (
            .O(N__45677),
            .I(N__45668));
    Span4Mux_h I__9799 (
            .O(N__45674),
            .I(N__45663));
    LocalMux I__9798 (
            .O(N__45671),
            .I(N__45663));
    LocalMux I__9797 (
            .O(N__45668),
            .I(N__45658));
    Span4Mux_v I__9796 (
            .O(N__45663),
            .I(N__45658));
    Odrv4 I__9795 (
            .O(N__45658),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ));
    InMux I__9794 (
            .O(N__45655),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ));
    CascadeMux I__9793 (
            .O(N__45652),
            .I(N__45648));
    CascadeMux I__9792 (
            .O(N__45651),
            .I(N__45645));
    InMux I__9791 (
            .O(N__45648),
            .I(N__45639));
    InMux I__9790 (
            .O(N__45645),
            .I(N__45639));
    InMux I__9789 (
            .O(N__45644),
            .I(N__45636));
    LocalMux I__9788 (
            .O(N__45639),
            .I(N__45633));
    LocalMux I__9787 (
            .O(N__45636),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    Odrv4 I__9786 (
            .O(N__45633),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ));
    InMux I__9785 (
            .O(N__45628),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ));
    InMux I__9784 (
            .O(N__45625),
            .I(N__45618));
    InMux I__9783 (
            .O(N__45624),
            .I(N__45618));
    InMux I__9782 (
            .O(N__45623),
            .I(N__45615));
    LocalMux I__9781 (
            .O(N__45618),
            .I(N__45612));
    LocalMux I__9780 (
            .O(N__45615),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    Odrv4 I__9779 (
            .O(N__45612),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ));
    InMux I__9778 (
            .O(N__45607),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ));
    CascadeMux I__9777 (
            .O(N__45604),
            .I(N__45600));
    InMux I__9776 (
            .O(N__45603),
            .I(N__45597));
    InMux I__9775 (
            .O(N__45600),
            .I(N__45593));
    LocalMux I__9774 (
            .O(N__45597),
            .I(N__45590));
    InMux I__9773 (
            .O(N__45596),
            .I(N__45587));
    LocalMux I__9772 (
            .O(N__45593),
            .I(N__45582));
    Span4Mux_h I__9771 (
            .O(N__45590),
            .I(N__45582));
    LocalMux I__9770 (
            .O(N__45587),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    Odrv4 I__9769 (
            .O(N__45582),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ));
    InMux I__9768 (
            .O(N__45577),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ));
    CascadeMux I__9767 (
            .O(N__45574),
            .I(N__45570));
    CascadeMux I__9766 (
            .O(N__45573),
            .I(N__45567));
    InMux I__9765 (
            .O(N__45570),
            .I(N__45562));
    InMux I__9764 (
            .O(N__45567),
            .I(N__45562));
    LocalMux I__9763 (
            .O(N__45562),
            .I(N__45558));
    InMux I__9762 (
            .O(N__45561),
            .I(N__45555));
    Span4Mux_h I__9761 (
            .O(N__45558),
            .I(N__45552));
    LocalMux I__9760 (
            .O(N__45555),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    Odrv4 I__9759 (
            .O(N__45552),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ));
    InMux I__9758 (
            .O(N__45547),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ));
    InMux I__9757 (
            .O(N__45544),
            .I(N__45537));
    InMux I__9756 (
            .O(N__45543),
            .I(N__45537));
    InMux I__9755 (
            .O(N__45542),
            .I(N__45534));
    LocalMux I__9754 (
            .O(N__45537),
            .I(N__45531));
    LocalMux I__9753 (
            .O(N__45534),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    Odrv4 I__9752 (
            .O(N__45531),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ));
    InMux I__9751 (
            .O(N__45526),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ));
    CascadeMux I__9750 (
            .O(N__45523),
            .I(N__45520));
    InMux I__9749 (
            .O(N__45520),
            .I(N__45516));
    InMux I__9748 (
            .O(N__45519),
            .I(N__45513));
    LocalMux I__9747 (
            .O(N__45516),
            .I(N__45507));
    LocalMux I__9746 (
            .O(N__45513),
            .I(N__45507));
    InMux I__9745 (
            .O(N__45512),
            .I(N__45504));
    Span4Mux_h I__9744 (
            .O(N__45507),
            .I(N__45501));
    LocalMux I__9743 (
            .O(N__45504),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    Odrv4 I__9742 (
            .O(N__45501),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ));
    InMux I__9741 (
            .O(N__45496),
            .I(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ));
    InMux I__9740 (
            .O(N__45493),
            .I(N__45489));
    CascadeMux I__9739 (
            .O(N__45492),
            .I(N__45486));
    LocalMux I__9738 (
            .O(N__45489),
            .I(N__45482));
    InMux I__9737 (
            .O(N__45486),
            .I(N__45479));
    InMux I__9736 (
            .O(N__45485),
            .I(N__45476));
    Span4Mux_v I__9735 (
            .O(N__45482),
            .I(N__45471));
    LocalMux I__9734 (
            .O(N__45479),
            .I(N__45471));
    LocalMux I__9733 (
            .O(N__45476),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    Odrv4 I__9732 (
            .O(N__45471),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ));
    InMux I__9731 (
            .O(N__45466),
            .I(bfn_18_8_0_));
    CascadeMux I__9730 (
            .O(N__45463),
            .I(N__45460));
    InMux I__9729 (
            .O(N__45460),
            .I(N__45457));
    LocalMux I__9728 (
            .O(N__45457),
            .I(N__45454));
    Odrv4 I__9727 (
            .O(N__45454),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ));
    InMux I__9726 (
            .O(N__45451),
            .I(N__45448));
    LocalMux I__9725 (
            .O(N__45448),
            .I(N__45445));
    Span4Mux_h I__9724 (
            .O(N__45445),
            .I(N__45442));
    Odrv4 I__9723 (
            .O(N__45442),
            .I(\current_shift_inst.un38_control_input_0_s0_28 ));
    InMux I__9722 (
            .O(N__45439),
            .I(\current_shift_inst.un38_control_input_cry_27_s0 ));
    InMux I__9721 (
            .O(N__45436),
            .I(N__45433));
    LocalMux I__9720 (
            .O(N__45433),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ));
    InMux I__9719 (
            .O(N__45430),
            .I(N__45427));
    LocalMux I__9718 (
            .O(N__45427),
            .I(N__45424));
    Odrv12 I__9717 (
            .O(N__45424),
            .I(\current_shift_inst.un38_control_input_0_s0_29 ));
    InMux I__9716 (
            .O(N__45421),
            .I(\current_shift_inst.un38_control_input_cry_28_s0 ));
    CascadeMux I__9715 (
            .O(N__45418),
            .I(N__45415));
    InMux I__9714 (
            .O(N__45415),
            .I(N__45412));
    LocalMux I__9713 (
            .O(N__45412),
            .I(N__45409));
    Span4Mux_h I__9712 (
            .O(N__45409),
            .I(N__45406));
    Span4Mux_v I__9711 (
            .O(N__45406),
            .I(N__45403));
    Span4Mux_v I__9710 (
            .O(N__45403),
            .I(N__45400));
    Odrv4 I__9709 (
            .O(N__45400),
            .I(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ));
    InMux I__9708 (
            .O(N__45397),
            .I(N__45394));
    LocalMux I__9707 (
            .O(N__45394),
            .I(N__45391));
    Odrv4 I__9706 (
            .O(N__45391),
            .I(\current_shift_inst.un38_control_input_0_s0_30 ));
    InMux I__9705 (
            .O(N__45388),
            .I(\current_shift_inst.un38_control_input_cry_29_s0 ));
    InMux I__9704 (
            .O(N__45385),
            .I(N__45382));
    LocalMux I__9703 (
            .O(N__45382),
            .I(N__45379));
    Span4Mux_v I__9702 (
            .O(N__45379),
            .I(N__45376));
    Span4Mux_v I__9701 (
            .O(N__45376),
            .I(N__45373));
    Odrv4 I__9700 (
            .O(N__45373),
            .I(\current_shift_inst.un38_control_input_axb_31_s0 ));
    InMux I__9699 (
            .O(N__45370),
            .I(\current_shift_inst.un38_control_input_cry_30_s0 ));
    InMux I__9698 (
            .O(N__45367),
            .I(N__45364));
    LocalMux I__9697 (
            .O(N__45364),
            .I(N__45361));
    Span4Mux_h I__9696 (
            .O(N__45361),
            .I(N__45358));
    Odrv4 I__9695 (
            .O(N__45358),
            .I(\current_shift_inst.control_input_axb_28 ));
    InMux I__9694 (
            .O(N__45355),
            .I(N__45352));
    LocalMux I__9693 (
            .O(N__45352),
            .I(elapsed_time_ns_1_RNI58DN9_0_27));
    CascadeMux I__9692 (
            .O(N__45349),
            .I(elapsed_time_ns_1_RNI58DN9_0_27_cascade_));
    InMux I__9691 (
            .O(N__45346),
            .I(N__45343));
    LocalMux I__9690 (
            .O(N__45343),
            .I(N__45340));
    Span4Mux_h I__9689 (
            .O(N__45340),
            .I(N__45337));
    Span4Mux_v I__9688 (
            .O(N__45337),
            .I(N__45334));
    Odrv4 I__9687 (
            .O(N__45334),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ));
    InMux I__9686 (
            .O(N__45331),
            .I(N__45327));
    InMux I__9685 (
            .O(N__45330),
            .I(N__45324));
    LocalMux I__9684 (
            .O(N__45327),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    LocalMux I__9683 (
            .O(N__45324),
            .I(elapsed_time_ns_1_RNI46CN9_0_17));
    InMux I__9682 (
            .O(N__45319),
            .I(N__45316));
    LocalMux I__9681 (
            .O(N__45316),
            .I(N__45312));
    InMux I__9680 (
            .O(N__45315),
            .I(N__45309));
    Span4Mux_h I__9679 (
            .O(N__45312),
            .I(N__45304));
    LocalMux I__9678 (
            .O(N__45309),
            .I(N__45304));
    Span4Mux_v I__9677 (
            .O(N__45304),
            .I(N__45300));
    InMux I__9676 (
            .O(N__45303),
            .I(N__45297));
    Odrv4 I__9675 (
            .O(N__45300),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    LocalMux I__9674 (
            .O(N__45297),
            .I(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ));
    InMux I__9673 (
            .O(N__45292),
            .I(bfn_18_7_0_));
    CascadeMux I__9672 (
            .O(N__45289),
            .I(N__45286));
    InMux I__9671 (
            .O(N__45286),
            .I(N__45283));
    LocalMux I__9670 (
            .O(N__45283),
            .I(N__45280));
    Odrv12 I__9669 (
            .O(N__45280),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ));
    InMux I__9668 (
            .O(N__45277),
            .I(N__45274));
    LocalMux I__9667 (
            .O(N__45274),
            .I(N__45271));
    Span4Mux_v I__9666 (
            .O(N__45271),
            .I(N__45268));
    Sp12to4 I__9665 (
            .O(N__45268),
            .I(N__45265));
    Odrv12 I__9664 (
            .O(N__45265),
            .I(\current_shift_inst.un38_control_input_0_s0_20 ));
    InMux I__9663 (
            .O(N__45262),
            .I(\current_shift_inst.un38_control_input_cry_19_s0 ));
    InMux I__9662 (
            .O(N__45259),
            .I(N__45256));
    LocalMux I__9661 (
            .O(N__45256),
            .I(N__45253));
    Odrv12 I__9660 (
            .O(N__45253),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ));
    InMux I__9659 (
            .O(N__45250),
            .I(N__45247));
    LocalMux I__9658 (
            .O(N__45247),
            .I(N__45244));
    Span4Mux_v I__9657 (
            .O(N__45244),
            .I(N__45241));
    Sp12to4 I__9656 (
            .O(N__45241),
            .I(N__45238));
    Odrv12 I__9655 (
            .O(N__45238),
            .I(\current_shift_inst.un38_control_input_0_s0_21 ));
    InMux I__9654 (
            .O(N__45235),
            .I(\current_shift_inst.un38_control_input_cry_20_s0 ));
    CascadeMux I__9653 (
            .O(N__45232),
            .I(N__45229));
    InMux I__9652 (
            .O(N__45229),
            .I(N__45226));
    LocalMux I__9651 (
            .O(N__45226),
            .I(N__45223));
    Span4Mux_h I__9650 (
            .O(N__45223),
            .I(N__45220));
    Span4Mux_v I__9649 (
            .O(N__45220),
            .I(N__45217));
    Odrv4 I__9648 (
            .O(N__45217),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ));
    InMux I__9647 (
            .O(N__45214),
            .I(N__45211));
    LocalMux I__9646 (
            .O(N__45211),
            .I(\current_shift_inst.un38_control_input_0_s0_22 ));
    InMux I__9645 (
            .O(N__45208),
            .I(\current_shift_inst.un38_control_input_cry_21_s0 ));
    InMux I__9644 (
            .O(N__45205),
            .I(N__45202));
    LocalMux I__9643 (
            .O(N__45202),
            .I(N__45199));
    Odrv12 I__9642 (
            .O(N__45199),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ));
    InMux I__9641 (
            .O(N__45196),
            .I(N__45193));
    LocalMux I__9640 (
            .O(N__45193),
            .I(\current_shift_inst.un38_control_input_0_s0_23 ));
    InMux I__9639 (
            .O(N__45190),
            .I(\current_shift_inst.un38_control_input_cry_22_s0 ));
    CascadeMux I__9638 (
            .O(N__45187),
            .I(N__45184));
    InMux I__9637 (
            .O(N__45184),
            .I(N__45181));
    LocalMux I__9636 (
            .O(N__45181),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ));
    InMux I__9635 (
            .O(N__45178),
            .I(N__45175));
    LocalMux I__9634 (
            .O(N__45175),
            .I(N__45172));
    Odrv4 I__9633 (
            .O(N__45172),
            .I(\current_shift_inst.un38_control_input_0_s0_24 ));
    InMux I__9632 (
            .O(N__45169),
            .I(bfn_17_21_0_));
    InMux I__9631 (
            .O(N__45166),
            .I(N__45163));
    LocalMux I__9630 (
            .O(N__45163),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ));
    InMux I__9629 (
            .O(N__45160),
            .I(N__45157));
    LocalMux I__9628 (
            .O(N__45157),
            .I(N__45154));
    Odrv4 I__9627 (
            .O(N__45154),
            .I(\current_shift_inst.un38_control_input_0_s0_25 ));
    InMux I__9626 (
            .O(N__45151),
            .I(\current_shift_inst.un38_control_input_cry_24_s0 ));
    CascadeMux I__9625 (
            .O(N__45148),
            .I(N__45145));
    InMux I__9624 (
            .O(N__45145),
            .I(N__45142));
    LocalMux I__9623 (
            .O(N__45142),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ));
    InMux I__9622 (
            .O(N__45139),
            .I(\current_shift_inst.un38_control_input_cry_25_s0 ));
    InMux I__9621 (
            .O(N__45136),
            .I(N__45133));
    LocalMux I__9620 (
            .O(N__45133),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ));
    InMux I__9619 (
            .O(N__45130),
            .I(N__45127));
    LocalMux I__9618 (
            .O(N__45127),
            .I(\current_shift_inst.un38_control_input_0_s0_27 ));
    InMux I__9617 (
            .O(N__45124),
            .I(\current_shift_inst.un38_control_input_cry_26_s0 ));
    CascadeMux I__9616 (
            .O(N__45121),
            .I(N__45118));
    InMux I__9615 (
            .O(N__45118),
            .I(N__45115));
    LocalMux I__9614 (
            .O(N__45115),
            .I(N__45112));
    Odrv12 I__9613 (
            .O(N__45112),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ));
    InMux I__9612 (
            .O(N__45109),
            .I(N__45106));
    LocalMux I__9611 (
            .O(N__45106),
            .I(\current_shift_inst.un38_control_input_0_s0_12 ));
    InMux I__9610 (
            .O(N__45103),
            .I(\current_shift_inst.un38_control_input_cry_11_s0 ));
    InMux I__9609 (
            .O(N__45100),
            .I(N__45097));
    LocalMux I__9608 (
            .O(N__45097),
            .I(N__45094));
    Odrv4 I__9607 (
            .O(N__45094),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ));
    InMux I__9606 (
            .O(N__45091),
            .I(N__45088));
    LocalMux I__9605 (
            .O(N__45088),
            .I(\current_shift_inst.un38_control_input_0_s0_13 ));
    InMux I__9604 (
            .O(N__45085),
            .I(\current_shift_inst.un38_control_input_cry_12_s0 ));
    CascadeMux I__9603 (
            .O(N__45082),
            .I(N__45079));
    InMux I__9602 (
            .O(N__45079),
            .I(N__45076));
    LocalMux I__9601 (
            .O(N__45076),
            .I(N__45073));
    Odrv12 I__9600 (
            .O(N__45073),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ));
    InMux I__9599 (
            .O(N__45070),
            .I(N__45067));
    LocalMux I__9598 (
            .O(N__45067),
            .I(\current_shift_inst.un38_control_input_0_s0_14 ));
    InMux I__9597 (
            .O(N__45064),
            .I(\current_shift_inst.un38_control_input_cry_13_s0 ));
    InMux I__9596 (
            .O(N__45061),
            .I(N__45058));
    LocalMux I__9595 (
            .O(N__45058),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ));
    InMux I__9594 (
            .O(N__45055),
            .I(N__45052));
    LocalMux I__9593 (
            .O(N__45052),
            .I(\current_shift_inst.un38_control_input_0_s0_15 ));
    InMux I__9592 (
            .O(N__45049),
            .I(\current_shift_inst.un38_control_input_cry_14_s0 ));
    CascadeMux I__9591 (
            .O(N__45046),
            .I(N__45043));
    InMux I__9590 (
            .O(N__45043),
            .I(N__45040));
    LocalMux I__9589 (
            .O(N__45040),
            .I(N__45037));
    Odrv12 I__9588 (
            .O(N__45037),
            .I(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ));
    InMux I__9587 (
            .O(N__45034),
            .I(N__45031));
    LocalMux I__9586 (
            .O(N__45031),
            .I(N__45028));
    Odrv4 I__9585 (
            .O(N__45028),
            .I(\current_shift_inst.un38_control_input_0_s0_16 ));
    InMux I__9584 (
            .O(N__45025),
            .I(bfn_17_20_0_));
    InMux I__9583 (
            .O(N__45022),
            .I(N__45019));
    LocalMux I__9582 (
            .O(N__45019),
            .I(N__45016));
    Span4Mux_v I__9581 (
            .O(N__45016),
            .I(N__45013));
    Odrv4 I__9580 (
            .O(N__45013),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ));
    InMux I__9579 (
            .O(N__45010),
            .I(N__45007));
    LocalMux I__9578 (
            .O(N__45007),
            .I(\current_shift_inst.un38_control_input_0_s0_17 ));
    InMux I__9577 (
            .O(N__45004),
            .I(\current_shift_inst.un38_control_input_cry_16_s0 ));
    CascadeMux I__9576 (
            .O(N__45001),
            .I(N__44998));
    InMux I__9575 (
            .O(N__44998),
            .I(N__44995));
    LocalMux I__9574 (
            .O(N__44995),
            .I(N__44992));
    Span12Mux_s9_h I__9573 (
            .O(N__44992),
            .I(N__44989));
    Odrv12 I__9572 (
            .O(N__44989),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ));
    InMux I__9571 (
            .O(N__44986),
            .I(N__44983));
    LocalMux I__9570 (
            .O(N__44983),
            .I(\current_shift_inst.un38_control_input_0_s0_18 ));
    InMux I__9569 (
            .O(N__44980),
            .I(\current_shift_inst.un38_control_input_cry_17_s0 ));
    InMux I__9568 (
            .O(N__44977),
            .I(N__44974));
    LocalMux I__9567 (
            .O(N__44974),
            .I(N__44971));
    Odrv4 I__9566 (
            .O(N__44971),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ));
    InMux I__9565 (
            .O(N__44968),
            .I(N__44965));
    LocalMux I__9564 (
            .O(N__44965),
            .I(N__44962));
    Span4Mux_h I__9563 (
            .O(N__44962),
            .I(N__44959));
    Odrv4 I__9562 (
            .O(N__44959),
            .I(\current_shift_inst.un38_control_input_0_s0_19 ));
    InMux I__9561 (
            .O(N__44956),
            .I(\current_shift_inst.un38_control_input_cry_18_s0 ));
    CascadeMux I__9560 (
            .O(N__44953),
            .I(N__44950));
    InMux I__9559 (
            .O(N__44950),
            .I(N__44947));
    LocalMux I__9558 (
            .O(N__44947),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ));
    InMux I__9557 (
            .O(N__44944),
            .I(N__44941));
    LocalMux I__9556 (
            .O(N__44941),
            .I(N__44938));
    Span4Mux_h I__9555 (
            .O(N__44938),
            .I(N__44935));
    Odrv4 I__9554 (
            .O(N__44935),
            .I(\current_shift_inst.un38_control_input_0_s0_4 ));
    InMux I__9553 (
            .O(N__44932),
            .I(\current_shift_inst.un38_control_input_cry_3_s0 ));
    InMux I__9552 (
            .O(N__44929),
            .I(N__44926));
    LocalMux I__9551 (
            .O(N__44926),
            .I(N__44923));
    Span4Mux_v I__9550 (
            .O(N__44923),
            .I(N__44920));
    Odrv4 I__9549 (
            .O(N__44920),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ));
    InMux I__9548 (
            .O(N__44917),
            .I(N__44914));
    LocalMux I__9547 (
            .O(N__44914),
            .I(N__44911));
    Span4Mux_v I__9546 (
            .O(N__44911),
            .I(N__44908));
    Odrv4 I__9545 (
            .O(N__44908),
            .I(\current_shift_inst.un38_control_input_0_s0_5 ));
    InMux I__9544 (
            .O(N__44905),
            .I(\current_shift_inst.un38_control_input_cry_4_s0 ));
    InMux I__9543 (
            .O(N__44902),
            .I(N__44899));
    LocalMux I__9542 (
            .O(N__44899),
            .I(N__44896));
    Span4Mux_v I__9541 (
            .O(N__44896),
            .I(N__44893));
    Odrv4 I__9540 (
            .O(N__44893),
            .I(\current_shift_inst.un38_control_input_0_s0_6 ));
    InMux I__9539 (
            .O(N__44890),
            .I(\current_shift_inst.un38_control_input_cry_5_s0 ));
    InMux I__9538 (
            .O(N__44887),
            .I(N__44884));
    LocalMux I__9537 (
            .O(N__44884),
            .I(N__44881));
    Span4Mux_h I__9536 (
            .O(N__44881),
            .I(N__44878));
    Odrv4 I__9535 (
            .O(N__44878),
            .I(\current_shift_inst.un38_control_input_0_s0_7 ));
    InMux I__9534 (
            .O(N__44875),
            .I(\current_shift_inst.un38_control_input_cry_6_s0 ));
    CascadeMux I__9533 (
            .O(N__44872),
            .I(N__44869));
    InMux I__9532 (
            .O(N__44869),
            .I(N__44866));
    LocalMux I__9531 (
            .O(N__44866),
            .I(N__44863));
    Span4Mux_v I__9530 (
            .O(N__44863),
            .I(N__44860));
    Odrv4 I__9529 (
            .O(N__44860),
            .I(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ));
    InMux I__9528 (
            .O(N__44857),
            .I(N__44854));
    LocalMux I__9527 (
            .O(N__44854),
            .I(N__44851));
    Span4Mux_v I__9526 (
            .O(N__44851),
            .I(N__44848));
    Odrv4 I__9525 (
            .O(N__44848),
            .I(\current_shift_inst.un38_control_input_0_s0_8 ));
    InMux I__9524 (
            .O(N__44845),
            .I(bfn_17_19_0_));
    InMux I__9523 (
            .O(N__44842),
            .I(N__44839));
    LocalMux I__9522 (
            .O(N__44839),
            .I(N__44836));
    Odrv12 I__9521 (
            .O(N__44836),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ));
    InMux I__9520 (
            .O(N__44833),
            .I(N__44830));
    LocalMux I__9519 (
            .O(N__44830),
            .I(N__44827));
    Span4Mux_h I__9518 (
            .O(N__44827),
            .I(N__44824));
    Odrv4 I__9517 (
            .O(N__44824),
            .I(\current_shift_inst.un38_control_input_0_s0_9 ));
    InMux I__9516 (
            .O(N__44821),
            .I(\current_shift_inst.un38_control_input_cry_8_s0 ));
    CascadeMux I__9515 (
            .O(N__44818),
            .I(N__44815));
    InMux I__9514 (
            .O(N__44815),
            .I(N__44812));
    LocalMux I__9513 (
            .O(N__44812),
            .I(N__44809));
    Span4Mux_v I__9512 (
            .O(N__44809),
            .I(N__44806));
    Odrv4 I__9511 (
            .O(N__44806),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ));
    InMux I__9510 (
            .O(N__44803),
            .I(N__44800));
    LocalMux I__9509 (
            .O(N__44800),
            .I(N__44797));
    Span4Mux_v I__9508 (
            .O(N__44797),
            .I(N__44794));
    Odrv4 I__9507 (
            .O(N__44794),
            .I(\current_shift_inst.un38_control_input_0_s0_10 ));
    InMux I__9506 (
            .O(N__44791),
            .I(\current_shift_inst.un38_control_input_cry_9_s0 ));
    InMux I__9505 (
            .O(N__44788),
            .I(N__44785));
    LocalMux I__9504 (
            .O(N__44785),
            .I(N__44782));
    Odrv12 I__9503 (
            .O(N__44782),
            .I(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ));
    InMux I__9502 (
            .O(N__44779),
            .I(N__44776));
    LocalMux I__9501 (
            .O(N__44776),
            .I(\current_shift_inst.un38_control_input_0_s0_11 ));
    InMux I__9500 (
            .O(N__44773),
            .I(\current_shift_inst.un38_control_input_cry_10_s0 ));
    CascadeMux I__9499 (
            .O(N__44770),
            .I(N__44767));
    InMux I__9498 (
            .O(N__44767),
            .I(N__44762));
    InMux I__9497 (
            .O(N__44766),
            .I(N__44756));
    InMux I__9496 (
            .O(N__44765),
            .I(N__44756));
    LocalMux I__9495 (
            .O(N__44762),
            .I(N__44753));
    InMux I__9494 (
            .O(N__44761),
            .I(N__44750));
    LocalMux I__9493 (
            .O(N__44756),
            .I(N__44747));
    Span4Mux_v I__9492 (
            .O(N__44753),
            .I(N__44744));
    LocalMux I__9491 (
            .O(N__44750),
            .I(N__44741));
    Span4Mux_h I__9490 (
            .O(N__44747),
            .I(N__44738));
    Odrv4 I__9489 (
            .O(N__44744),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv12 I__9488 (
            .O(N__44741),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    Odrv4 I__9487 (
            .O(N__44738),
            .I(\current_shift_inst.elapsed_time_ns_s1_26 ));
    InMux I__9486 (
            .O(N__44731),
            .I(N__44727));
    CascadeMux I__9485 (
            .O(N__44730),
            .I(N__44724));
    LocalMux I__9484 (
            .O(N__44727),
            .I(N__44720));
    InMux I__9483 (
            .O(N__44724),
            .I(N__44717));
    InMux I__9482 (
            .O(N__44723),
            .I(N__44714));
    Odrv12 I__9481 (
            .O(N__44720),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9480 (
            .O(N__44717),
            .I(\current_shift_inst.un4_control_input1_26 ));
    LocalMux I__9479 (
            .O(N__44714),
            .I(\current_shift_inst.un4_control_input1_26 ));
    InMux I__9478 (
            .O(N__44707),
            .I(N__44700));
    InMux I__9477 (
            .O(N__44706),
            .I(N__44700));
    CascadeMux I__9476 (
            .O(N__44705),
            .I(N__44697));
    LocalMux I__9475 (
            .O(N__44700),
            .I(N__44694));
    InMux I__9474 (
            .O(N__44697),
            .I(N__44691));
    Span4Mux_h I__9473 (
            .O(N__44694),
            .I(N__44688));
    LocalMux I__9472 (
            .O(N__44691),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    Odrv4 I__9471 (
            .O(N__44688),
            .I(\current_shift_inst.un4_control_input1_31_THRU_CO ));
    InMux I__9470 (
            .O(N__44683),
            .I(N__44677));
    InMux I__9469 (
            .O(N__44682),
            .I(N__44677));
    LocalMux I__9468 (
            .O(N__44677),
            .I(N__44673));
    InMux I__9467 (
            .O(N__44676),
            .I(N__44670));
    Span4Mux_h I__9466 (
            .O(N__44673),
            .I(N__44664));
    LocalMux I__9465 (
            .O(N__44670),
            .I(N__44664));
    InMux I__9464 (
            .O(N__44669),
            .I(N__44661));
    Odrv4 I__9463 (
            .O(N__44664),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    LocalMux I__9462 (
            .O(N__44661),
            .I(\current_shift_inst.elapsed_time_ns_s1_21 ));
    InMux I__9461 (
            .O(N__44656),
            .I(N__44649));
    InMux I__9460 (
            .O(N__44655),
            .I(N__44649));
    InMux I__9459 (
            .O(N__44654),
            .I(N__44646));
    LocalMux I__9458 (
            .O(N__44649),
            .I(N__44643));
    LocalMux I__9457 (
            .O(N__44646),
            .I(N__44640));
    Odrv4 I__9456 (
            .O(N__44643),
            .I(\current_shift_inst.un4_control_input1_21 ));
    Odrv4 I__9455 (
            .O(N__44640),
            .I(\current_shift_inst.un4_control_input1_21 ));
    InMux I__9454 (
            .O(N__44635),
            .I(N__44632));
    LocalMux I__9453 (
            .O(N__44632),
            .I(N__44629));
    Odrv12 I__9452 (
            .O(N__44629),
            .I(\current_shift_inst.un38_control_input_cry_0_s0_sf ));
    CascadeMux I__9451 (
            .O(N__44626),
            .I(N__44623));
    InMux I__9450 (
            .O(N__44623),
            .I(N__44620));
    LocalMux I__9449 (
            .O(N__44620),
            .I(N__44617));
    Span4Mux_h I__9448 (
            .O(N__44617),
            .I(N__44614));
    Span4Mux_v I__9447 (
            .O(N__44614),
            .I(N__44611));
    Odrv4 I__9446 (
            .O(N__44611),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ));
    CascadeMux I__9445 (
            .O(N__44608),
            .I(N__44605));
    InMux I__9444 (
            .O(N__44605),
            .I(N__44602));
    LocalMux I__9443 (
            .O(N__44602),
            .I(N__44599));
    Span4Mux_h I__9442 (
            .O(N__44599),
            .I(N__44596));
    Odrv4 I__9441 (
            .O(N__44596),
            .I(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ));
    InMux I__9440 (
            .O(N__44593),
            .I(N__44590));
    LocalMux I__9439 (
            .O(N__44590),
            .I(N__44587));
    Odrv12 I__9438 (
            .O(N__44587),
            .I(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ));
    InMux I__9437 (
            .O(N__44584),
            .I(N__44581));
    LocalMux I__9436 (
            .O(N__44581),
            .I(\current_shift_inst.un38_control_input_0_s0_3 ));
    InMux I__9435 (
            .O(N__44578),
            .I(\current_shift_inst.un38_control_input_cry_2_s0 ));
    InMux I__9434 (
            .O(N__44575),
            .I(N__44569));
    InMux I__9433 (
            .O(N__44574),
            .I(N__44569));
    LocalMux I__9432 (
            .O(N__44569),
            .I(N__44565));
    InMux I__9431 (
            .O(N__44568),
            .I(N__44562));
    Span4Mux_v I__9430 (
            .O(N__44565),
            .I(N__44556));
    LocalMux I__9429 (
            .O(N__44562),
            .I(N__44556));
    InMux I__9428 (
            .O(N__44561),
            .I(N__44553));
    Odrv4 I__9427 (
            .O(N__44556),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    LocalMux I__9426 (
            .O(N__44553),
            .I(\current_shift_inst.elapsed_time_ns_s1_22 ));
    CascadeMux I__9425 (
            .O(N__44548),
            .I(N__44544));
    InMux I__9424 (
            .O(N__44547),
            .I(N__44540));
    InMux I__9423 (
            .O(N__44544),
            .I(N__44535));
    InMux I__9422 (
            .O(N__44543),
            .I(N__44535));
    LocalMux I__9421 (
            .O(N__44540),
            .I(N__44532));
    LocalMux I__9420 (
            .O(N__44535),
            .I(\current_shift_inst.un4_control_input1_22 ));
    Odrv4 I__9419 (
            .O(N__44532),
            .I(\current_shift_inst.un4_control_input1_22 ));
    CascadeMux I__9418 (
            .O(N__44527),
            .I(N__44523));
    CascadeMux I__9417 (
            .O(N__44526),
            .I(N__44520));
    InMux I__9416 (
            .O(N__44523),
            .I(N__44517));
    InMux I__9415 (
            .O(N__44520),
            .I(N__44514));
    LocalMux I__9414 (
            .O(N__44517),
            .I(N__44510));
    LocalMux I__9413 (
            .O(N__44514),
            .I(N__44507));
    InMux I__9412 (
            .O(N__44513),
            .I(N__44504));
    Span4Mux_v I__9411 (
            .O(N__44510),
            .I(N__44498));
    Span4Mux_v I__9410 (
            .O(N__44507),
            .I(N__44498));
    LocalMux I__9409 (
            .O(N__44504),
            .I(N__44495));
    InMux I__9408 (
            .O(N__44503),
            .I(N__44492));
    Odrv4 I__9407 (
            .O(N__44498),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    Odrv4 I__9406 (
            .O(N__44495),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    LocalMux I__9405 (
            .O(N__44492),
            .I(\current_shift_inst.elapsed_time_ns_s1_5 ));
    InMux I__9404 (
            .O(N__44485),
            .I(N__44481));
    InMux I__9403 (
            .O(N__44484),
            .I(N__44478));
    LocalMux I__9402 (
            .O(N__44481),
            .I(N__44474));
    LocalMux I__9401 (
            .O(N__44478),
            .I(N__44471));
    InMux I__9400 (
            .O(N__44477),
            .I(N__44468));
    Odrv12 I__9399 (
            .O(N__44474),
            .I(\current_shift_inst.un4_control_input1_5 ));
    Odrv4 I__9398 (
            .O(N__44471),
            .I(\current_shift_inst.un4_control_input1_5 ));
    LocalMux I__9397 (
            .O(N__44468),
            .I(\current_shift_inst.un4_control_input1_5 ));
    InMux I__9396 (
            .O(N__44461),
            .I(N__44457));
    InMux I__9395 (
            .O(N__44460),
            .I(N__44454));
    LocalMux I__9394 (
            .O(N__44457),
            .I(N__44450));
    LocalMux I__9393 (
            .O(N__44454),
            .I(N__44447));
    InMux I__9392 (
            .O(N__44453),
            .I(N__44444));
    Span4Mux_h I__9391 (
            .O(N__44450),
            .I(N__44440));
    Span4Mux_v I__9390 (
            .O(N__44447),
            .I(N__44435));
    LocalMux I__9389 (
            .O(N__44444),
            .I(N__44435));
    InMux I__9388 (
            .O(N__44443),
            .I(N__44432));
    Odrv4 I__9387 (
            .O(N__44440),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    Odrv4 I__9386 (
            .O(N__44435),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    LocalMux I__9385 (
            .O(N__44432),
            .I(\current_shift_inst.elapsed_time_ns_s1_16 ));
    CascadeMux I__9384 (
            .O(N__44425),
            .I(N__44422));
    InMux I__9383 (
            .O(N__44422),
            .I(N__44418));
    InMux I__9382 (
            .O(N__44421),
            .I(N__44415));
    LocalMux I__9381 (
            .O(N__44418),
            .I(N__44411));
    LocalMux I__9380 (
            .O(N__44415),
            .I(N__44408));
    InMux I__9379 (
            .O(N__44414),
            .I(N__44405));
    Span4Mux_h I__9378 (
            .O(N__44411),
            .I(N__44398));
    Span4Mux_v I__9377 (
            .O(N__44408),
            .I(N__44398));
    LocalMux I__9376 (
            .O(N__44405),
            .I(N__44398));
    Odrv4 I__9375 (
            .O(N__44398),
            .I(\current_shift_inst.un4_control_input1_16 ));
    CascadeMux I__9374 (
            .O(N__44395),
            .I(N__44392));
    InMux I__9373 (
            .O(N__44392),
            .I(N__44387));
    InMux I__9372 (
            .O(N__44391),
            .I(N__44384));
    CascadeMux I__9371 (
            .O(N__44390),
            .I(N__44381));
    LocalMux I__9370 (
            .O(N__44387),
            .I(N__44378));
    LocalMux I__9369 (
            .O(N__44384),
            .I(N__44375));
    InMux I__9368 (
            .O(N__44381),
            .I(N__44372));
    Span4Mux_v I__9367 (
            .O(N__44378),
            .I(N__44366));
    Span4Mux_v I__9366 (
            .O(N__44375),
            .I(N__44366));
    LocalMux I__9365 (
            .O(N__44372),
            .I(N__44363));
    InMux I__9364 (
            .O(N__44371),
            .I(N__44360));
    Odrv4 I__9363 (
            .O(N__44366),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    Odrv12 I__9362 (
            .O(N__44363),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    LocalMux I__9361 (
            .O(N__44360),
            .I(\current_shift_inst.elapsed_time_ns_s1_28 ));
    InMux I__9360 (
            .O(N__44353),
            .I(N__44350));
    LocalMux I__9359 (
            .O(N__44350),
            .I(N__44345));
    InMux I__9358 (
            .O(N__44349),
            .I(N__44342));
    InMux I__9357 (
            .O(N__44348),
            .I(N__44339));
    Span4Mux_v I__9356 (
            .O(N__44345),
            .I(N__44334));
    LocalMux I__9355 (
            .O(N__44342),
            .I(N__44334));
    LocalMux I__9354 (
            .O(N__44339),
            .I(\current_shift_inst.un4_control_input1_28 ));
    Odrv4 I__9353 (
            .O(N__44334),
            .I(\current_shift_inst.un4_control_input1_28 ));
    CascadeMux I__9352 (
            .O(N__44329),
            .I(N__44325));
    InMux I__9351 (
            .O(N__44328),
            .I(N__44321));
    InMux I__9350 (
            .O(N__44325),
            .I(N__44315));
    InMux I__9349 (
            .O(N__44324),
            .I(N__44315));
    LocalMux I__9348 (
            .O(N__44321),
            .I(N__44312));
    InMux I__9347 (
            .O(N__44320),
            .I(N__44309));
    LocalMux I__9346 (
            .O(N__44315),
            .I(N__44306));
    Span4Mux_v I__9345 (
            .O(N__44312),
            .I(N__44299));
    LocalMux I__9344 (
            .O(N__44309),
            .I(N__44299));
    Span4Mux_v I__9343 (
            .O(N__44306),
            .I(N__44299));
    Odrv4 I__9342 (
            .O(N__44299),
            .I(\current_shift_inst.elapsed_time_ns_s1_27 ));
    InMux I__9341 (
            .O(N__44296),
            .I(N__44293));
    LocalMux I__9340 (
            .O(N__44293),
            .I(N__44288));
    InMux I__9339 (
            .O(N__44292),
            .I(N__44285));
    InMux I__9338 (
            .O(N__44291),
            .I(N__44282));
    Span4Mux_v I__9337 (
            .O(N__44288),
            .I(N__44277));
    LocalMux I__9336 (
            .O(N__44285),
            .I(N__44277));
    LocalMux I__9335 (
            .O(N__44282),
            .I(\current_shift_inst.un4_control_input1_27 ));
    Odrv4 I__9334 (
            .O(N__44277),
            .I(\current_shift_inst.un4_control_input1_27 ));
    InMux I__9333 (
            .O(N__44272),
            .I(N__44266));
    InMux I__9332 (
            .O(N__44271),
            .I(N__44266));
    LocalMux I__9331 (
            .O(N__44266),
            .I(N__44261));
    InMux I__9330 (
            .O(N__44265),
            .I(N__44258));
    InMux I__9329 (
            .O(N__44264),
            .I(N__44255));
    Odrv12 I__9328 (
            .O(N__44261),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__9327 (
            .O(N__44258),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    LocalMux I__9326 (
            .O(N__44255),
            .I(\current_shift_inst.elapsed_time_ns_s1_10 ));
    CascadeMux I__9325 (
            .O(N__44248),
            .I(N__44244));
    InMux I__9324 (
            .O(N__44247),
            .I(N__44238));
    InMux I__9323 (
            .O(N__44244),
            .I(N__44238));
    InMux I__9322 (
            .O(N__44243),
            .I(N__44235));
    LocalMux I__9321 (
            .O(N__44238),
            .I(\current_shift_inst.un4_control_input1_10 ));
    LocalMux I__9320 (
            .O(N__44235),
            .I(\current_shift_inst.un4_control_input1_10 ));
    InMux I__9319 (
            .O(N__44230),
            .I(N__44227));
    LocalMux I__9318 (
            .O(N__44227),
            .I(N__44223));
    InMux I__9317 (
            .O(N__44226),
            .I(N__44220));
    Span4Mux_h I__9316 (
            .O(N__44223),
            .I(N__44217));
    LocalMux I__9315 (
            .O(N__44220),
            .I(N__44214));
    Span4Mux_v I__9314 (
            .O(N__44217),
            .I(N__44210));
    Span4Mux_v I__9313 (
            .O(N__44214),
            .I(N__44207));
    InMux I__9312 (
            .O(N__44213),
            .I(N__44204));
    Odrv4 I__9311 (
            .O(N__44210),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    Odrv4 I__9310 (
            .O(N__44207),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    LocalMux I__9309 (
            .O(N__44204),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ));
    CEMux I__9308 (
            .O(N__44197),
            .I(N__44176));
    CEMux I__9307 (
            .O(N__44196),
            .I(N__44176));
    CEMux I__9306 (
            .O(N__44195),
            .I(N__44176));
    CEMux I__9305 (
            .O(N__44194),
            .I(N__44176));
    CEMux I__9304 (
            .O(N__44193),
            .I(N__44176));
    CEMux I__9303 (
            .O(N__44192),
            .I(N__44176));
    CEMux I__9302 (
            .O(N__44191),
            .I(N__44176));
    GlobalMux I__9301 (
            .O(N__44176),
            .I(N__44173));
    gio2CtrlBuf I__9300 (
            .O(N__44173),
            .I(\current_shift_inst.timer_s1.N_163_i_g ));
    CascadeMux I__9299 (
            .O(N__44170),
            .I(N__44167));
    InMux I__9298 (
            .O(N__44167),
            .I(N__44161));
    InMux I__9297 (
            .O(N__44166),
            .I(N__44161));
    LocalMux I__9296 (
            .O(N__44161),
            .I(N__44157));
    InMux I__9295 (
            .O(N__44160),
            .I(N__44154));
    Odrv4 I__9294 (
            .O(N__44157),
            .I(\current_shift_inst.un4_control_input1_3 ));
    LocalMux I__9293 (
            .O(N__44154),
            .I(\current_shift_inst.un4_control_input1_3 ));
    InMux I__9292 (
            .O(N__44149),
            .I(N__44144));
    InMux I__9291 (
            .O(N__44148),
            .I(N__44139));
    InMux I__9290 (
            .O(N__44147),
            .I(N__44139));
    LocalMux I__9289 (
            .O(N__44144),
            .I(N__44136));
    LocalMux I__9288 (
            .O(N__44139),
            .I(N__44132));
    Span4Mux_v I__9287 (
            .O(N__44136),
            .I(N__44129));
    InMux I__9286 (
            .O(N__44135),
            .I(N__44126));
    Odrv4 I__9285 (
            .O(N__44132),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    Odrv4 I__9284 (
            .O(N__44129),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    LocalMux I__9283 (
            .O(N__44126),
            .I(\current_shift_inst.elapsed_time_ns_s1_3 ));
    InMux I__9282 (
            .O(N__44119),
            .I(N__44115));
    CascadeMux I__9281 (
            .O(N__44118),
            .I(N__44111));
    LocalMux I__9280 (
            .O(N__44115),
            .I(N__44108));
    InMux I__9279 (
            .O(N__44114),
            .I(N__44105));
    InMux I__9278 (
            .O(N__44111),
            .I(N__44102));
    Odrv4 I__9277 (
            .O(N__44108),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__9276 (
            .O(N__44105),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    LocalMux I__9275 (
            .O(N__44102),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1 ));
    InMux I__9274 (
            .O(N__44095),
            .I(N__44092));
    LocalMux I__9273 (
            .O(N__44092),
            .I(\current_shift_inst.un4_control_input1_1 ));
    CascadeMux I__9272 (
            .O(N__44089),
            .I(\current_shift_inst.un4_control_input1_1_cascade_ ));
    InMux I__9271 (
            .O(N__44086),
            .I(N__44082));
    InMux I__9270 (
            .O(N__44085),
            .I(N__44079));
    LocalMux I__9269 (
            .O(N__44082),
            .I(N__44072));
    LocalMux I__9268 (
            .O(N__44079),
            .I(N__44072));
    InMux I__9267 (
            .O(N__44078),
            .I(N__44067));
    InMux I__9266 (
            .O(N__44077),
            .I(N__44067));
    Odrv4 I__9265 (
            .O(N__44072),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    LocalMux I__9264 (
            .O(N__44067),
            .I(\current_shift_inst.elapsed_time_ns_s1_1 ));
    CascadeMux I__9263 (
            .O(N__44062),
            .I(N__44058));
    CascadeMux I__9262 (
            .O(N__44061),
            .I(N__44055));
    InMux I__9261 (
            .O(N__44058),
            .I(N__44052));
    InMux I__9260 (
            .O(N__44055),
            .I(N__44049));
    LocalMux I__9259 (
            .O(N__44052),
            .I(N__44046));
    LocalMux I__9258 (
            .O(N__44049),
            .I(N__44039));
    Span4Mux_v I__9257 (
            .O(N__44046),
            .I(N__44039));
    InMux I__9256 (
            .O(N__44045),
            .I(N__44036));
    InMux I__9255 (
            .O(N__44044),
            .I(N__44033));
    Odrv4 I__9254 (
            .O(N__44039),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__9253 (
            .O(N__44036),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    LocalMux I__9252 (
            .O(N__44033),
            .I(\current_shift_inst.elapsed_time_ns_s1_13 ));
    InMux I__9251 (
            .O(N__44026),
            .I(N__44023));
    LocalMux I__9250 (
            .O(N__44023),
            .I(N__44018));
    InMux I__9249 (
            .O(N__44022),
            .I(N__44015));
    InMux I__9248 (
            .O(N__44021),
            .I(N__44012));
    Odrv4 I__9247 (
            .O(N__44018),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9246 (
            .O(N__44015),
            .I(\current_shift_inst.un4_control_input1_13 ));
    LocalMux I__9245 (
            .O(N__44012),
            .I(\current_shift_inst.un4_control_input1_13 ));
    InMux I__9244 (
            .O(N__44005),
            .I(N__44002));
    LocalMux I__9243 (
            .O(N__44002),
            .I(\current_shift_inst.un4_control_input_1_axb_18 ));
    InMux I__9242 (
            .O(N__43999),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ));
    InMux I__9241 (
            .O(N__43996),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ));
    InMux I__9240 (
            .O(N__43993),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ));
    InMux I__9239 (
            .O(N__43990),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ));
    InMux I__9238 (
            .O(N__43987),
            .I(bfn_17_13_0_));
    InMux I__9237 (
            .O(N__43984),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__9236 (
            .O(N__43981),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__9235 (
            .O(N__43978),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__9234 (
            .O(N__43975),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ));
    CEMux I__9233 (
            .O(N__43972),
            .I(N__43967));
    CEMux I__9232 (
            .O(N__43971),
            .I(N__43964));
    CEMux I__9231 (
            .O(N__43970),
            .I(N__43960));
    LocalMux I__9230 (
            .O(N__43967),
            .I(N__43956));
    LocalMux I__9229 (
            .O(N__43964),
            .I(N__43953));
    CEMux I__9228 (
            .O(N__43963),
            .I(N__43950));
    LocalMux I__9227 (
            .O(N__43960),
            .I(N__43947));
    CEMux I__9226 (
            .O(N__43959),
            .I(N__43944));
    Span4Mux_v I__9225 (
            .O(N__43956),
            .I(N__43941));
    Span4Mux_h I__9224 (
            .O(N__43953),
            .I(N__43938));
    LocalMux I__9223 (
            .O(N__43950),
            .I(N__43935));
    Span4Mux_h I__9222 (
            .O(N__43947),
            .I(N__43930));
    LocalMux I__9221 (
            .O(N__43944),
            .I(N__43930));
    Span4Mux_h I__9220 (
            .O(N__43941),
            .I(N__43927));
    Span4Mux_h I__9219 (
            .O(N__43938),
            .I(N__43924));
    Span4Mux_h I__9218 (
            .O(N__43935),
            .I(N__43921));
    Span4Mux_h I__9217 (
            .O(N__43930),
            .I(N__43918));
    Odrv4 I__9216 (
            .O(N__43927),
            .I(\delay_measurement_inst.delay_hc_timer.N_165_i ));
    Odrv4 I__9215 (
            .O(N__43924),
            .I(\delay_measurement_inst.delay_hc_timer.N_165_i ));
    Odrv4 I__9214 (
            .O(N__43921),
            .I(\delay_measurement_inst.delay_hc_timer.N_165_i ));
    Odrv4 I__9213 (
            .O(N__43918),
            .I(\delay_measurement_inst.delay_hc_timer.N_165_i ));
    InMux I__9212 (
            .O(N__43909),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__9211 (
            .O(N__43906),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ));
    InMux I__9210 (
            .O(N__43903),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ));
    InMux I__9209 (
            .O(N__43900),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ));
    InMux I__9208 (
            .O(N__43897),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ));
    InMux I__9207 (
            .O(N__43894),
            .I(bfn_17_12_0_));
    InMux I__9206 (
            .O(N__43891),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ));
    InMux I__9205 (
            .O(N__43888),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ));
    InMux I__9204 (
            .O(N__43885),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__9203 (
            .O(N__43882),
            .I(N__43879));
    LocalMux I__9202 (
            .O(N__43879),
            .I(N__43875));
    InMux I__9201 (
            .O(N__43878),
            .I(N__43872));
    Odrv4 I__9200 (
            .O(N__43875),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    LocalMux I__9199 (
            .O(N__43872),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ));
    InMux I__9198 (
            .O(N__43867),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ));
    InMux I__9197 (
            .O(N__43864),
            .I(N__43860));
    InMux I__9196 (
            .O(N__43863),
            .I(N__43857));
    LocalMux I__9195 (
            .O(N__43860),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    LocalMux I__9194 (
            .O(N__43857),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ));
    InMux I__9193 (
            .O(N__43852),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ));
    InMux I__9192 (
            .O(N__43849),
            .I(N__43845));
    InMux I__9191 (
            .O(N__43848),
            .I(N__43842));
    LocalMux I__9190 (
            .O(N__43845),
            .I(N__43839));
    LocalMux I__9189 (
            .O(N__43842),
            .I(N__43836));
    Span4Mux_v I__9188 (
            .O(N__43839),
            .I(N__43833));
    Odrv12 I__9187 (
            .O(N__43836),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    Odrv4 I__9186 (
            .O(N__43833),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ));
    InMux I__9185 (
            .O(N__43828),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__9184 (
            .O(N__43825),
            .I(N__43822));
    InMux I__9183 (
            .O(N__43822),
            .I(N__43818));
    InMux I__9182 (
            .O(N__43821),
            .I(N__43815));
    LocalMux I__9181 (
            .O(N__43818),
            .I(N__43812));
    LocalMux I__9180 (
            .O(N__43815),
            .I(N__43809));
    Span4Mux_v I__9179 (
            .O(N__43812),
            .I(N__43806));
    Odrv4 I__9178 (
            .O(N__43809),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    Odrv4 I__9177 (
            .O(N__43806),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ));
    InMux I__9176 (
            .O(N__43801),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ));
    InMux I__9175 (
            .O(N__43798),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ));
    InMux I__9174 (
            .O(N__43795),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ));
    InMux I__9173 (
            .O(N__43792),
            .I(bfn_17_11_0_));
    InMux I__9172 (
            .O(N__43789),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ));
    InMux I__9171 (
            .O(N__43786),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ));
    InMux I__9170 (
            .O(N__43783),
            .I(N__43780));
    LocalMux I__9169 (
            .O(N__43780),
            .I(elapsed_time_ns_1_RNII43T9_0_6));
    CascadeMux I__9168 (
            .O(N__43777),
            .I(elapsed_time_ns_1_RNII43T9_0_6_cascade_));
    InMux I__9167 (
            .O(N__43774),
            .I(N__43771));
    LocalMux I__9166 (
            .O(N__43771),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ));
    InMux I__9165 (
            .O(N__43768),
            .I(N__43765));
    LocalMux I__9164 (
            .O(N__43765),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11));
    CascadeMux I__9163 (
            .O(N__43762),
            .I(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_));
    InMux I__9162 (
            .O(N__43759),
            .I(N__43756));
    LocalMux I__9161 (
            .O(N__43756),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ));
    InMux I__9160 (
            .O(N__43753),
            .I(N__43747));
    InMux I__9159 (
            .O(N__43752),
            .I(N__43747));
    LocalMux I__9158 (
            .O(N__43747),
            .I(elapsed_time_ns_1_RNI24CN9_0_15));
    InMux I__9157 (
            .O(N__43744),
            .I(N__43741));
    LocalMux I__9156 (
            .O(N__43741),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ));
    InMux I__9155 (
            .O(N__43738),
            .I(N__43732));
    InMux I__9154 (
            .O(N__43737),
            .I(N__43732));
    LocalMux I__9153 (
            .O(N__43732),
            .I(elapsed_time_ns_1_RNIV0CN9_0_12));
    InMux I__9152 (
            .O(N__43729),
            .I(N__43726));
    LocalMux I__9151 (
            .O(N__43726),
            .I(N__43722));
    InMux I__9150 (
            .O(N__43725),
            .I(N__43719));
    Span4Mux_v I__9149 (
            .O(N__43722),
            .I(N__43714));
    LocalMux I__9148 (
            .O(N__43719),
            .I(N__43714));
    Odrv4 I__9147 (
            .O(N__43714),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ));
    InMux I__9146 (
            .O(N__43711),
            .I(N__43707));
    CascadeMux I__9145 (
            .O(N__43710),
            .I(N__43704));
    LocalMux I__9144 (
            .O(N__43707),
            .I(N__43701));
    InMux I__9143 (
            .O(N__43704),
            .I(N__43698));
    Span4Mux_v I__9142 (
            .O(N__43701),
            .I(N__43693));
    LocalMux I__9141 (
            .O(N__43698),
            .I(N__43693));
    Odrv4 I__9140 (
            .O(N__43693),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ));
    InMux I__9139 (
            .O(N__43690),
            .I(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__9138 (
            .O(N__43687),
            .I(N__43684));
    LocalMux I__9137 (
            .O(N__43684),
            .I(elapsed_time_ns_1_RNITUBN9_0_10));
    CascadeMux I__9136 (
            .O(N__43681),
            .I(elapsed_time_ns_1_RNITUBN9_0_10_cascade_));
    InMux I__9135 (
            .O(N__43678),
            .I(N__43675));
    LocalMux I__9134 (
            .O(N__43675),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ));
    InMux I__9133 (
            .O(N__43672),
            .I(N__43669));
    LocalMux I__9132 (
            .O(N__43669),
            .I(elapsed_time_ns_1_RNIK63T9_0_8));
    CascadeMux I__9131 (
            .O(N__43666),
            .I(elapsed_time_ns_1_RNIK63T9_0_8_cascade_));
    InMux I__9130 (
            .O(N__43663),
            .I(N__43660));
    LocalMux I__9129 (
            .O(N__43660),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ));
    InMux I__9128 (
            .O(N__43657),
            .I(N__43651));
    InMux I__9127 (
            .O(N__43656),
            .I(N__43651));
    LocalMux I__9126 (
            .O(N__43651),
            .I(elapsed_time_ns_1_RNI35CN9_0_16));
    InMux I__9125 (
            .O(N__43648),
            .I(N__43645));
    LocalMux I__9124 (
            .O(N__43645),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ));
    InMux I__9123 (
            .O(N__43642),
            .I(N__43639));
    LocalMux I__9122 (
            .O(N__43639),
            .I(elapsed_time_ns_1_RNIL73T9_0_9));
    CascadeMux I__9121 (
            .O(N__43636),
            .I(elapsed_time_ns_1_RNIL73T9_0_9_cascade_));
    InMux I__9120 (
            .O(N__43633),
            .I(N__43630));
    LocalMux I__9119 (
            .O(N__43630),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ));
    InMux I__9118 (
            .O(N__43627),
            .I(N__43624));
    LocalMux I__9117 (
            .O(N__43624),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ));
    InMux I__9116 (
            .O(N__43621),
            .I(N__43616));
    InMux I__9115 (
            .O(N__43620),
            .I(N__43613));
    InMux I__9114 (
            .O(N__43619),
            .I(N__43610));
    LocalMux I__9113 (
            .O(N__43616),
            .I(N__43605));
    LocalMux I__9112 (
            .O(N__43613),
            .I(N__43605));
    LocalMux I__9111 (
            .O(N__43610),
            .I(N__43602));
    Odrv12 I__9110 (
            .O(N__43605),
            .I(\current_shift_inst.un4_control_input1_25 ));
    Odrv4 I__9109 (
            .O(N__43602),
            .I(\current_shift_inst.un4_control_input1_25 ));
    InMux I__9108 (
            .O(N__43597),
            .I(N__43594));
    LocalMux I__9107 (
            .O(N__43594),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7));
    CascadeMux I__9106 (
            .O(N__43591),
            .I(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_));
    InMux I__9105 (
            .O(N__43588),
            .I(N__43585));
    LocalMux I__9104 (
            .O(N__43585),
            .I(N__43582));
    Odrv4 I__9103 (
            .O(N__43582),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ));
    InMux I__9102 (
            .O(N__43579),
            .I(N__43575));
    InMux I__9101 (
            .O(N__43578),
            .I(N__43572));
    LocalMux I__9100 (
            .O(N__43575),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    LocalMux I__9099 (
            .O(N__43572),
            .I(elapsed_time_ns_1_RNI25DN9_0_24));
    InMux I__9098 (
            .O(N__43567),
            .I(N__43564));
    LocalMux I__9097 (
            .O(N__43564),
            .I(N__43561));
    Span4Mux_v I__9096 (
            .O(N__43561),
            .I(N__43558));
    Odrv4 I__9095 (
            .O(N__43558),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ));
    InMux I__9094 (
            .O(N__43555),
            .I(N__43552));
    LocalMux I__9093 (
            .O(N__43552),
            .I(N__43549));
    Span4Mux_v I__9092 (
            .O(N__43549),
            .I(N__43546));
    Odrv4 I__9091 (
            .O(N__43546),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ));
    InMux I__9090 (
            .O(N__43543),
            .I(N__43540));
    LocalMux I__9089 (
            .O(N__43540),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20));
    CascadeMux I__9088 (
            .O(N__43537),
            .I(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_));
    InMux I__9087 (
            .O(N__43534),
            .I(N__43531));
    LocalMux I__9086 (
            .O(N__43531),
            .I(N__43528));
    Odrv4 I__9085 (
            .O(N__43528),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ));
    InMux I__9084 (
            .O(N__43525),
            .I(N__43522));
    LocalMux I__9083 (
            .O(N__43522),
            .I(elapsed_time_ns_1_RNIH33T9_0_5));
    CascadeMux I__9082 (
            .O(N__43519),
            .I(elapsed_time_ns_1_RNIH33T9_0_5_cascade_));
    InMux I__9081 (
            .O(N__43516),
            .I(N__43513));
    LocalMux I__9080 (
            .O(N__43513),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ));
    InMux I__9079 (
            .O(N__43510),
            .I(N__43507));
    LocalMux I__9078 (
            .O(N__43507),
            .I(N__43504));
    Odrv4 I__9077 (
            .O(N__43504),
            .I(\current_shift_inst.control_input_axb_19 ));
    CascadeMux I__9076 (
            .O(N__43501),
            .I(N__43497));
    InMux I__9075 (
            .O(N__43500),
            .I(N__43494));
    InMux I__9074 (
            .O(N__43497),
            .I(N__43491));
    LocalMux I__9073 (
            .O(N__43494),
            .I(N__43484));
    LocalMux I__9072 (
            .O(N__43491),
            .I(N__43484));
    InMux I__9071 (
            .O(N__43490),
            .I(N__43481));
    InMux I__9070 (
            .O(N__43489),
            .I(N__43478));
    Span4Mux_v I__9069 (
            .O(N__43484),
            .I(N__43471));
    LocalMux I__9068 (
            .O(N__43481),
            .I(N__43471));
    LocalMux I__9067 (
            .O(N__43478),
            .I(N__43471));
    Odrv4 I__9066 (
            .O(N__43471),
            .I(\current_shift_inst.elapsed_time_ns_s1_30 ));
    InMux I__9065 (
            .O(N__43468),
            .I(N__43464));
    InMux I__9064 (
            .O(N__43467),
            .I(N__43461));
    LocalMux I__9063 (
            .O(N__43464),
            .I(N__43457));
    LocalMux I__9062 (
            .O(N__43461),
            .I(N__43454));
    InMux I__9061 (
            .O(N__43460),
            .I(N__43451));
    Span4Mux_v I__9060 (
            .O(N__43457),
            .I(N__43448));
    Span4Mux_v I__9059 (
            .O(N__43454),
            .I(N__43443));
    LocalMux I__9058 (
            .O(N__43451),
            .I(N__43443));
    Odrv4 I__9057 (
            .O(N__43448),
            .I(\current_shift_inst.un4_control_input1_30 ));
    Odrv4 I__9056 (
            .O(N__43443),
            .I(\current_shift_inst.un4_control_input1_30 ));
    InMux I__9055 (
            .O(N__43438),
            .I(N__43435));
    LocalMux I__9054 (
            .O(N__43435),
            .I(N__43432));
    Odrv12 I__9053 (
            .O(N__43432),
            .I(\current_shift_inst.un4_control_input_1_axb_26 ));
    InMux I__9052 (
            .O(N__43429),
            .I(N__43426));
    LocalMux I__9051 (
            .O(N__43426),
            .I(N__43423));
    Odrv4 I__9050 (
            .O(N__43423),
            .I(\current_shift_inst.control_input_axb_20 ));
    CascadeMux I__9049 (
            .O(N__43420),
            .I(N__43416));
    CascadeMux I__9048 (
            .O(N__43419),
            .I(N__43413));
    InMux I__9047 (
            .O(N__43416),
            .I(N__43410));
    InMux I__9046 (
            .O(N__43413),
            .I(N__43407));
    LocalMux I__9045 (
            .O(N__43410),
            .I(N__43403));
    LocalMux I__9044 (
            .O(N__43407),
            .I(N__43400));
    InMux I__9043 (
            .O(N__43406),
            .I(N__43397));
    Span4Mux_v I__9042 (
            .O(N__43403),
            .I(N__43389));
    Span4Mux_v I__9041 (
            .O(N__43400),
            .I(N__43389));
    LocalMux I__9040 (
            .O(N__43397),
            .I(N__43389));
    InMux I__9039 (
            .O(N__43396),
            .I(N__43386));
    Odrv4 I__9038 (
            .O(N__43389),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    LocalMux I__9037 (
            .O(N__43386),
            .I(\current_shift_inst.elapsed_time_ns_s1_29 ));
    InMux I__9036 (
            .O(N__43381),
            .I(N__43376));
    InMux I__9035 (
            .O(N__43380),
            .I(N__43373));
    InMux I__9034 (
            .O(N__43379),
            .I(N__43370));
    LocalMux I__9033 (
            .O(N__43376),
            .I(N__43365));
    LocalMux I__9032 (
            .O(N__43373),
            .I(N__43365));
    LocalMux I__9031 (
            .O(N__43370),
            .I(N__43362));
    Odrv12 I__9030 (
            .O(N__43365),
            .I(\current_shift_inst.un4_control_input1_29 ));
    Odrv4 I__9029 (
            .O(N__43362),
            .I(\current_shift_inst.un4_control_input1_29 ));
    InMux I__9028 (
            .O(N__43357),
            .I(N__43354));
    LocalMux I__9027 (
            .O(N__43354),
            .I(N__43351));
    Span4Mux_h I__9026 (
            .O(N__43351),
            .I(N__43348));
    Odrv4 I__9025 (
            .O(N__43348),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ));
    InMux I__9024 (
            .O(N__43345),
            .I(N__43342));
    LocalMux I__9023 (
            .O(N__43342),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ));
    CascadeMux I__9022 (
            .O(N__43339),
            .I(N__43336));
    InMux I__9021 (
            .O(N__43336),
            .I(N__43333));
    LocalMux I__9020 (
            .O(N__43333),
            .I(N__43330));
    Span4Mux_h I__9019 (
            .O(N__43330),
            .I(N__43327));
    Odrv4 I__9018 (
            .O(N__43327),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ));
    InMux I__9017 (
            .O(N__43324),
            .I(N__43321));
    LocalMux I__9016 (
            .O(N__43321),
            .I(N__43318));
    Span4Mux_h I__9015 (
            .O(N__43318),
            .I(N__43315));
    Odrv4 I__9014 (
            .O(N__43315),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ));
    InMux I__9013 (
            .O(N__43312),
            .I(N__43309));
    LocalMux I__9012 (
            .O(N__43309),
            .I(N__43306));
    Span4Mux_h I__9011 (
            .O(N__43306),
            .I(N__43303));
    Odrv4 I__9010 (
            .O(N__43303),
            .I(\current_shift_inst.control_input_axb_11 ));
    InMux I__9009 (
            .O(N__43300),
            .I(N__43297));
    LocalMux I__9008 (
            .O(N__43297),
            .I(N__43294));
    Odrv4 I__9007 (
            .O(N__43294),
            .I(\current_shift_inst.control_input_axb_8 ));
    InMux I__9006 (
            .O(N__43291),
            .I(N__43288));
    LocalMux I__9005 (
            .O(N__43288),
            .I(N__43285));
    Odrv4 I__9004 (
            .O(N__43285),
            .I(\current_shift_inst.control_input_axb_14 ));
    InMux I__9003 (
            .O(N__43282),
            .I(N__43279));
    LocalMux I__9002 (
            .O(N__43279),
            .I(N__43276));
    Odrv4 I__9001 (
            .O(N__43276),
            .I(\current_shift_inst.control_input_axb_15 ));
    InMux I__9000 (
            .O(N__43273),
            .I(N__43270));
    LocalMux I__8999 (
            .O(N__43270),
            .I(N__43267));
    Odrv4 I__8998 (
            .O(N__43267),
            .I(\current_shift_inst.control_input_axb_12 ));
    InMux I__8997 (
            .O(N__43264),
            .I(N__43261));
    LocalMux I__8996 (
            .O(N__43261),
            .I(N__43258));
    Span4Mux_h I__8995 (
            .O(N__43258),
            .I(N__43255));
    Odrv4 I__8994 (
            .O(N__43255),
            .I(\current_shift_inst.control_input_axb_24 ));
    InMux I__8993 (
            .O(N__43252),
            .I(N__43249));
    LocalMux I__8992 (
            .O(N__43249),
            .I(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ));
    InMux I__8991 (
            .O(N__43246),
            .I(N__43243));
    LocalMux I__8990 (
            .O(N__43243),
            .I(N__43240));
    Odrv4 I__8989 (
            .O(N__43240),
            .I(\current_shift_inst.un4_control_input_1_axb_29 ));
    InMux I__8988 (
            .O(N__43237),
            .I(N__43224));
    InMux I__8987 (
            .O(N__43236),
            .I(N__43224));
    InMux I__8986 (
            .O(N__43235),
            .I(N__43207));
    InMux I__8985 (
            .O(N__43234),
            .I(N__43207));
    InMux I__8984 (
            .O(N__43233),
            .I(N__43207));
    InMux I__8983 (
            .O(N__43232),
            .I(N__43207));
    InMux I__8982 (
            .O(N__43231),
            .I(N__43207));
    InMux I__8981 (
            .O(N__43230),
            .I(N__43202));
    InMux I__8980 (
            .O(N__43229),
            .I(N__43202));
    LocalMux I__8979 (
            .O(N__43224),
            .I(N__43199));
    InMux I__8978 (
            .O(N__43223),
            .I(N__43192));
    InMux I__8977 (
            .O(N__43222),
            .I(N__43192));
    InMux I__8976 (
            .O(N__43221),
            .I(N__43192));
    InMux I__8975 (
            .O(N__43220),
            .I(N__43185));
    InMux I__8974 (
            .O(N__43219),
            .I(N__43185));
    InMux I__8973 (
            .O(N__43218),
            .I(N__43185));
    LocalMux I__8972 (
            .O(N__43207),
            .I(N__43170));
    LocalMux I__8971 (
            .O(N__43202),
            .I(N__43170));
    Span4Mux_v I__8970 (
            .O(N__43199),
            .I(N__43163));
    LocalMux I__8969 (
            .O(N__43192),
            .I(N__43163));
    LocalMux I__8968 (
            .O(N__43185),
            .I(N__43163));
    InMux I__8967 (
            .O(N__43184),
            .I(N__43154));
    InMux I__8966 (
            .O(N__43183),
            .I(N__43154));
    InMux I__8965 (
            .O(N__43182),
            .I(N__43154));
    InMux I__8964 (
            .O(N__43181),
            .I(N__43154));
    InMux I__8963 (
            .O(N__43180),
            .I(N__43147));
    InMux I__8962 (
            .O(N__43179),
            .I(N__43147));
    InMux I__8961 (
            .O(N__43178),
            .I(N__43147));
    InMux I__8960 (
            .O(N__43177),
            .I(N__43144));
    InMux I__8959 (
            .O(N__43176),
            .I(N__43139));
    InMux I__8958 (
            .O(N__43175),
            .I(N__43139));
    Odrv12 I__8957 (
            .O(N__43170),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    Odrv4 I__8956 (
            .O(N__43163),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8955 (
            .O(N__43154),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8954 (
            .O(N__43147),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8953 (
            .O(N__43144),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    LocalMux I__8952 (
            .O(N__43139),
            .I(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ));
    CascadeMux I__8951 (
            .O(N__43126),
            .I(N__43123));
    InMux I__8950 (
            .O(N__43123),
            .I(N__43120));
    LocalMux I__8949 (
            .O(N__43120),
            .I(N__43117));
    Odrv4 I__8948 (
            .O(N__43117),
            .I(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ));
    InMux I__8947 (
            .O(N__43114),
            .I(N__43111));
    LocalMux I__8946 (
            .O(N__43111),
            .I(N__43108));
    Span4Mux_h I__8945 (
            .O(N__43108),
            .I(N__43105));
    Odrv4 I__8944 (
            .O(N__43105),
            .I(\current_shift_inst.control_input_axb_9 ));
    InMux I__8943 (
            .O(N__43102),
            .I(N__43099));
    LocalMux I__8942 (
            .O(N__43099),
            .I(N__43096));
    Odrv4 I__8941 (
            .O(N__43096),
            .I(\current_shift_inst.control_input_axb_0 ));
    CascadeMux I__8940 (
            .O(N__43093),
            .I(\current_shift_inst.control_input_axb_0_cascade_ ));
    CascadeMux I__8939 (
            .O(N__43090),
            .I(N__43086));
    InMux I__8938 (
            .O(N__43089),
            .I(N__43082));
    InMux I__8937 (
            .O(N__43086),
            .I(N__43079));
    InMux I__8936 (
            .O(N__43085),
            .I(N__43076));
    LocalMux I__8935 (
            .O(N__43082),
            .I(N__43071));
    LocalMux I__8934 (
            .O(N__43079),
            .I(N__43071));
    LocalMux I__8933 (
            .O(N__43076),
            .I(\current_shift_inst.N_1379_i ));
    Odrv4 I__8932 (
            .O(N__43071),
            .I(\current_shift_inst.N_1379_i ));
    InMux I__8931 (
            .O(N__43066),
            .I(N__43063));
    LocalMux I__8930 (
            .O(N__43063),
            .I(N__43060));
    Span4Mux_h I__8929 (
            .O(N__43060),
            .I(N__43057));
    Odrv4 I__8928 (
            .O(N__43057),
            .I(\current_shift_inst.control_input_axb_10 ));
    CascadeMux I__8927 (
            .O(N__43054),
            .I(N__43051));
    InMux I__8926 (
            .O(N__43051),
            .I(N__43048));
    LocalMux I__8925 (
            .O(N__43048),
            .I(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ));
    InMux I__8924 (
            .O(N__43045),
            .I(N__43042));
    LocalMux I__8923 (
            .O(N__43042),
            .I(N__43039));
    Odrv4 I__8922 (
            .O(N__43039),
            .I(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ));
    CascadeMux I__8921 (
            .O(N__43036),
            .I(N__43033));
    InMux I__8920 (
            .O(N__43033),
            .I(N__43030));
    LocalMux I__8919 (
            .O(N__43030),
            .I(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ));
    CascadeMux I__8918 (
            .O(N__43027),
            .I(N__43024));
    InMux I__8917 (
            .O(N__43024),
            .I(N__43021));
    LocalMux I__8916 (
            .O(N__43021),
            .I(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ));
    CascadeMux I__8915 (
            .O(N__43018),
            .I(N__43015));
    InMux I__8914 (
            .O(N__43015),
            .I(N__43012));
    LocalMux I__8913 (
            .O(N__43012),
            .I(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ));
    InMux I__8912 (
            .O(N__43009),
            .I(N__43006));
    LocalMux I__8911 (
            .O(N__43006),
            .I(\current_shift_inst.un4_control_input_1_axb_25 ));
    CascadeMux I__8910 (
            .O(N__43003),
            .I(N__43000));
    InMux I__8909 (
            .O(N__43000),
            .I(N__42997));
    LocalMux I__8908 (
            .O(N__42997),
            .I(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ));
    CascadeMux I__8907 (
            .O(N__42994),
            .I(N__42991));
    InMux I__8906 (
            .O(N__42991),
            .I(N__42988));
    LocalMux I__8905 (
            .O(N__42988),
            .I(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ));
    CascadeMux I__8904 (
            .O(N__42985),
            .I(N__42982));
    InMux I__8903 (
            .O(N__42982),
            .I(N__42979));
    LocalMux I__8902 (
            .O(N__42979),
            .I(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ));
    InMux I__8901 (
            .O(N__42976),
            .I(N__42973));
    LocalMux I__8900 (
            .O(N__42973),
            .I(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ));
    InMux I__8899 (
            .O(N__42970),
            .I(\current_shift_inst.un4_control_input_1_cry_25 ));
    InMux I__8898 (
            .O(N__42967),
            .I(N__42964));
    LocalMux I__8897 (
            .O(N__42964),
            .I(N__42961));
    Span4Mux_h I__8896 (
            .O(N__42961),
            .I(N__42958));
    Odrv4 I__8895 (
            .O(N__42958),
            .I(\current_shift_inst.un4_control_input_1_axb_27 ));
    InMux I__8894 (
            .O(N__42955),
            .I(\current_shift_inst.un4_control_input_1_cry_26 ));
    InMux I__8893 (
            .O(N__42952),
            .I(N__42949));
    LocalMux I__8892 (
            .O(N__42949),
            .I(N__42946));
    Span4Mux_h I__8891 (
            .O(N__42946),
            .I(N__42943));
    Odrv4 I__8890 (
            .O(N__42943),
            .I(\current_shift_inst.un4_control_input_1_axb_28 ));
    InMux I__8889 (
            .O(N__42940),
            .I(\current_shift_inst.un4_control_input_1_cry_27 ));
    InMux I__8888 (
            .O(N__42937),
            .I(\current_shift_inst.un4_control_input_1_cry_28 ));
    InMux I__8887 (
            .O(N__42934),
            .I(\current_shift_inst.un4_control_input1_31 ));
    InMux I__8886 (
            .O(N__42931),
            .I(N__42928));
    LocalMux I__8885 (
            .O(N__42928),
            .I(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ));
    CascadeMux I__8884 (
            .O(N__42925),
            .I(N__42922));
    InMux I__8883 (
            .O(N__42922),
            .I(N__42919));
    LocalMux I__8882 (
            .O(N__42919),
            .I(N__42916));
    Odrv4 I__8881 (
            .O(N__42916),
            .I(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ));
    CascadeMux I__8880 (
            .O(N__42913),
            .I(N__42910));
    InMux I__8879 (
            .O(N__42910),
            .I(N__42907));
    LocalMux I__8878 (
            .O(N__42907),
            .I(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ));
    InMux I__8877 (
            .O(N__42904),
            .I(\current_shift_inst.un4_control_input_1_cry_17 ));
    InMux I__8876 (
            .O(N__42901),
            .I(N__42898));
    LocalMux I__8875 (
            .O(N__42898),
            .I(N__42895));
    Odrv12 I__8874 (
            .O(N__42895),
            .I(\current_shift_inst.un4_control_input_1_axb_19 ));
    InMux I__8873 (
            .O(N__42892),
            .I(\current_shift_inst.un4_control_input_1_cry_18 ));
    InMux I__8872 (
            .O(N__42889),
            .I(N__42886));
    LocalMux I__8871 (
            .O(N__42886),
            .I(N__42883));
    Span4Mux_h I__8870 (
            .O(N__42883),
            .I(N__42880));
    Odrv4 I__8869 (
            .O(N__42880),
            .I(\current_shift_inst.un4_control_input_1_axb_20 ));
    InMux I__8868 (
            .O(N__42877),
            .I(\current_shift_inst.un4_control_input_1_cry_19 ));
    InMux I__8867 (
            .O(N__42874),
            .I(N__42871));
    LocalMux I__8866 (
            .O(N__42871),
            .I(N__42868));
    Span4Mux_h I__8865 (
            .O(N__42868),
            .I(N__42865));
    Odrv4 I__8864 (
            .O(N__42865),
            .I(\current_shift_inst.un4_control_input_1_axb_21 ));
    InMux I__8863 (
            .O(N__42862),
            .I(\current_shift_inst.un4_control_input_1_cry_20 ));
    InMux I__8862 (
            .O(N__42859),
            .I(N__42856));
    LocalMux I__8861 (
            .O(N__42856),
            .I(N__42853));
    Span4Mux_h I__8860 (
            .O(N__42853),
            .I(N__42850));
    Odrv4 I__8859 (
            .O(N__42850),
            .I(\current_shift_inst.un4_control_input_1_axb_22 ));
    InMux I__8858 (
            .O(N__42847),
            .I(\current_shift_inst.un4_control_input_1_cry_21 ));
    InMux I__8857 (
            .O(N__42844),
            .I(N__42841));
    LocalMux I__8856 (
            .O(N__42841),
            .I(N__42838));
    Span4Mux_h I__8855 (
            .O(N__42838),
            .I(N__42835));
    Odrv4 I__8854 (
            .O(N__42835),
            .I(\current_shift_inst.un4_control_input_1_axb_23 ));
    InMux I__8853 (
            .O(N__42832),
            .I(\current_shift_inst.un4_control_input_1_cry_22 ));
    InMux I__8852 (
            .O(N__42829),
            .I(\current_shift_inst.un4_control_input_1_cry_23 ));
    InMux I__8851 (
            .O(N__42826),
            .I(bfn_16_16_0_));
    InMux I__8850 (
            .O(N__42823),
            .I(N__42820));
    LocalMux I__8849 (
            .O(N__42820),
            .I(\current_shift_inst.un4_control_input_1_axb_9 ));
    InMux I__8848 (
            .O(N__42817),
            .I(bfn_16_14_0_));
    InMux I__8847 (
            .O(N__42814),
            .I(N__42811));
    LocalMux I__8846 (
            .O(N__42811),
            .I(\current_shift_inst.un4_control_input_1_axb_10 ));
    InMux I__8845 (
            .O(N__42808),
            .I(\current_shift_inst.un4_control_input_1_cry_9 ));
    InMux I__8844 (
            .O(N__42805),
            .I(N__42802));
    LocalMux I__8843 (
            .O(N__42802),
            .I(N__42799));
    Span4Mux_h I__8842 (
            .O(N__42799),
            .I(N__42796));
    Odrv4 I__8841 (
            .O(N__42796),
            .I(\current_shift_inst.un4_control_input_1_axb_11 ));
    InMux I__8840 (
            .O(N__42793),
            .I(\current_shift_inst.un4_control_input_1_cry_10 ));
    InMux I__8839 (
            .O(N__42790),
            .I(N__42787));
    LocalMux I__8838 (
            .O(N__42787),
            .I(N__42784));
    Span4Mux_v I__8837 (
            .O(N__42784),
            .I(N__42781));
    Odrv4 I__8836 (
            .O(N__42781),
            .I(\current_shift_inst.un4_control_input_1_axb_12 ));
    InMux I__8835 (
            .O(N__42778),
            .I(\current_shift_inst.un4_control_input_1_cry_11 ));
    InMux I__8834 (
            .O(N__42775),
            .I(N__42772));
    LocalMux I__8833 (
            .O(N__42772),
            .I(\current_shift_inst.un4_control_input_1_axb_13 ));
    InMux I__8832 (
            .O(N__42769),
            .I(\current_shift_inst.un4_control_input_1_cry_12 ));
    InMux I__8831 (
            .O(N__42766),
            .I(N__42763));
    LocalMux I__8830 (
            .O(N__42763),
            .I(\current_shift_inst.un4_control_input_1_axb_14 ));
    InMux I__8829 (
            .O(N__42760),
            .I(\current_shift_inst.un4_control_input_1_cry_13 ));
    InMux I__8828 (
            .O(N__42757),
            .I(N__42754));
    LocalMux I__8827 (
            .O(N__42754),
            .I(N__42751));
    Span4Mux_h I__8826 (
            .O(N__42751),
            .I(N__42748));
    Odrv4 I__8825 (
            .O(N__42748),
            .I(\current_shift_inst.un4_control_input_1_axb_15 ));
    InMux I__8824 (
            .O(N__42745),
            .I(\current_shift_inst.un4_control_input_1_cry_14 ));
    InMux I__8823 (
            .O(N__42742),
            .I(N__42739));
    LocalMux I__8822 (
            .O(N__42739),
            .I(\current_shift_inst.un4_control_input_1_axb_16 ));
    InMux I__8821 (
            .O(N__42736),
            .I(\current_shift_inst.un4_control_input_1_cry_15 ));
    InMux I__8820 (
            .O(N__42733),
            .I(N__42730));
    LocalMux I__8819 (
            .O(N__42730),
            .I(N__42727));
    Odrv12 I__8818 (
            .O(N__42727),
            .I(\current_shift_inst.un4_control_input_1_axb_17 ));
    InMux I__8817 (
            .O(N__42724),
            .I(bfn_16_15_0_));
    InMux I__8816 (
            .O(N__42721),
            .I(N__42718));
    LocalMux I__8815 (
            .O(N__42718),
            .I(\current_shift_inst.un4_control_input_1_axb_1 ));
    InMux I__8814 (
            .O(N__42715),
            .I(N__42712));
    LocalMux I__8813 (
            .O(N__42712),
            .I(\current_shift_inst.un4_control_input_1_axb_2 ));
    InMux I__8812 (
            .O(N__42709),
            .I(\current_shift_inst.un4_control_input_1_cry_1 ));
    InMux I__8811 (
            .O(N__42706),
            .I(N__42703));
    LocalMux I__8810 (
            .O(N__42703),
            .I(\current_shift_inst.un4_control_input_1_axb_3 ));
    InMux I__8809 (
            .O(N__42700),
            .I(\current_shift_inst.un4_control_input_1_cry_2 ));
    InMux I__8808 (
            .O(N__42697),
            .I(N__42694));
    LocalMux I__8807 (
            .O(N__42694),
            .I(\current_shift_inst.un4_control_input_1_axb_4 ));
    InMux I__8806 (
            .O(N__42691),
            .I(\current_shift_inst.un4_control_input_1_cry_3 ));
    InMux I__8805 (
            .O(N__42688),
            .I(N__42685));
    LocalMux I__8804 (
            .O(N__42685),
            .I(\current_shift_inst.un4_control_input_1_axb_5 ));
    InMux I__8803 (
            .O(N__42682),
            .I(\current_shift_inst.un4_control_input_1_cry_4 ));
    InMux I__8802 (
            .O(N__42679),
            .I(N__42676));
    LocalMux I__8801 (
            .O(N__42676),
            .I(\current_shift_inst.un4_control_input_1_axb_6 ));
    InMux I__8800 (
            .O(N__42673),
            .I(\current_shift_inst.un4_control_input_1_cry_5 ));
    InMux I__8799 (
            .O(N__42670),
            .I(N__42667));
    LocalMux I__8798 (
            .O(N__42667),
            .I(\current_shift_inst.un4_control_input_1_axb_7 ));
    InMux I__8797 (
            .O(N__42664),
            .I(\current_shift_inst.un4_control_input_1_cry_6 ));
    InMux I__8796 (
            .O(N__42661),
            .I(N__42658));
    LocalMux I__8795 (
            .O(N__42658),
            .I(N__42655));
    Span4Mux_h I__8794 (
            .O(N__42655),
            .I(N__42652));
    Odrv4 I__8793 (
            .O(N__42652),
            .I(\current_shift_inst.un4_control_input_1_axb_8 ));
    InMux I__8792 (
            .O(N__42649),
            .I(\current_shift_inst.un4_control_input_1_cry_7 ));
    InMux I__8791 (
            .O(N__42646),
            .I(N__42643));
    LocalMux I__8790 (
            .O(N__42643),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ));
    InMux I__8789 (
            .O(N__42640),
            .I(N__42636));
    InMux I__8788 (
            .O(N__42639),
            .I(N__42632));
    LocalMux I__8787 (
            .O(N__42636),
            .I(N__42627));
    InMux I__8786 (
            .O(N__42635),
            .I(N__42624));
    LocalMux I__8785 (
            .O(N__42632),
            .I(N__42621));
    InMux I__8784 (
            .O(N__42631),
            .I(N__42618));
    InMux I__8783 (
            .O(N__42630),
            .I(N__42615));
    Odrv4 I__8782 (
            .O(N__42627),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__8781 (
            .O(N__42624),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    Odrv12 I__8780 (
            .O(N__42621),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__8779 (
            .O(N__42618),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    LocalMux I__8778 (
            .O(N__42615),
            .I(elapsed_time_ns_1_RNI04EN9_0_31));
    InMux I__8777 (
            .O(N__42604),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ));
    InMux I__8776 (
            .O(N__42601),
            .I(N__42598));
    LocalMux I__8775 (
            .O(N__42598),
            .I(N__42594));
    InMux I__8774 (
            .O(N__42597),
            .I(N__42591));
    Span4Mux_h I__8773 (
            .O(N__42594),
            .I(N__42588));
    LocalMux I__8772 (
            .O(N__42591),
            .I(N__42585));
    Odrv4 I__8771 (
            .O(N__42588),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_28));
    Odrv12 I__8770 (
            .O(N__42585),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_28));
    InMux I__8769 (
            .O(N__42580),
            .I(N__42577));
    LocalMux I__8768 (
            .O(N__42577),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ));
    CascadeMux I__8767 (
            .O(N__42574),
            .I(N__42571));
    InMux I__8766 (
            .O(N__42571),
            .I(N__42568));
    LocalMux I__8765 (
            .O(N__42568),
            .I(N__42565));
    Span4Mux_v I__8764 (
            .O(N__42565),
            .I(N__42562));
    Odrv4 I__8763 (
            .O(N__42562),
            .I(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ));
    CascadeMux I__8762 (
            .O(N__42559),
            .I(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ));
    InMux I__8761 (
            .O(N__42556),
            .I(N__42552));
    CascadeMux I__8760 (
            .O(N__42555),
            .I(N__42549));
    LocalMux I__8759 (
            .O(N__42552),
            .I(N__42546));
    InMux I__8758 (
            .O(N__42549),
            .I(N__42543));
    Span4Mux_v I__8757 (
            .O(N__42546),
            .I(N__42540));
    LocalMux I__8756 (
            .O(N__42543),
            .I(N__42537));
    Span4Mux_h I__8755 (
            .O(N__42540),
            .I(N__42532));
    Span4Mux_v I__8754 (
            .O(N__42537),
            .I(N__42532));
    Odrv4 I__8753 (
            .O(N__42532),
            .I(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ));
    InMux I__8752 (
            .O(N__42529),
            .I(N__42526));
    LocalMux I__8751 (
            .O(N__42526),
            .I(N__42522));
    InMux I__8750 (
            .O(N__42525),
            .I(N__42518));
    Span4Mux_h I__8749 (
            .O(N__42522),
            .I(N__42515));
    InMux I__8748 (
            .O(N__42521),
            .I(N__42512));
    LocalMux I__8747 (
            .O(N__42518),
            .I(N__42509));
    Odrv4 I__8746 (
            .O(N__42515),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    LocalMux I__8745 (
            .O(N__42512),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    Odrv12 I__8744 (
            .O(N__42509),
            .I(\current_shift_inst.timer_s1.counterZ0Z_0 ));
    InMux I__8743 (
            .O(N__42502),
            .I(N__42499));
    LocalMux I__8742 (
            .O(N__42499),
            .I(N__42495));
    InMux I__8741 (
            .O(N__42498),
            .I(N__42492));
    Odrv4 I__8740 (
            .O(N__42495),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ));
    LocalMux I__8739 (
            .O(N__42492),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ));
    InMux I__8738 (
            .O(N__42487),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ));
    InMux I__8737 (
            .O(N__42484),
            .I(N__42480));
    InMux I__8736 (
            .O(N__42483),
            .I(N__42477));
    LocalMux I__8735 (
            .O(N__42480),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ));
    LocalMux I__8734 (
            .O(N__42477),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ));
    InMux I__8733 (
            .O(N__42472),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ));
    InMux I__8732 (
            .O(N__42469),
            .I(N__42466));
    LocalMux I__8731 (
            .O(N__42466),
            .I(N__42463));
    Odrv4 I__8730 (
            .O(N__42463),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ));
    InMux I__8729 (
            .O(N__42460),
            .I(N__42456));
    InMux I__8728 (
            .O(N__42459),
            .I(N__42453));
    LocalMux I__8727 (
            .O(N__42456),
            .I(N__42450));
    LocalMux I__8726 (
            .O(N__42453),
            .I(N__42447));
    Odrv4 I__8725 (
            .O(N__42450),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ));
    Odrv4 I__8724 (
            .O(N__42447),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ));
    InMux I__8723 (
            .O(N__42442),
            .I(bfn_16_11_0_));
    InMux I__8722 (
            .O(N__42439),
            .I(N__42435));
    InMux I__8721 (
            .O(N__42438),
            .I(N__42432));
    LocalMux I__8720 (
            .O(N__42435),
            .I(N__42427));
    LocalMux I__8719 (
            .O(N__42432),
            .I(N__42427));
    Odrv4 I__8718 (
            .O(N__42427),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ));
    InMux I__8717 (
            .O(N__42424),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ));
    InMux I__8716 (
            .O(N__42421),
            .I(N__42417));
    InMux I__8715 (
            .O(N__42420),
            .I(N__42414));
    LocalMux I__8714 (
            .O(N__42417),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ));
    LocalMux I__8713 (
            .O(N__42414),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ));
    InMux I__8712 (
            .O(N__42409),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ));
    InMux I__8711 (
            .O(N__42406),
            .I(N__42402));
    InMux I__8710 (
            .O(N__42405),
            .I(N__42399));
    LocalMux I__8709 (
            .O(N__42402),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ));
    LocalMux I__8708 (
            .O(N__42399),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ));
    InMux I__8707 (
            .O(N__42394),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ));
    InMux I__8706 (
            .O(N__42391),
            .I(N__42388));
    LocalMux I__8705 (
            .O(N__42388),
            .I(N__42385));
    Odrv12 I__8704 (
            .O(N__42385),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ));
    InMux I__8703 (
            .O(N__42382),
            .I(N__42378));
    InMux I__8702 (
            .O(N__42381),
            .I(N__42375));
    LocalMux I__8701 (
            .O(N__42378),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ));
    LocalMux I__8700 (
            .O(N__42375),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ));
    InMux I__8699 (
            .O(N__42370),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ));
    InMux I__8698 (
            .O(N__42367),
            .I(N__42364));
    LocalMux I__8697 (
            .O(N__42364),
            .I(N__42361));
    Span4Mux_h I__8696 (
            .O(N__42361),
            .I(N__42358));
    Odrv4 I__8695 (
            .O(N__42358),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ));
    InMux I__8694 (
            .O(N__42355),
            .I(N__42351));
    InMux I__8693 (
            .O(N__42354),
            .I(N__42348));
    LocalMux I__8692 (
            .O(N__42351),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ));
    LocalMux I__8691 (
            .O(N__42348),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ));
    InMux I__8690 (
            .O(N__42343),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ));
    InMux I__8689 (
            .O(N__42340),
            .I(N__42336));
    InMux I__8688 (
            .O(N__42339),
            .I(N__42333));
    LocalMux I__8687 (
            .O(N__42336),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ));
    LocalMux I__8686 (
            .O(N__42333),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ));
    InMux I__8685 (
            .O(N__42328),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ));
    InMux I__8684 (
            .O(N__42325),
            .I(N__42321));
    InMux I__8683 (
            .O(N__42324),
            .I(N__42318));
    LocalMux I__8682 (
            .O(N__42321),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ));
    LocalMux I__8681 (
            .O(N__42318),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ));
    InMux I__8680 (
            .O(N__42313),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ));
    InMux I__8679 (
            .O(N__42310),
            .I(N__42306));
    InMux I__8678 (
            .O(N__42309),
            .I(N__42303));
    LocalMux I__8677 (
            .O(N__42306),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ));
    LocalMux I__8676 (
            .O(N__42303),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ));
    InMux I__8675 (
            .O(N__42298),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ));
    InMux I__8674 (
            .O(N__42295),
            .I(N__42291));
    InMux I__8673 (
            .O(N__42294),
            .I(N__42288));
    LocalMux I__8672 (
            .O(N__42291),
            .I(N__42285));
    LocalMux I__8671 (
            .O(N__42288),
            .I(N__42282));
    Odrv4 I__8670 (
            .O(N__42285),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ));
    Odrv4 I__8669 (
            .O(N__42282),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ));
    InMux I__8668 (
            .O(N__42277),
            .I(bfn_16_10_0_));
    InMux I__8667 (
            .O(N__42274),
            .I(N__42270));
    InMux I__8666 (
            .O(N__42273),
            .I(N__42267));
    LocalMux I__8665 (
            .O(N__42270),
            .I(N__42262));
    LocalMux I__8664 (
            .O(N__42267),
            .I(N__42262));
    Odrv4 I__8663 (
            .O(N__42262),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ));
    InMux I__8662 (
            .O(N__42259),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ));
    InMux I__8661 (
            .O(N__42256),
            .I(N__42252));
    InMux I__8660 (
            .O(N__42255),
            .I(N__42249));
    LocalMux I__8659 (
            .O(N__42252),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ));
    LocalMux I__8658 (
            .O(N__42249),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ));
    InMux I__8657 (
            .O(N__42244),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ));
    InMux I__8656 (
            .O(N__42241),
            .I(N__42237));
    InMux I__8655 (
            .O(N__42240),
            .I(N__42234));
    LocalMux I__8654 (
            .O(N__42237),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ));
    LocalMux I__8653 (
            .O(N__42234),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ));
    InMux I__8652 (
            .O(N__42229),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ));
    InMux I__8651 (
            .O(N__42226),
            .I(N__42223));
    LocalMux I__8650 (
            .O(N__42223),
            .I(N__42220));
    Span4Mux_h I__8649 (
            .O(N__42220),
            .I(N__42216));
    InMux I__8648 (
            .O(N__42219),
            .I(N__42213));
    Span4Mux_h I__8647 (
            .O(N__42216),
            .I(N__42210));
    LocalMux I__8646 (
            .O(N__42213),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ));
    Odrv4 I__8645 (
            .O(N__42210),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ));
    InMux I__8644 (
            .O(N__42205),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ));
    InMux I__8643 (
            .O(N__42202),
            .I(N__42199));
    LocalMux I__8642 (
            .O(N__42199),
            .I(N__42196));
    Span4Mux_h I__8641 (
            .O(N__42196),
            .I(N__42193));
    Odrv4 I__8640 (
            .O(N__42193),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ));
    InMux I__8639 (
            .O(N__42190),
            .I(N__42186));
    InMux I__8638 (
            .O(N__42189),
            .I(N__42183));
    LocalMux I__8637 (
            .O(N__42186),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ));
    LocalMux I__8636 (
            .O(N__42183),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ));
    InMux I__8635 (
            .O(N__42178),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ));
    InMux I__8634 (
            .O(N__42175),
            .I(N__42171));
    InMux I__8633 (
            .O(N__42174),
            .I(N__42168));
    LocalMux I__8632 (
            .O(N__42171),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ));
    LocalMux I__8631 (
            .O(N__42168),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ));
    InMux I__8630 (
            .O(N__42163),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ));
    InMux I__8629 (
            .O(N__42160),
            .I(N__42156));
    InMux I__8628 (
            .O(N__42159),
            .I(N__42153));
    LocalMux I__8627 (
            .O(N__42156),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ));
    LocalMux I__8626 (
            .O(N__42153),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ));
    InMux I__8625 (
            .O(N__42148),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ));
    InMux I__8624 (
            .O(N__42145),
            .I(N__42141));
    InMux I__8623 (
            .O(N__42144),
            .I(N__42138));
    LocalMux I__8622 (
            .O(N__42141),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ));
    LocalMux I__8621 (
            .O(N__42138),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ));
    InMux I__8620 (
            .O(N__42133),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ));
    InMux I__8619 (
            .O(N__42130),
            .I(N__42126));
    InMux I__8618 (
            .O(N__42129),
            .I(N__42123));
    LocalMux I__8617 (
            .O(N__42126),
            .I(N__42120));
    LocalMux I__8616 (
            .O(N__42123),
            .I(N__42117));
    Odrv4 I__8615 (
            .O(N__42120),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ));
    Odrv4 I__8614 (
            .O(N__42117),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ));
    InMux I__8613 (
            .O(N__42112),
            .I(bfn_16_9_0_));
    InMux I__8612 (
            .O(N__42109),
            .I(N__42105));
    InMux I__8611 (
            .O(N__42108),
            .I(N__42102));
    LocalMux I__8610 (
            .O(N__42105),
            .I(N__42097));
    LocalMux I__8609 (
            .O(N__42102),
            .I(N__42097));
    Span4Mux_v I__8608 (
            .O(N__42097),
            .I(N__42094));
    Odrv4 I__8607 (
            .O(N__42094),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ));
    InMux I__8606 (
            .O(N__42091),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ));
    InMux I__8605 (
            .O(N__42088),
            .I(N__42084));
    InMux I__8604 (
            .O(N__42087),
            .I(N__42081));
    LocalMux I__8603 (
            .O(N__42084),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ));
    LocalMux I__8602 (
            .O(N__42081),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ));
    InMux I__8601 (
            .O(N__42076),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ));
    InMux I__8600 (
            .O(N__42073),
            .I(N__42069));
    InMux I__8599 (
            .O(N__42072),
            .I(N__42066));
    LocalMux I__8598 (
            .O(N__42069),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ));
    LocalMux I__8597 (
            .O(N__42066),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ));
    InMux I__8596 (
            .O(N__42061),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ));
    InMux I__8595 (
            .O(N__42058),
            .I(N__42054));
    InMux I__8594 (
            .O(N__42057),
            .I(N__42051));
    LocalMux I__8593 (
            .O(N__42054),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ));
    LocalMux I__8592 (
            .O(N__42051),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ));
    InMux I__8591 (
            .O(N__42046),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ));
    CEMux I__8590 (
            .O(N__42043),
            .I(N__42040));
    LocalMux I__8589 (
            .O(N__42040),
            .I(N__42034));
    CEMux I__8588 (
            .O(N__42039),
            .I(N__42029));
    CEMux I__8587 (
            .O(N__42038),
            .I(N__42026));
    CEMux I__8586 (
            .O(N__42037),
            .I(N__42023));
    Span4Mux_h I__8585 (
            .O(N__42034),
            .I(N__42019));
    CEMux I__8584 (
            .O(N__42033),
            .I(N__42016));
    CEMux I__8583 (
            .O(N__42032),
            .I(N__42013));
    LocalMux I__8582 (
            .O(N__42029),
            .I(N__42010));
    LocalMux I__8581 (
            .O(N__42026),
            .I(N__42007));
    LocalMux I__8580 (
            .O(N__42023),
            .I(N__42004));
    CEMux I__8579 (
            .O(N__42022),
            .I(N__42001));
    Span4Mux_v I__8578 (
            .O(N__42019),
            .I(N__41996));
    LocalMux I__8577 (
            .O(N__42016),
            .I(N__41996));
    LocalMux I__8576 (
            .O(N__42013),
            .I(N__41993));
    Span4Mux_h I__8575 (
            .O(N__42010),
            .I(N__41990));
    Span4Mux_h I__8574 (
            .O(N__42007),
            .I(N__41983));
    Span4Mux_v I__8573 (
            .O(N__42004),
            .I(N__41983));
    LocalMux I__8572 (
            .O(N__42001),
            .I(N__41983));
    Span4Mux_h I__8571 (
            .O(N__41996),
            .I(N__41978));
    Span4Mux_h I__8570 (
            .O(N__41993),
            .I(N__41978));
    Span4Mux_v I__8569 (
            .O(N__41990),
            .I(N__41973));
    Span4Mux_v I__8568 (
            .O(N__41983),
            .I(N__41973));
    Odrv4 I__8567 (
            .O(N__41978),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__8566 (
            .O(N__41973),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ));
    CascadeMux I__8565 (
            .O(N__41968),
            .I(elapsed_time_ns_1_RNI04EN9_0_31_cascade_));
    InMux I__8564 (
            .O(N__41965),
            .I(N__41962));
    LocalMux I__8563 (
            .O(N__41962),
            .I(N__41959));
    Span12Mux_s6_v I__8562 (
            .O(N__41959),
            .I(N__41956));
    Odrv12 I__8561 (
            .O(N__41956),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ));
    CEMux I__8560 (
            .O(N__41953),
            .I(N__41949));
    CEMux I__8559 (
            .O(N__41952),
            .I(N__41944));
    LocalMux I__8558 (
            .O(N__41949),
            .I(N__41941));
    CEMux I__8557 (
            .O(N__41948),
            .I(N__41938));
    CEMux I__8556 (
            .O(N__41947),
            .I(N__41935));
    LocalMux I__8555 (
            .O(N__41944),
            .I(N__41929));
    Span4Mux_h I__8554 (
            .O(N__41941),
            .I(N__41922));
    LocalMux I__8553 (
            .O(N__41938),
            .I(N__41922));
    LocalMux I__8552 (
            .O(N__41935),
            .I(N__41922));
    CEMux I__8551 (
            .O(N__41934),
            .I(N__41919));
    CEMux I__8550 (
            .O(N__41933),
            .I(N__41916));
    CEMux I__8549 (
            .O(N__41932),
            .I(N__41912));
    Span4Mux_h I__8548 (
            .O(N__41929),
            .I(N__41905));
    Span4Mux_v I__8547 (
            .O(N__41922),
            .I(N__41905));
    LocalMux I__8546 (
            .O(N__41919),
            .I(N__41905));
    LocalMux I__8545 (
            .O(N__41916),
            .I(N__41902));
    CEMux I__8544 (
            .O(N__41915),
            .I(N__41899));
    LocalMux I__8543 (
            .O(N__41912),
            .I(N__41896));
    Span4Mux_h I__8542 (
            .O(N__41905),
            .I(N__41893));
    Span4Mux_h I__8541 (
            .O(N__41902),
            .I(N__41890));
    LocalMux I__8540 (
            .O(N__41899),
            .I(N__41887));
    Span4Mux_h I__8539 (
            .O(N__41896),
            .I(N__41884));
    Odrv4 I__8538 (
            .O(N__41893),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__8537 (
            .O(N__41890),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__8536 (
            .O(N__41887),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    Odrv4 I__8535 (
            .O(N__41884),
            .I(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ));
    CascadeMux I__8534 (
            .O(N__41875),
            .I(N__41872));
    InMux I__8533 (
            .O(N__41872),
            .I(N__41869));
    LocalMux I__8532 (
            .O(N__41869),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ));
    InMux I__8531 (
            .O(N__41866),
            .I(N__41863));
    LocalMux I__8530 (
            .O(N__41863),
            .I(N__41859));
    InMux I__8529 (
            .O(N__41862),
            .I(N__41856));
    Span4Mux_h I__8528 (
            .O(N__41859),
            .I(N__41853));
    LocalMux I__8527 (
            .O(N__41856),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    Odrv4 I__8526 (
            .O(N__41853),
            .I(elapsed_time_ns_1_RNIE03T9_0_2));
    InMux I__8525 (
            .O(N__41848),
            .I(N__41845));
    LocalMux I__8524 (
            .O(N__41845),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ));
    InMux I__8523 (
            .O(N__41842),
            .I(N__41839));
    LocalMux I__8522 (
            .O(N__41839),
            .I(N__41836));
    Odrv4 I__8521 (
            .O(N__41836),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ));
    InMux I__8520 (
            .O(N__41833),
            .I(N__41828));
    CascadeMux I__8519 (
            .O(N__41832),
            .I(N__41825));
    InMux I__8518 (
            .O(N__41831),
            .I(N__41822));
    LocalMux I__8517 (
            .O(N__41828),
            .I(N__41819));
    InMux I__8516 (
            .O(N__41825),
            .I(N__41816));
    LocalMux I__8515 (
            .O(N__41822),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    Odrv4 I__8514 (
            .O(N__41819),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    LocalMux I__8513 (
            .O(N__41816),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ));
    InMux I__8512 (
            .O(N__41809),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ));
    InMux I__8511 (
            .O(N__41806),
            .I(N__41803));
    LocalMux I__8510 (
            .O(N__41803),
            .I(N__41800));
    Odrv4 I__8509 (
            .O(N__41800),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ));
    InMux I__8508 (
            .O(N__41797),
            .I(N__41793));
    InMux I__8507 (
            .O(N__41796),
            .I(N__41790));
    LocalMux I__8506 (
            .O(N__41793),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ));
    LocalMux I__8505 (
            .O(N__41790),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ));
    InMux I__8504 (
            .O(N__41785),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ));
    InMux I__8503 (
            .O(N__41782),
            .I(N__41778));
    InMux I__8502 (
            .O(N__41781),
            .I(N__41775));
    LocalMux I__8501 (
            .O(N__41778),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ));
    LocalMux I__8500 (
            .O(N__41775),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ));
    InMux I__8499 (
            .O(N__41770),
            .I(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ));
    InMux I__8498 (
            .O(N__41767),
            .I(N__41764));
    LocalMux I__8497 (
            .O(N__41764),
            .I(\current_shift_inst.control_input_axb_29 ));
    InMux I__8496 (
            .O(N__41761),
            .I(N__41757));
    InMux I__8495 (
            .O(N__41760),
            .I(N__41754));
    LocalMux I__8494 (
            .O(N__41757),
            .I(N__41751));
    LocalMux I__8493 (
            .O(N__41754),
            .I(N__41748));
    Span4Mux_h I__8492 (
            .O(N__41751),
            .I(N__41745));
    Odrv4 I__8491 (
            .O(N__41748),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    Odrv4 I__8490 (
            .O(N__41745),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ));
    InMux I__8489 (
            .O(N__41740),
            .I(N__41736));
    InMux I__8488 (
            .O(N__41739),
            .I(N__41733));
    LocalMux I__8487 (
            .O(N__41736),
            .I(N__41730));
    LocalMux I__8486 (
            .O(N__41733),
            .I(N__41727));
    Span4Mux_h I__8485 (
            .O(N__41730),
            .I(N__41724));
    Odrv12 I__8484 (
            .O(N__41727),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    Odrv4 I__8483 (
            .O(N__41724),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ));
    CascadeMux I__8482 (
            .O(N__41719),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ));
    InMux I__8481 (
            .O(N__41716),
            .I(N__41710));
    InMux I__8480 (
            .O(N__41715),
            .I(N__41710));
    LocalMux I__8479 (
            .O(N__41710),
            .I(N__41707));
    Odrv4 I__8478 (
            .O(N__41707),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ));
    InMux I__8477 (
            .O(N__41704),
            .I(N__41700));
    InMux I__8476 (
            .O(N__41703),
            .I(N__41697));
    LocalMux I__8475 (
            .O(N__41700),
            .I(N__41692));
    LocalMux I__8474 (
            .O(N__41697),
            .I(N__41692));
    Odrv12 I__8473 (
            .O(N__41692),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ));
    InMux I__8472 (
            .O(N__41689),
            .I(N__41683));
    InMux I__8471 (
            .O(N__41688),
            .I(N__41683));
    LocalMux I__8470 (
            .O(N__41683),
            .I(N__41680));
    Odrv4 I__8469 (
            .O(N__41680),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ));
    CascadeMux I__8468 (
            .O(N__41677),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ));
    InMux I__8467 (
            .O(N__41674),
            .I(N__41671));
    LocalMux I__8466 (
            .O(N__41671),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ));
    InMux I__8465 (
            .O(N__41668),
            .I(N__41665));
    LocalMux I__8464 (
            .O(N__41665),
            .I(\current_shift_inst.control_input_axb_18 ));
    InMux I__8463 (
            .O(N__41662),
            .I(N__41658));
    InMux I__8462 (
            .O(N__41661),
            .I(N__41655));
    LocalMux I__8461 (
            .O(N__41658),
            .I(N__41650));
    LocalMux I__8460 (
            .O(N__41655),
            .I(N__41650));
    Odrv12 I__8459 (
            .O(N__41650),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ));
    InMux I__8458 (
            .O(N__41647),
            .I(N__41643));
    InMux I__8457 (
            .O(N__41646),
            .I(N__41640));
    LocalMux I__8456 (
            .O(N__41643),
            .I(N__41635));
    LocalMux I__8455 (
            .O(N__41640),
            .I(N__41635));
    Odrv4 I__8454 (
            .O(N__41635),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ));
    CascadeMux I__8453 (
            .O(N__41632),
            .I(N__41629));
    InMux I__8452 (
            .O(N__41629),
            .I(N__41626));
    LocalMux I__8451 (
            .O(N__41626),
            .I(N__41622));
    InMux I__8450 (
            .O(N__41625),
            .I(N__41619));
    Span4Mux_h I__8449 (
            .O(N__41622),
            .I(N__41614));
    LocalMux I__8448 (
            .O(N__41619),
            .I(N__41614));
    Odrv4 I__8447 (
            .O(N__41614),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ));
    InMux I__8446 (
            .O(N__41611),
            .I(N__41608));
    LocalMux I__8445 (
            .O(N__41608),
            .I(N__41604));
    InMux I__8444 (
            .O(N__41607),
            .I(N__41601));
    Span4Mux_h I__8443 (
            .O(N__41604),
            .I(N__41598));
    LocalMux I__8442 (
            .O(N__41601),
            .I(N__41595));
    Odrv4 I__8441 (
            .O(N__41598),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    Odrv12 I__8440 (
            .O(N__41595),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ));
    InMux I__8439 (
            .O(N__41590),
            .I(N__41587));
    LocalMux I__8438 (
            .O(N__41587),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ));
    InMux I__8437 (
            .O(N__41584),
            .I(N__41581));
    LocalMux I__8436 (
            .O(N__41581),
            .I(N__41578));
    Span4Mux_h I__8435 (
            .O(N__41578),
            .I(N__41575));
    Odrv4 I__8434 (
            .O(N__41575),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ));
    CascadeMux I__8433 (
            .O(N__41572),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ));
    InMux I__8432 (
            .O(N__41569),
            .I(N__41566));
    LocalMux I__8431 (
            .O(N__41566),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ));
    InMux I__8430 (
            .O(N__41563),
            .I(N__41560));
    LocalMux I__8429 (
            .O(N__41560),
            .I(N__41556));
    InMux I__8428 (
            .O(N__41559),
            .I(N__41553));
    Span4Mux_h I__8427 (
            .O(N__41556),
            .I(N__41550));
    LocalMux I__8426 (
            .O(N__41553),
            .I(N__41547));
    Odrv4 I__8425 (
            .O(N__41550),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_15));
    Odrv4 I__8424 (
            .O(N__41547),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_15));
    InMux I__8423 (
            .O(N__41542),
            .I(N__41539));
    LocalMux I__8422 (
            .O(N__41539),
            .I(N__41536));
    Odrv4 I__8421 (
            .O(N__41536),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ));
    InMux I__8420 (
            .O(N__41533),
            .I(N__41530));
    LocalMux I__8419 (
            .O(N__41530),
            .I(\current_shift_inst.control_input_axb_7 ));
    InMux I__8418 (
            .O(N__41527),
            .I(N__41524));
    LocalMux I__8417 (
            .O(N__41524),
            .I(\current_shift_inst.control_input_axb_13 ));
    InMux I__8416 (
            .O(N__41521),
            .I(N__41518));
    LocalMux I__8415 (
            .O(N__41518),
            .I(\current_shift_inst.control_input_axb_21 ));
    InMux I__8414 (
            .O(N__41515),
            .I(N__41512));
    LocalMux I__8413 (
            .O(N__41512),
            .I(\current_shift_inst.control_input_axb_26 ));
    InMux I__8412 (
            .O(N__41509),
            .I(N__41506));
    LocalMux I__8411 (
            .O(N__41506),
            .I(\current_shift_inst.control_input_axb_22 ));
    InMux I__8410 (
            .O(N__41503),
            .I(N__41500));
    LocalMux I__8409 (
            .O(N__41500),
            .I(\current_shift_inst.control_input_axb_17 ));
    InMux I__8408 (
            .O(N__41497),
            .I(N__41494));
    LocalMux I__8407 (
            .O(N__41494),
            .I(\current_shift_inst.control_input_axb_16 ));
    InMux I__8406 (
            .O(N__41491),
            .I(N__41488));
    LocalMux I__8405 (
            .O(N__41488),
            .I(\current_shift_inst.control_input_axb_25 ));
    InMux I__8404 (
            .O(N__41485),
            .I(N__41482));
    LocalMux I__8403 (
            .O(N__41482),
            .I(\current_shift_inst.control_input_axb_27 ));
    CascadeMux I__8402 (
            .O(N__41479),
            .I(N__41476));
    InMux I__8401 (
            .O(N__41476),
            .I(N__41473));
    LocalMux I__8400 (
            .O(N__41473),
            .I(N__41470));
    Span4Mux_v I__8399 (
            .O(N__41470),
            .I(N__41467));
    Odrv4 I__8398 (
            .O(N__41467),
            .I(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ));
    InMux I__8397 (
            .O(N__41464),
            .I(\current_shift_inst.un10_control_input_cry_30 ));
    InMux I__8396 (
            .O(N__41461),
            .I(N__41458));
    LocalMux I__8395 (
            .O(N__41458),
            .I(\current_shift_inst.control_input_axb_1 ));
    InMux I__8394 (
            .O(N__41455),
            .I(N__41452));
    LocalMux I__8393 (
            .O(N__41452),
            .I(\current_shift_inst.control_input_axb_2 ));
    InMux I__8392 (
            .O(N__41449),
            .I(N__41446));
    LocalMux I__8391 (
            .O(N__41446),
            .I(\current_shift_inst.control_input_axb_3 ));
    InMux I__8390 (
            .O(N__41443),
            .I(N__41440));
    LocalMux I__8389 (
            .O(N__41440),
            .I(\current_shift_inst.control_input_axb_4 ));
    InMux I__8388 (
            .O(N__41437),
            .I(N__41434));
    LocalMux I__8387 (
            .O(N__41434),
            .I(\current_shift_inst.control_input_axb_5 ));
    InMux I__8386 (
            .O(N__41431),
            .I(N__41428));
    LocalMux I__8385 (
            .O(N__41428),
            .I(\current_shift_inst.control_input_axb_6 ));
    InMux I__8384 (
            .O(N__41425),
            .I(N__41422));
    LocalMux I__8383 (
            .O(N__41422),
            .I(N__41419));
    Odrv12 I__8382 (
            .O(N__41419),
            .I(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ));
    CascadeMux I__8381 (
            .O(N__41416),
            .I(N__41413));
    InMux I__8380 (
            .O(N__41413),
            .I(N__41410));
    LocalMux I__8379 (
            .O(N__41410),
            .I(N__41407));
    Odrv4 I__8378 (
            .O(N__41407),
            .I(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ));
    InMux I__8377 (
            .O(N__41404),
            .I(N__41401));
    LocalMux I__8376 (
            .O(N__41401),
            .I(N__41398));
    Odrv4 I__8375 (
            .O(N__41398),
            .I(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ));
    CascadeMux I__8374 (
            .O(N__41395),
            .I(N__41392));
    InMux I__8373 (
            .O(N__41392),
            .I(N__41389));
    LocalMux I__8372 (
            .O(N__41389),
            .I(N__41386));
    Odrv4 I__8371 (
            .O(N__41386),
            .I(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ));
    CascadeMux I__8370 (
            .O(N__41383),
            .I(N__41380));
    InMux I__8369 (
            .O(N__41380),
            .I(N__41377));
    LocalMux I__8368 (
            .O(N__41377),
            .I(N__41374));
    Odrv4 I__8367 (
            .O(N__41374),
            .I(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ));
    InMux I__8366 (
            .O(N__41371),
            .I(N__41368));
    LocalMux I__8365 (
            .O(N__41368),
            .I(N__41365));
    Odrv12 I__8364 (
            .O(N__41365),
            .I(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ));
    CascadeMux I__8363 (
            .O(N__41362),
            .I(N__41359));
    InMux I__8362 (
            .O(N__41359),
            .I(N__41356));
    LocalMux I__8361 (
            .O(N__41356),
            .I(N__41353));
    Odrv4 I__8360 (
            .O(N__41353),
            .I(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ));
    InMux I__8359 (
            .O(N__41350),
            .I(N__41347));
    LocalMux I__8358 (
            .O(N__41347),
            .I(N__41344));
    Odrv4 I__8357 (
            .O(N__41344),
            .I(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ));
    CascadeMux I__8356 (
            .O(N__41341),
            .I(N__41338));
    InMux I__8355 (
            .O(N__41338),
            .I(N__41335));
    LocalMux I__8354 (
            .O(N__41335),
            .I(N__41332));
    Odrv4 I__8353 (
            .O(N__41332),
            .I(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ));
    CascadeMux I__8352 (
            .O(N__41329),
            .I(N__41326));
    InMux I__8351 (
            .O(N__41326),
            .I(N__41323));
    LocalMux I__8350 (
            .O(N__41323),
            .I(N__41320));
    Odrv4 I__8349 (
            .O(N__41320),
            .I(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ));
    InMux I__8348 (
            .O(N__41317),
            .I(N__41314));
    LocalMux I__8347 (
            .O(N__41314),
            .I(N__41311));
    Odrv12 I__8346 (
            .O(N__41311),
            .I(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ));
    CascadeMux I__8345 (
            .O(N__41308),
            .I(N__41305));
    InMux I__8344 (
            .O(N__41305),
            .I(N__41302));
    LocalMux I__8343 (
            .O(N__41302),
            .I(N__41299));
    Odrv12 I__8342 (
            .O(N__41299),
            .I(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ));
    CascadeMux I__8341 (
            .O(N__41296),
            .I(N__41293));
    InMux I__8340 (
            .O(N__41293),
            .I(N__41290));
    LocalMux I__8339 (
            .O(N__41290),
            .I(N__41287));
    Odrv12 I__8338 (
            .O(N__41287),
            .I(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ));
    InMux I__8337 (
            .O(N__41284),
            .I(N__41281));
    LocalMux I__8336 (
            .O(N__41281),
            .I(N__41278));
    Odrv12 I__8335 (
            .O(N__41278),
            .I(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ));
    InMux I__8334 (
            .O(N__41275),
            .I(N__41272));
    LocalMux I__8333 (
            .O(N__41272),
            .I(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ));
    InMux I__8332 (
            .O(N__41269),
            .I(N__41265));
    InMux I__8331 (
            .O(N__41268),
            .I(N__41262));
    LocalMux I__8330 (
            .O(N__41265),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    LocalMux I__8329 (
            .O(N__41262),
            .I(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ));
    InMux I__8328 (
            .O(N__41257),
            .I(N__41253));
    InMux I__8327 (
            .O(N__41256),
            .I(N__41250));
    LocalMux I__8326 (
            .O(N__41253),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    LocalMux I__8325 (
            .O(N__41250),
            .I(elapsed_time_ns_1_RNIF13T9_0_3));
    InMux I__8324 (
            .O(N__41245),
            .I(N__41240));
    InMux I__8323 (
            .O(N__41244),
            .I(N__41237));
    InMux I__8322 (
            .O(N__41243),
            .I(N__41234));
    LocalMux I__8321 (
            .O(N__41240),
            .I(N__41231));
    LocalMux I__8320 (
            .O(N__41237),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    LocalMux I__8319 (
            .O(N__41234),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    Odrv12 I__8318 (
            .O(N__41231),
            .I(\current_shift_inst.timer_s1.counterZ0Z_1 ));
    InMux I__8317 (
            .O(N__41224),
            .I(N__41221));
    LocalMux I__8316 (
            .O(N__41221),
            .I(N__41218));
    Span4Mux_h I__8315 (
            .O(N__41218),
            .I(N__41214));
    InMux I__8314 (
            .O(N__41217),
            .I(N__41211));
    Odrv4 I__8313 (
            .O(N__41214),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_21));
    LocalMux I__8312 (
            .O(N__41211),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_21));
    InMux I__8311 (
            .O(N__41206),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ));
    InMux I__8310 (
            .O(N__41203),
            .I(N__41200));
    LocalMux I__8309 (
            .O(N__41200),
            .I(N__41197));
    Span4Mux_h I__8308 (
            .O(N__41197),
            .I(N__41193));
    InMux I__8307 (
            .O(N__41196),
            .I(N__41190));
    Odrv4 I__8306 (
            .O(N__41193),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_22));
    LocalMux I__8305 (
            .O(N__41190),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_22));
    InMux I__8304 (
            .O(N__41185),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ));
    InMux I__8303 (
            .O(N__41182),
            .I(N__41179));
    LocalMux I__8302 (
            .O(N__41179),
            .I(N__41176));
    Span4Mux_h I__8301 (
            .O(N__41176),
            .I(N__41172));
    InMux I__8300 (
            .O(N__41175),
            .I(N__41169));
    Odrv4 I__8299 (
            .O(N__41172),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_23));
    LocalMux I__8298 (
            .O(N__41169),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_23));
    InMux I__8297 (
            .O(N__41164),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ));
    InMux I__8296 (
            .O(N__41161),
            .I(N__41158));
    LocalMux I__8295 (
            .O(N__41158),
            .I(N__41154));
    InMux I__8294 (
            .O(N__41157),
            .I(N__41151));
    Odrv12 I__8293 (
            .O(N__41154),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_24));
    LocalMux I__8292 (
            .O(N__41151),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_24));
    InMux I__8291 (
            .O(N__41146),
            .I(bfn_15_10_0_));
    InMux I__8290 (
            .O(N__41143),
            .I(N__41140));
    LocalMux I__8289 (
            .O(N__41140),
            .I(N__41137));
    Span12Mux_s9_v I__8288 (
            .O(N__41137),
            .I(N__41133));
    InMux I__8287 (
            .O(N__41136),
            .I(N__41130));
    Odrv12 I__8286 (
            .O(N__41133),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_25));
    LocalMux I__8285 (
            .O(N__41130),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_25));
    InMux I__8284 (
            .O(N__41125),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ));
    InMux I__8283 (
            .O(N__41122),
            .I(N__41119));
    LocalMux I__8282 (
            .O(N__41119),
            .I(N__41115));
    InMux I__8281 (
            .O(N__41118),
            .I(N__41112));
    Odrv4 I__8280 (
            .O(N__41115),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_26));
    LocalMux I__8279 (
            .O(N__41112),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_26));
    InMux I__8278 (
            .O(N__41107),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ));
    InMux I__8277 (
            .O(N__41104),
            .I(N__41101));
    LocalMux I__8276 (
            .O(N__41101),
            .I(N__41097));
    InMux I__8275 (
            .O(N__41100),
            .I(N__41094));
    Odrv4 I__8274 (
            .O(N__41097),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_27));
    LocalMux I__8273 (
            .O(N__41094),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_27));
    InMux I__8272 (
            .O(N__41089),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ));
    InMux I__8271 (
            .O(N__41086),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ));
    InMux I__8270 (
            .O(N__41083),
            .I(N__41080));
    LocalMux I__8269 (
            .O(N__41080),
            .I(N__41076));
    InMux I__8268 (
            .O(N__41079),
            .I(N__41073));
    Span4Mux_h I__8267 (
            .O(N__41076),
            .I(N__41070));
    LocalMux I__8266 (
            .O(N__41073),
            .I(N__41067));
    Odrv4 I__8265 (
            .O(N__41070),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_13));
    Odrv4 I__8264 (
            .O(N__41067),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_13));
    InMux I__8263 (
            .O(N__41062),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ));
    InMux I__8262 (
            .O(N__41059),
            .I(N__41056));
    LocalMux I__8261 (
            .O(N__41056),
            .I(N__41052));
    InMux I__8260 (
            .O(N__41055),
            .I(N__41049));
    Span4Mux_h I__8259 (
            .O(N__41052),
            .I(N__41046));
    LocalMux I__8258 (
            .O(N__41049),
            .I(N__41043));
    Odrv4 I__8257 (
            .O(N__41046),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_14));
    Odrv4 I__8256 (
            .O(N__41043),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_14));
    InMux I__8255 (
            .O(N__41038),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ));
    InMux I__8254 (
            .O(N__41035),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ));
    InMux I__8253 (
            .O(N__41032),
            .I(N__41028));
    InMux I__8252 (
            .O(N__41031),
            .I(N__41025));
    LocalMux I__8251 (
            .O(N__41028),
            .I(N__41022));
    LocalMux I__8250 (
            .O(N__41025),
            .I(N__41019));
    Span4Mux_h I__8249 (
            .O(N__41022),
            .I(N__41016));
    Span4Mux_h I__8248 (
            .O(N__41019),
            .I(N__41013));
    Odrv4 I__8247 (
            .O(N__41016),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_16));
    Odrv4 I__8246 (
            .O(N__41013),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_16));
    InMux I__8245 (
            .O(N__41008),
            .I(bfn_15_9_0_));
    InMux I__8244 (
            .O(N__41005),
            .I(N__41001));
    InMux I__8243 (
            .O(N__41004),
            .I(N__40998));
    LocalMux I__8242 (
            .O(N__41001),
            .I(N__40995));
    LocalMux I__8241 (
            .O(N__40998),
            .I(N__40992));
    Span4Mux_h I__8240 (
            .O(N__40995),
            .I(N__40989));
    Span4Mux_h I__8239 (
            .O(N__40992),
            .I(N__40986));
    Odrv4 I__8238 (
            .O(N__40989),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_17));
    Odrv4 I__8237 (
            .O(N__40986),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_17));
    InMux I__8236 (
            .O(N__40981),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ));
    InMux I__8235 (
            .O(N__40978),
            .I(N__40974));
    InMux I__8234 (
            .O(N__40977),
            .I(N__40971));
    LocalMux I__8233 (
            .O(N__40974),
            .I(N__40966));
    LocalMux I__8232 (
            .O(N__40971),
            .I(N__40966));
    Span4Mux_h I__8231 (
            .O(N__40966),
            .I(N__40963));
    Odrv4 I__8230 (
            .O(N__40963),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_18));
    InMux I__8229 (
            .O(N__40960),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ));
    InMux I__8228 (
            .O(N__40957),
            .I(N__40953));
    InMux I__8227 (
            .O(N__40956),
            .I(N__40950));
    LocalMux I__8226 (
            .O(N__40953),
            .I(N__40947));
    LocalMux I__8225 (
            .O(N__40950),
            .I(N__40944));
    Span4Mux_h I__8224 (
            .O(N__40947),
            .I(N__40941));
    Span4Mux_v I__8223 (
            .O(N__40944),
            .I(N__40938));
    Odrv4 I__8222 (
            .O(N__40941),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_19));
    Odrv4 I__8221 (
            .O(N__40938),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_19));
    InMux I__8220 (
            .O(N__40933),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ));
    InMux I__8219 (
            .O(N__40930),
            .I(N__40927));
    LocalMux I__8218 (
            .O(N__40927),
            .I(N__40924));
    Span4Mux_v I__8217 (
            .O(N__40924),
            .I(N__40920));
    InMux I__8216 (
            .O(N__40923),
            .I(N__40917));
    Odrv4 I__8215 (
            .O(N__40920),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_20));
    LocalMux I__8214 (
            .O(N__40917),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_20));
    InMux I__8213 (
            .O(N__40912),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ));
    InMux I__8212 (
            .O(N__40909),
            .I(N__40906));
    LocalMux I__8211 (
            .O(N__40906),
            .I(N__40902));
    InMux I__8210 (
            .O(N__40905),
            .I(N__40899));
    Span4Mux_h I__8209 (
            .O(N__40902),
            .I(N__40896));
    LocalMux I__8208 (
            .O(N__40899),
            .I(N__40893));
    Odrv4 I__8207 (
            .O(N__40896),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_4));
    Odrv4 I__8206 (
            .O(N__40893),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_4));
    InMux I__8205 (
            .O(N__40888),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ));
    InMux I__8204 (
            .O(N__40885),
            .I(N__40882));
    LocalMux I__8203 (
            .O(N__40882),
            .I(N__40878));
    InMux I__8202 (
            .O(N__40881),
            .I(N__40875));
    Span4Mux_h I__8201 (
            .O(N__40878),
            .I(N__40872));
    LocalMux I__8200 (
            .O(N__40875),
            .I(N__40869));
    Odrv4 I__8199 (
            .O(N__40872),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_5));
    Odrv4 I__8198 (
            .O(N__40869),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_5));
    InMux I__8197 (
            .O(N__40864),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ));
    InMux I__8196 (
            .O(N__40861),
            .I(N__40858));
    LocalMux I__8195 (
            .O(N__40858),
            .I(N__40854));
    InMux I__8194 (
            .O(N__40857),
            .I(N__40851));
    Span4Mux_h I__8193 (
            .O(N__40854),
            .I(N__40848));
    LocalMux I__8192 (
            .O(N__40851),
            .I(N__40845));
    Odrv4 I__8191 (
            .O(N__40848),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_6));
    Odrv4 I__8190 (
            .O(N__40845),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_6));
    InMux I__8189 (
            .O(N__40840),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ));
    InMux I__8188 (
            .O(N__40837),
            .I(N__40834));
    LocalMux I__8187 (
            .O(N__40834),
            .I(N__40830));
    InMux I__8186 (
            .O(N__40833),
            .I(N__40827));
    Span4Mux_h I__8185 (
            .O(N__40830),
            .I(N__40824));
    LocalMux I__8184 (
            .O(N__40827),
            .I(N__40821));
    Odrv4 I__8183 (
            .O(N__40824),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_7));
    Odrv4 I__8182 (
            .O(N__40821),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_7));
    InMux I__8181 (
            .O(N__40816),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ));
    InMux I__8180 (
            .O(N__40813),
            .I(N__40809));
    InMux I__8179 (
            .O(N__40812),
            .I(N__40806));
    LocalMux I__8178 (
            .O(N__40809),
            .I(N__40803));
    LocalMux I__8177 (
            .O(N__40806),
            .I(N__40798));
    Span4Mux_h I__8176 (
            .O(N__40803),
            .I(N__40798));
    Odrv4 I__8175 (
            .O(N__40798),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_8));
    InMux I__8174 (
            .O(N__40795),
            .I(bfn_15_8_0_));
    InMux I__8173 (
            .O(N__40792),
            .I(N__40789));
    LocalMux I__8172 (
            .O(N__40789),
            .I(N__40785));
    InMux I__8171 (
            .O(N__40788),
            .I(N__40782));
    Span4Mux_h I__8170 (
            .O(N__40785),
            .I(N__40779));
    LocalMux I__8169 (
            .O(N__40782),
            .I(N__40776));
    Odrv4 I__8168 (
            .O(N__40779),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_9));
    Odrv4 I__8167 (
            .O(N__40776),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_9));
    InMux I__8166 (
            .O(N__40771),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ));
    InMux I__8165 (
            .O(N__40768),
            .I(N__40765));
    LocalMux I__8164 (
            .O(N__40765),
            .I(N__40761));
    InMux I__8163 (
            .O(N__40764),
            .I(N__40758));
    Span4Mux_v I__8162 (
            .O(N__40761),
            .I(N__40755));
    LocalMux I__8161 (
            .O(N__40758),
            .I(N__40752));
    Odrv4 I__8160 (
            .O(N__40755),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_10));
    Odrv4 I__8159 (
            .O(N__40752),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_10));
    InMux I__8158 (
            .O(N__40747),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ));
    InMux I__8157 (
            .O(N__40744),
            .I(N__40741));
    LocalMux I__8156 (
            .O(N__40741),
            .I(N__40737));
    InMux I__8155 (
            .O(N__40740),
            .I(N__40734));
    Span4Mux_v I__8154 (
            .O(N__40737),
            .I(N__40731));
    LocalMux I__8153 (
            .O(N__40734),
            .I(N__40728));
    Odrv4 I__8152 (
            .O(N__40731),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_11));
    Odrv4 I__8151 (
            .O(N__40728),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_11));
    InMux I__8150 (
            .O(N__40723),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ));
    InMux I__8149 (
            .O(N__40720),
            .I(N__40717));
    LocalMux I__8148 (
            .O(N__40717),
            .I(N__40713));
    InMux I__8147 (
            .O(N__40716),
            .I(N__40710));
    Span4Mux_h I__8146 (
            .O(N__40713),
            .I(N__40707));
    LocalMux I__8145 (
            .O(N__40710),
            .I(N__40704));
    Odrv4 I__8144 (
            .O(N__40707),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_12));
    Odrv4 I__8143 (
            .O(N__40704),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_12));
    InMux I__8142 (
            .O(N__40699),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ));
    InMux I__8141 (
            .O(N__40696),
            .I(N__40693));
    LocalMux I__8140 (
            .O(N__40693),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ));
    CascadeMux I__8139 (
            .O(N__40690),
            .I(N__40687));
    InMux I__8138 (
            .O(N__40687),
            .I(N__40684));
    LocalMux I__8137 (
            .O(N__40684),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ));
    InMux I__8136 (
            .O(N__40681),
            .I(N__40678));
    LocalMux I__8135 (
            .O(N__40678),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ));
    InMux I__8134 (
            .O(N__40675),
            .I(N__40672));
    LocalMux I__8133 (
            .O(N__40672),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ));
    InMux I__8132 (
            .O(N__40669),
            .I(N__40666));
    LocalMux I__8131 (
            .O(N__40666),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ));
    InMux I__8130 (
            .O(N__40663),
            .I(N__40660));
    LocalMux I__8129 (
            .O(N__40660),
            .I(\phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ));
    InMux I__8128 (
            .O(N__40657),
            .I(N__40654));
    LocalMux I__8127 (
            .O(N__40654),
            .I(N__40650));
    InMux I__8126 (
            .O(N__40653),
            .I(N__40647));
    Span4Mux_v I__8125 (
            .O(N__40650),
            .I(N__40644));
    LocalMux I__8124 (
            .O(N__40647),
            .I(N__40641));
    Odrv4 I__8123 (
            .O(N__40644),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_1));
    Odrv4 I__8122 (
            .O(N__40641),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_1));
    InMux I__8121 (
            .O(N__40636),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ));
    InMux I__8120 (
            .O(N__40633),
            .I(N__40630));
    LocalMux I__8119 (
            .O(N__40630),
            .I(N__40626));
    InMux I__8118 (
            .O(N__40629),
            .I(N__40623));
    Span4Mux_v I__8117 (
            .O(N__40626),
            .I(N__40620));
    LocalMux I__8116 (
            .O(N__40623),
            .I(N__40617));
    Odrv4 I__8115 (
            .O(N__40620),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_2));
    Odrv4 I__8114 (
            .O(N__40617),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_2));
    InMux I__8113 (
            .O(N__40612),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ));
    InMux I__8112 (
            .O(N__40609),
            .I(N__40606));
    LocalMux I__8111 (
            .O(N__40606),
            .I(N__40602));
    InMux I__8110 (
            .O(N__40605),
            .I(N__40599));
    Span4Mux_v I__8109 (
            .O(N__40602),
            .I(N__40596));
    LocalMux I__8108 (
            .O(N__40599),
            .I(N__40593));
    Odrv4 I__8107 (
            .O(N__40596),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_3));
    Odrv4 I__8106 (
            .O(N__40593),
            .I(phase_controller_inst1_stoper_hc_target_ticks_1_i_3));
    InMux I__8105 (
            .O(N__40588),
            .I(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ));
    CascadeMux I__8104 (
            .O(N__40585),
            .I(N__40582));
    InMux I__8103 (
            .O(N__40582),
            .I(N__40579));
    LocalMux I__8102 (
            .O(N__40579),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ));
    InMux I__8101 (
            .O(N__40576),
            .I(N__40573));
    LocalMux I__8100 (
            .O(N__40573),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ));
    InMux I__8099 (
            .O(N__40570),
            .I(N__40567));
    LocalMux I__8098 (
            .O(N__40567),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ));
    CascadeMux I__8097 (
            .O(N__40564),
            .I(N__40561));
    InMux I__8096 (
            .O(N__40561),
            .I(N__40558));
    LocalMux I__8095 (
            .O(N__40558),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ));
    InMux I__8094 (
            .O(N__40555),
            .I(N__40552));
    LocalMux I__8093 (
            .O(N__40552),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ));
    InMux I__8092 (
            .O(N__40549),
            .I(N__40546));
    LocalMux I__8091 (
            .O(N__40546),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ));
    InMux I__8090 (
            .O(N__40543),
            .I(N__40540));
    LocalMux I__8089 (
            .O(N__40540),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ));
    InMux I__8088 (
            .O(N__40537),
            .I(N__40534));
    LocalMux I__8087 (
            .O(N__40534),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ));
    InMux I__8086 (
            .O(N__40531),
            .I(N__40528));
    LocalMux I__8085 (
            .O(N__40528),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ));
    CascadeMux I__8084 (
            .O(N__40525),
            .I(\current_shift_inst.control_input_31_cascade_ ));
    CascadeMux I__8083 (
            .O(N__40522),
            .I(N__40519));
    InMux I__8082 (
            .O(N__40519),
            .I(N__40516));
    LocalMux I__8081 (
            .O(N__40516),
            .I(N__40513));
    Odrv4 I__8080 (
            .O(N__40513),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ));
    CascadeMux I__8079 (
            .O(N__40510),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ));
    InMux I__8078 (
            .O(N__40507),
            .I(N__40504));
    LocalMux I__8077 (
            .O(N__40504),
            .I(N__40500));
    InMux I__8076 (
            .O(N__40503),
            .I(N__40497));
    Span4Mux_h I__8075 (
            .O(N__40500),
            .I(N__40494));
    LocalMux I__8074 (
            .O(N__40497),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    Odrv4 I__8073 (
            .O(N__40494),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ));
    CascadeMux I__8072 (
            .O(N__40489),
            .I(N__40486));
    InMux I__8071 (
            .O(N__40486),
            .I(N__40483));
    LocalMux I__8070 (
            .O(N__40483),
            .I(N__40479));
    InMux I__8069 (
            .O(N__40482),
            .I(N__40476));
    Span4Mux_h I__8068 (
            .O(N__40479),
            .I(N__40473));
    LocalMux I__8067 (
            .O(N__40476),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    Odrv4 I__8066 (
            .O(N__40473),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ));
    CascadeMux I__8065 (
            .O(N__40468),
            .I(N__40464));
    InMux I__8064 (
            .O(N__40467),
            .I(N__40461));
    InMux I__8063 (
            .O(N__40464),
            .I(N__40458));
    LocalMux I__8062 (
            .O(N__40461),
            .I(N__40455));
    LocalMux I__8061 (
            .O(N__40458),
            .I(N__40450));
    Span4Mux_v I__8060 (
            .O(N__40455),
            .I(N__40450));
    Odrv4 I__8059 (
            .O(N__40450),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ));
    CascadeMux I__8058 (
            .O(N__40447),
            .I(N__40444));
    InMux I__8057 (
            .O(N__40444),
            .I(N__40441));
    LocalMux I__8056 (
            .O(N__40441),
            .I(N__40437));
    InMux I__8055 (
            .O(N__40440),
            .I(N__40434));
    Span4Mux_h I__8054 (
            .O(N__40437),
            .I(N__40431));
    LocalMux I__8053 (
            .O(N__40434),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    Odrv4 I__8052 (
            .O(N__40431),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ));
    InMux I__8051 (
            .O(N__40426),
            .I(N__40423));
    LocalMux I__8050 (
            .O(N__40423),
            .I(N__40419));
    InMux I__8049 (
            .O(N__40422),
            .I(N__40416));
    Span4Mux_v I__8048 (
            .O(N__40419),
            .I(N__40411));
    LocalMux I__8047 (
            .O(N__40416),
            .I(N__40411));
    Odrv4 I__8046 (
            .O(N__40411),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ));
    InMux I__8045 (
            .O(N__40408),
            .I(N__40402));
    InMux I__8044 (
            .O(N__40407),
            .I(N__40402));
    LocalMux I__8043 (
            .O(N__40402),
            .I(N__40399));
    Odrv4 I__8042 (
            .O(N__40399),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ));
    CascadeMux I__8041 (
            .O(N__40396),
            .I(N__40393));
    InMux I__8040 (
            .O(N__40393),
            .I(N__40387));
    InMux I__8039 (
            .O(N__40392),
            .I(N__40387));
    LocalMux I__8038 (
            .O(N__40387),
            .I(N__40384));
    Span4Mux_h I__8037 (
            .O(N__40384),
            .I(N__40381));
    Odrv4 I__8036 (
            .O(N__40381),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ));
    InMux I__8035 (
            .O(N__40378),
            .I(N__40372));
    InMux I__8034 (
            .O(N__40377),
            .I(N__40372));
    LocalMux I__8033 (
            .O(N__40372),
            .I(N__40369));
    Odrv12 I__8032 (
            .O(N__40369),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ));
    ClkMux I__8031 (
            .O(N__40366),
            .I(N__40363));
    GlobalMux I__8030 (
            .O(N__40363),
            .I(N__40360));
    gio2CtrlBuf I__8029 (
            .O(N__40360),
            .I(delay_hc_input_c_g));
    CascadeMux I__8028 (
            .O(N__40357),
            .I(N__40354));
    InMux I__8027 (
            .O(N__40354),
            .I(N__40351));
    LocalMux I__8026 (
            .O(N__40351),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ));
    InMux I__8025 (
            .O(N__40348),
            .I(N__40345));
    LocalMux I__8024 (
            .O(N__40345),
            .I(N__40342));
    Odrv4 I__8023 (
            .O(N__40342),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ));
    InMux I__8022 (
            .O(N__40339),
            .I(\current_shift_inst.control_input_cry_22 ));
    InMux I__8021 (
            .O(N__40336),
            .I(N__40333));
    LocalMux I__8020 (
            .O(N__40333),
            .I(N__40330));
    Odrv4 I__8019 (
            .O(N__40330),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ));
    InMux I__8018 (
            .O(N__40327),
            .I(bfn_14_22_0_));
    InMux I__8017 (
            .O(N__40324),
            .I(N__40321));
    LocalMux I__8016 (
            .O(N__40321),
            .I(N__40318));
    Odrv4 I__8015 (
            .O(N__40318),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ));
    InMux I__8014 (
            .O(N__40315),
            .I(\current_shift_inst.control_input_cry_24 ));
    InMux I__8013 (
            .O(N__40312),
            .I(N__40309));
    LocalMux I__8012 (
            .O(N__40309),
            .I(N__40306));
    Odrv4 I__8011 (
            .O(N__40306),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ));
    InMux I__8010 (
            .O(N__40303),
            .I(\current_shift_inst.control_input_cry_25 ));
    InMux I__8009 (
            .O(N__40300),
            .I(N__40297));
    LocalMux I__8008 (
            .O(N__40297),
            .I(N__40294));
    Odrv4 I__8007 (
            .O(N__40294),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ));
    InMux I__8006 (
            .O(N__40291),
            .I(\current_shift_inst.control_input_cry_26 ));
    InMux I__8005 (
            .O(N__40288),
            .I(N__40285));
    LocalMux I__8004 (
            .O(N__40285),
            .I(N__40282));
    Odrv4 I__8003 (
            .O(N__40282),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ));
    InMux I__8002 (
            .O(N__40279),
            .I(\current_shift_inst.control_input_cry_27 ));
    InMux I__8001 (
            .O(N__40276),
            .I(N__40273));
    LocalMux I__8000 (
            .O(N__40273),
            .I(N__40270));
    Odrv4 I__7999 (
            .O(N__40270),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ));
    InMux I__7998 (
            .O(N__40267),
            .I(\current_shift_inst.control_input_cry_28 ));
    InMux I__7997 (
            .O(N__40264),
            .I(\current_shift_inst.control_input_cry_29 ));
    InMux I__7996 (
            .O(N__40261),
            .I(N__40258));
    LocalMux I__7995 (
            .O(N__40258),
            .I(N__40255));
    Odrv4 I__7994 (
            .O(N__40255),
            .I(\current_shift_inst.control_input_31 ));
    InMux I__7993 (
            .O(N__40252),
            .I(N__40249));
    LocalMux I__7992 (
            .O(N__40249),
            .I(N__40246));
    Odrv4 I__7991 (
            .O(N__40246),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ));
    InMux I__7990 (
            .O(N__40243),
            .I(\current_shift_inst.control_input_cry_14 ));
    InMux I__7989 (
            .O(N__40240),
            .I(N__40237));
    LocalMux I__7988 (
            .O(N__40237),
            .I(N__40234));
    Odrv4 I__7987 (
            .O(N__40234),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ));
    InMux I__7986 (
            .O(N__40231),
            .I(bfn_14_21_0_));
    InMux I__7985 (
            .O(N__40228),
            .I(N__40225));
    LocalMux I__7984 (
            .O(N__40225),
            .I(N__40222));
    Odrv4 I__7983 (
            .O(N__40222),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ));
    InMux I__7982 (
            .O(N__40219),
            .I(\current_shift_inst.control_input_cry_16 ));
    InMux I__7981 (
            .O(N__40216),
            .I(N__40213));
    LocalMux I__7980 (
            .O(N__40213),
            .I(N__40210));
    Odrv4 I__7979 (
            .O(N__40210),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ));
    InMux I__7978 (
            .O(N__40207),
            .I(\current_shift_inst.control_input_cry_17 ));
    InMux I__7977 (
            .O(N__40204),
            .I(N__40201));
    LocalMux I__7976 (
            .O(N__40201),
            .I(N__40198));
    Odrv4 I__7975 (
            .O(N__40198),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ));
    InMux I__7974 (
            .O(N__40195),
            .I(\current_shift_inst.control_input_cry_18 ));
    InMux I__7973 (
            .O(N__40192),
            .I(N__40189));
    LocalMux I__7972 (
            .O(N__40189),
            .I(N__40186));
    Odrv4 I__7971 (
            .O(N__40186),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ));
    InMux I__7970 (
            .O(N__40183),
            .I(\current_shift_inst.control_input_cry_19 ));
    InMux I__7969 (
            .O(N__40180),
            .I(N__40177));
    LocalMux I__7968 (
            .O(N__40177),
            .I(N__40174));
    Odrv4 I__7967 (
            .O(N__40174),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ));
    InMux I__7966 (
            .O(N__40171),
            .I(\current_shift_inst.control_input_cry_20 ));
    CascadeMux I__7965 (
            .O(N__40168),
            .I(N__40165));
    InMux I__7964 (
            .O(N__40165),
            .I(N__40162));
    LocalMux I__7963 (
            .O(N__40162),
            .I(N__40159));
    Odrv4 I__7962 (
            .O(N__40159),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ));
    InMux I__7961 (
            .O(N__40156),
            .I(\current_shift_inst.control_input_cry_21 ));
    CascadeMux I__7960 (
            .O(N__40153),
            .I(N__40150));
    InMux I__7959 (
            .O(N__40150),
            .I(N__40147));
    LocalMux I__7958 (
            .O(N__40147),
            .I(N__40144));
    Odrv4 I__7957 (
            .O(N__40144),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ));
    InMux I__7956 (
            .O(N__40141),
            .I(\current_shift_inst.control_input_cry_5 ));
    InMux I__7955 (
            .O(N__40138),
            .I(N__40135));
    LocalMux I__7954 (
            .O(N__40135),
            .I(N__40132));
    Odrv4 I__7953 (
            .O(N__40132),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ));
    InMux I__7952 (
            .O(N__40129),
            .I(\current_shift_inst.control_input_cry_6 ));
    InMux I__7951 (
            .O(N__40126),
            .I(N__40123));
    LocalMux I__7950 (
            .O(N__40123),
            .I(N__40120));
    Odrv4 I__7949 (
            .O(N__40120),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ));
    InMux I__7948 (
            .O(N__40117),
            .I(bfn_14_20_0_));
    InMux I__7947 (
            .O(N__40114),
            .I(N__40111));
    LocalMux I__7946 (
            .O(N__40111),
            .I(N__40108));
    Odrv4 I__7945 (
            .O(N__40108),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ));
    InMux I__7944 (
            .O(N__40105),
            .I(\current_shift_inst.control_input_cry_8 ));
    InMux I__7943 (
            .O(N__40102),
            .I(N__40099));
    LocalMux I__7942 (
            .O(N__40099),
            .I(N__40096));
    Odrv4 I__7941 (
            .O(N__40096),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ));
    InMux I__7940 (
            .O(N__40093),
            .I(\current_shift_inst.control_input_cry_9 ));
    InMux I__7939 (
            .O(N__40090),
            .I(N__40087));
    LocalMux I__7938 (
            .O(N__40087),
            .I(N__40084));
    Odrv4 I__7937 (
            .O(N__40084),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ));
    InMux I__7936 (
            .O(N__40081),
            .I(\current_shift_inst.control_input_cry_10 ));
    InMux I__7935 (
            .O(N__40078),
            .I(N__40075));
    LocalMux I__7934 (
            .O(N__40075),
            .I(N__40072));
    Odrv4 I__7933 (
            .O(N__40072),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ));
    InMux I__7932 (
            .O(N__40069),
            .I(\current_shift_inst.control_input_cry_11 ));
    InMux I__7931 (
            .O(N__40066),
            .I(N__40063));
    LocalMux I__7930 (
            .O(N__40063),
            .I(N__40060));
    Odrv4 I__7929 (
            .O(N__40060),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ));
    InMux I__7928 (
            .O(N__40057),
            .I(\current_shift_inst.control_input_cry_12 ));
    CascadeMux I__7927 (
            .O(N__40054),
            .I(N__40051));
    InMux I__7926 (
            .O(N__40051),
            .I(N__40048));
    LocalMux I__7925 (
            .O(N__40048),
            .I(N__40045));
    Odrv4 I__7924 (
            .O(N__40045),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ));
    InMux I__7923 (
            .O(N__40042),
            .I(\current_shift_inst.control_input_cry_13 ));
    InMux I__7922 (
            .O(N__40039),
            .I(N__40036));
    LocalMux I__7921 (
            .O(N__40036),
            .I(N__40033));
    Odrv4 I__7920 (
            .O(N__40033),
            .I(\current_shift_inst.elapsed_time_ns_s1_fast_31 ));
    InMux I__7919 (
            .O(N__40030),
            .I(N__40027));
    LocalMux I__7918 (
            .O(N__40027),
            .I(N__40024));
    Odrv4 I__7917 (
            .O(N__40024),
            .I(\current_shift_inst.control_input_1 ));
    InMux I__7916 (
            .O(N__40021),
            .I(N__40018));
    LocalMux I__7915 (
            .O(N__40018),
            .I(N__40015));
    Odrv4 I__7914 (
            .O(N__40015),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ));
    InMux I__7913 (
            .O(N__40012),
            .I(\current_shift_inst.control_input_cry_0 ));
    InMux I__7912 (
            .O(N__40009),
            .I(N__40006));
    LocalMux I__7911 (
            .O(N__40006),
            .I(N__40003));
    Odrv4 I__7910 (
            .O(N__40003),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ));
    InMux I__7909 (
            .O(N__40000),
            .I(\current_shift_inst.control_input_cry_1 ));
    InMux I__7908 (
            .O(N__39997),
            .I(N__39994));
    LocalMux I__7907 (
            .O(N__39994),
            .I(N__39991));
    Odrv4 I__7906 (
            .O(N__39991),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ));
    InMux I__7905 (
            .O(N__39988),
            .I(\current_shift_inst.control_input_cry_2 ));
    InMux I__7904 (
            .O(N__39985),
            .I(N__39982));
    LocalMux I__7903 (
            .O(N__39982),
            .I(N__39979));
    Span4Mux_h I__7902 (
            .O(N__39979),
            .I(N__39976));
    Odrv4 I__7901 (
            .O(N__39976),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ));
    InMux I__7900 (
            .O(N__39973),
            .I(\current_shift_inst.control_input_cry_3 ));
    InMux I__7899 (
            .O(N__39970),
            .I(N__39967));
    LocalMux I__7898 (
            .O(N__39967),
            .I(N__39964));
    Odrv4 I__7897 (
            .O(N__39964),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ));
    InMux I__7896 (
            .O(N__39961),
            .I(\current_shift_inst.control_input_cry_4 ));
    CascadeMux I__7895 (
            .O(N__39958),
            .I(N__39954));
    CascadeMux I__7894 (
            .O(N__39957),
            .I(N__39951));
    InMux I__7893 (
            .O(N__39954),
            .I(N__39945));
    InMux I__7892 (
            .O(N__39951),
            .I(N__39945));
    InMux I__7891 (
            .O(N__39950),
            .I(N__39942));
    LocalMux I__7890 (
            .O(N__39945),
            .I(N__39939));
    LocalMux I__7889 (
            .O(N__39942),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    Odrv12 I__7888 (
            .O(N__39939),
            .I(\current_shift_inst.timer_s1.counterZ0Z_21 ));
    InMux I__7887 (
            .O(N__39934),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ));
    InMux I__7886 (
            .O(N__39931),
            .I(N__39925));
    InMux I__7885 (
            .O(N__39930),
            .I(N__39925));
    LocalMux I__7884 (
            .O(N__39925),
            .I(N__39921));
    InMux I__7883 (
            .O(N__39924),
            .I(N__39918));
    Span4Mux_v I__7882 (
            .O(N__39921),
            .I(N__39915));
    LocalMux I__7881 (
            .O(N__39918),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    Odrv4 I__7880 (
            .O(N__39915),
            .I(\current_shift_inst.timer_s1.counterZ0Z_22 ));
    InMux I__7879 (
            .O(N__39910),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__7878 (
            .O(N__39907),
            .I(N__39904));
    InMux I__7877 (
            .O(N__39904),
            .I(N__39900));
    InMux I__7876 (
            .O(N__39903),
            .I(N__39897));
    LocalMux I__7875 (
            .O(N__39900),
            .I(N__39891));
    LocalMux I__7874 (
            .O(N__39897),
            .I(N__39891));
    InMux I__7873 (
            .O(N__39896),
            .I(N__39888));
    Span4Mux_v I__7872 (
            .O(N__39891),
            .I(N__39885));
    LocalMux I__7871 (
            .O(N__39888),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    Odrv4 I__7870 (
            .O(N__39885),
            .I(\current_shift_inst.timer_s1.counterZ0Z_23 ));
    InMux I__7869 (
            .O(N__39880),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__7868 (
            .O(N__39877),
            .I(N__39873));
    CascadeMux I__7867 (
            .O(N__39876),
            .I(N__39870));
    InMux I__7866 (
            .O(N__39873),
            .I(N__39866));
    InMux I__7865 (
            .O(N__39870),
            .I(N__39863));
    InMux I__7864 (
            .O(N__39869),
            .I(N__39860));
    LocalMux I__7863 (
            .O(N__39866),
            .I(N__39855));
    LocalMux I__7862 (
            .O(N__39863),
            .I(N__39855));
    LocalMux I__7861 (
            .O(N__39860),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    Odrv12 I__7860 (
            .O(N__39855),
            .I(\current_shift_inst.timer_s1.counterZ0Z_24 ));
    InMux I__7859 (
            .O(N__39850),
            .I(bfn_14_18_0_));
    CascadeMux I__7858 (
            .O(N__39847),
            .I(N__39844));
    InMux I__7857 (
            .O(N__39844),
            .I(N__39841));
    LocalMux I__7856 (
            .O(N__39841),
            .I(N__39836));
    InMux I__7855 (
            .O(N__39840),
            .I(N__39833));
    InMux I__7854 (
            .O(N__39839),
            .I(N__39830));
    Sp12to4 I__7853 (
            .O(N__39836),
            .I(N__39825));
    LocalMux I__7852 (
            .O(N__39833),
            .I(N__39825));
    LocalMux I__7851 (
            .O(N__39830),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    Odrv12 I__7850 (
            .O(N__39825),
            .I(\current_shift_inst.timer_s1.counterZ0Z_25 ));
    InMux I__7849 (
            .O(N__39820),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ));
    InMux I__7848 (
            .O(N__39817),
            .I(N__39813));
    InMux I__7847 (
            .O(N__39816),
            .I(N__39810));
    LocalMux I__7846 (
            .O(N__39813),
            .I(N__39807));
    LocalMux I__7845 (
            .O(N__39810),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    Odrv12 I__7844 (
            .O(N__39807),
            .I(\current_shift_inst.timer_s1.counterZ0Z_28 ));
    CascadeMux I__7843 (
            .O(N__39802),
            .I(N__39799));
    InMux I__7842 (
            .O(N__39799),
            .I(N__39794));
    InMux I__7841 (
            .O(N__39798),
            .I(N__39791));
    InMux I__7840 (
            .O(N__39797),
            .I(N__39788));
    LocalMux I__7839 (
            .O(N__39794),
            .I(N__39783));
    LocalMux I__7838 (
            .O(N__39791),
            .I(N__39783));
    LocalMux I__7837 (
            .O(N__39788),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    Odrv12 I__7836 (
            .O(N__39783),
            .I(\current_shift_inst.timer_s1.counterZ0Z_26 ));
    InMux I__7835 (
            .O(N__39778),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ));
    InMux I__7834 (
            .O(N__39775),
            .I(N__39772));
    LocalMux I__7833 (
            .O(N__39772),
            .I(N__39768));
    InMux I__7832 (
            .O(N__39771),
            .I(N__39765));
    Span4Mux_v I__7831 (
            .O(N__39768),
            .I(N__39762));
    LocalMux I__7830 (
            .O(N__39765),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    Odrv4 I__7829 (
            .O(N__39762),
            .I(\current_shift_inst.timer_s1.counterZ0Z_29 ));
    CascadeMux I__7828 (
            .O(N__39757),
            .I(N__39754));
    InMux I__7827 (
            .O(N__39754),
            .I(N__39749));
    InMux I__7826 (
            .O(N__39753),
            .I(N__39746));
    InMux I__7825 (
            .O(N__39752),
            .I(N__39743));
    LocalMux I__7824 (
            .O(N__39749),
            .I(N__39738));
    LocalMux I__7823 (
            .O(N__39746),
            .I(N__39738));
    LocalMux I__7822 (
            .O(N__39743),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    Odrv12 I__7821 (
            .O(N__39738),
            .I(\current_shift_inst.timer_s1.counterZ0Z_27 ));
    InMux I__7820 (
            .O(N__39733),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ));
    InMux I__7819 (
            .O(N__39730),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__7818 (
            .O(N__39727),
            .I(N__39723));
    CascadeMux I__7817 (
            .O(N__39726),
            .I(N__39720));
    InMux I__7816 (
            .O(N__39723),
            .I(N__39714));
    InMux I__7815 (
            .O(N__39720),
            .I(N__39714));
    InMux I__7814 (
            .O(N__39719),
            .I(N__39711));
    LocalMux I__7813 (
            .O(N__39714),
            .I(N__39708));
    LocalMux I__7812 (
            .O(N__39711),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    Odrv12 I__7811 (
            .O(N__39708),
            .I(\current_shift_inst.timer_s1.counterZ0Z_13 ));
    InMux I__7810 (
            .O(N__39703),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__7809 (
            .O(N__39700),
            .I(N__39696));
    CascadeMux I__7808 (
            .O(N__39699),
            .I(N__39693));
    InMux I__7807 (
            .O(N__39696),
            .I(N__39688));
    InMux I__7806 (
            .O(N__39693),
            .I(N__39688));
    LocalMux I__7805 (
            .O(N__39688),
            .I(N__39684));
    InMux I__7804 (
            .O(N__39687),
            .I(N__39681));
    Span4Mux_v I__7803 (
            .O(N__39684),
            .I(N__39678));
    LocalMux I__7802 (
            .O(N__39681),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    Odrv4 I__7801 (
            .O(N__39678),
            .I(\current_shift_inst.timer_s1.counterZ0Z_14 ));
    InMux I__7800 (
            .O(N__39673),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__7799 (
            .O(N__39670),
            .I(N__39667));
    InMux I__7798 (
            .O(N__39667),
            .I(N__39662));
    InMux I__7797 (
            .O(N__39666),
            .I(N__39659));
    InMux I__7796 (
            .O(N__39665),
            .I(N__39656));
    LocalMux I__7795 (
            .O(N__39662),
            .I(N__39651));
    LocalMux I__7794 (
            .O(N__39659),
            .I(N__39651));
    LocalMux I__7793 (
            .O(N__39656),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    Odrv12 I__7792 (
            .O(N__39651),
            .I(\current_shift_inst.timer_s1.counterZ0Z_15 ));
    InMux I__7791 (
            .O(N__39646),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__7790 (
            .O(N__39643),
            .I(N__39640));
    InMux I__7789 (
            .O(N__39640),
            .I(N__39637));
    LocalMux I__7788 (
            .O(N__39637),
            .I(N__39632));
    InMux I__7787 (
            .O(N__39636),
            .I(N__39629));
    InMux I__7786 (
            .O(N__39635),
            .I(N__39626));
    Sp12to4 I__7785 (
            .O(N__39632),
            .I(N__39621));
    LocalMux I__7784 (
            .O(N__39629),
            .I(N__39621));
    LocalMux I__7783 (
            .O(N__39626),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    Odrv12 I__7782 (
            .O(N__39621),
            .I(\current_shift_inst.timer_s1.counterZ0Z_16 ));
    InMux I__7781 (
            .O(N__39616),
            .I(bfn_14_17_0_));
    CascadeMux I__7780 (
            .O(N__39613),
            .I(N__39610));
    InMux I__7779 (
            .O(N__39610),
            .I(N__39607));
    LocalMux I__7778 (
            .O(N__39607),
            .I(N__39602));
    InMux I__7777 (
            .O(N__39606),
            .I(N__39599));
    InMux I__7776 (
            .O(N__39605),
            .I(N__39596));
    Sp12to4 I__7775 (
            .O(N__39602),
            .I(N__39591));
    LocalMux I__7774 (
            .O(N__39599),
            .I(N__39591));
    LocalMux I__7773 (
            .O(N__39596),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    Odrv12 I__7772 (
            .O(N__39591),
            .I(\current_shift_inst.timer_s1.counterZ0Z_17 ));
    InMux I__7771 (
            .O(N__39586),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ));
    InMux I__7770 (
            .O(N__39583),
            .I(N__39576));
    InMux I__7769 (
            .O(N__39582),
            .I(N__39576));
    InMux I__7768 (
            .O(N__39581),
            .I(N__39573));
    LocalMux I__7767 (
            .O(N__39576),
            .I(N__39570));
    LocalMux I__7766 (
            .O(N__39573),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    Odrv12 I__7765 (
            .O(N__39570),
            .I(\current_shift_inst.timer_s1.counterZ0Z_18 ));
    InMux I__7764 (
            .O(N__39565),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ));
    InMux I__7763 (
            .O(N__39562),
            .I(N__39555));
    InMux I__7762 (
            .O(N__39561),
            .I(N__39555));
    InMux I__7761 (
            .O(N__39560),
            .I(N__39552));
    LocalMux I__7760 (
            .O(N__39555),
            .I(N__39549));
    LocalMux I__7759 (
            .O(N__39552),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    Odrv12 I__7758 (
            .O(N__39549),
            .I(\current_shift_inst.timer_s1.counterZ0Z_19 ));
    InMux I__7757 (
            .O(N__39544),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ));
    CascadeMux I__7756 (
            .O(N__39541),
            .I(N__39537));
    CascadeMux I__7755 (
            .O(N__39540),
            .I(N__39534));
    InMux I__7754 (
            .O(N__39537),
            .I(N__39528));
    InMux I__7753 (
            .O(N__39534),
            .I(N__39528));
    InMux I__7752 (
            .O(N__39533),
            .I(N__39525));
    LocalMux I__7751 (
            .O(N__39528),
            .I(N__39522));
    LocalMux I__7750 (
            .O(N__39525),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    Odrv12 I__7749 (
            .O(N__39522),
            .I(\current_shift_inst.timer_s1.counterZ0Z_20 ));
    InMux I__7748 (
            .O(N__39517),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ));
    InMux I__7747 (
            .O(N__39514),
            .I(N__39508));
    InMux I__7746 (
            .O(N__39513),
            .I(N__39508));
    LocalMux I__7745 (
            .O(N__39508),
            .I(N__39504));
    InMux I__7744 (
            .O(N__39507),
            .I(N__39501));
    Span4Mux_v I__7743 (
            .O(N__39504),
            .I(N__39498));
    LocalMux I__7742 (
            .O(N__39501),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    Odrv4 I__7741 (
            .O(N__39498),
            .I(\current_shift_inst.timer_s1.counterZ0Z_4 ));
    InMux I__7740 (
            .O(N__39493),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__7739 (
            .O(N__39490),
            .I(N__39486));
    CascadeMux I__7738 (
            .O(N__39489),
            .I(N__39483));
    InMux I__7737 (
            .O(N__39486),
            .I(N__39477));
    InMux I__7736 (
            .O(N__39483),
            .I(N__39477));
    InMux I__7735 (
            .O(N__39482),
            .I(N__39474));
    LocalMux I__7734 (
            .O(N__39477),
            .I(N__39471));
    LocalMux I__7733 (
            .O(N__39474),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    Odrv12 I__7732 (
            .O(N__39471),
            .I(\current_shift_inst.timer_s1.counterZ0Z_5 ));
    InMux I__7731 (
            .O(N__39466),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__7730 (
            .O(N__39463),
            .I(N__39459));
    CascadeMux I__7729 (
            .O(N__39462),
            .I(N__39456));
    InMux I__7728 (
            .O(N__39459),
            .I(N__39451));
    InMux I__7727 (
            .O(N__39456),
            .I(N__39451));
    LocalMux I__7726 (
            .O(N__39451),
            .I(N__39447));
    InMux I__7725 (
            .O(N__39450),
            .I(N__39444));
    Span4Mux_v I__7724 (
            .O(N__39447),
            .I(N__39441));
    LocalMux I__7723 (
            .O(N__39444),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    Odrv4 I__7722 (
            .O(N__39441),
            .I(\current_shift_inst.timer_s1.counterZ0Z_6 ));
    InMux I__7721 (
            .O(N__39436),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__7720 (
            .O(N__39433),
            .I(N__39430));
    InMux I__7719 (
            .O(N__39430),
            .I(N__39426));
    InMux I__7718 (
            .O(N__39429),
            .I(N__39423));
    LocalMux I__7717 (
            .O(N__39426),
            .I(N__39417));
    LocalMux I__7716 (
            .O(N__39423),
            .I(N__39417));
    InMux I__7715 (
            .O(N__39422),
            .I(N__39414));
    Span4Mux_v I__7714 (
            .O(N__39417),
            .I(N__39411));
    LocalMux I__7713 (
            .O(N__39414),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    Odrv4 I__7712 (
            .O(N__39411),
            .I(\current_shift_inst.timer_s1.counterZ0Z_7 ));
    InMux I__7711 (
            .O(N__39406),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__7710 (
            .O(N__39403),
            .I(N__39400));
    InMux I__7709 (
            .O(N__39400),
            .I(N__39395));
    InMux I__7708 (
            .O(N__39399),
            .I(N__39392));
    InMux I__7707 (
            .O(N__39398),
            .I(N__39389));
    LocalMux I__7706 (
            .O(N__39395),
            .I(N__39384));
    LocalMux I__7705 (
            .O(N__39392),
            .I(N__39384));
    LocalMux I__7704 (
            .O(N__39389),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    Odrv12 I__7703 (
            .O(N__39384),
            .I(\current_shift_inst.timer_s1.counterZ0Z_8 ));
    InMux I__7702 (
            .O(N__39379),
            .I(bfn_14_16_0_));
    CascadeMux I__7701 (
            .O(N__39376),
            .I(N__39373));
    InMux I__7700 (
            .O(N__39373),
            .I(N__39370));
    LocalMux I__7699 (
            .O(N__39370),
            .I(N__39365));
    InMux I__7698 (
            .O(N__39369),
            .I(N__39362));
    InMux I__7697 (
            .O(N__39368),
            .I(N__39359));
    Sp12to4 I__7696 (
            .O(N__39365),
            .I(N__39354));
    LocalMux I__7695 (
            .O(N__39362),
            .I(N__39354));
    LocalMux I__7694 (
            .O(N__39359),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    Odrv12 I__7693 (
            .O(N__39354),
            .I(\current_shift_inst.timer_s1.counterZ0Z_9 ));
    InMux I__7692 (
            .O(N__39349),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__7691 (
            .O(N__39346),
            .I(N__39343));
    InMux I__7690 (
            .O(N__39343),
            .I(N__39339));
    InMux I__7689 (
            .O(N__39342),
            .I(N__39336));
    LocalMux I__7688 (
            .O(N__39339),
            .I(N__39330));
    LocalMux I__7687 (
            .O(N__39336),
            .I(N__39330));
    InMux I__7686 (
            .O(N__39335),
            .I(N__39327));
    Span4Mux_v I__7685 (
            .O(N__39330),
            .I(N__39324));
    LocalMux I__7684 (
            .O(N__39327),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    Odrv4 I__7683 (
            .O(N__39324),
            .I(\current_shift_inst.timer_s1.counterZ0Z_10 ));
    InMux I__7682 (
            .O(N__39319),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ));
    InMux I__7681 (
            .O(N__39316),
            .I(N__39310));
    InMux I__7680 (
            .O(N__39315),
            .I(N__39310));
    LocalMux I__7679 (
            .O(N__39310),
            .I(N__39306));
    InMux I__7678 (
            .O(N__39309),
            .I(N__39303));
    Span4Mux_v I__7677 (
            .O(N__39306),
            .I(N__39300));
    LocalMux I__7676 (
            .O(N__39303),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    Odrv4 I__7675 (
            .O(N__39300),
            .I(\current_shift_inst.timer_s1.counterZ0Z_11 ));
    InMux I__7674 (
            .O(N__39295),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ));
    InMux I__7673 (
            .O(N__39292),
            .I(N__39286));
    InMux I__7672 (
            .O(N__39291),
            .I(N__39286));
    LocalMux I__7671 (
            .O(N__39286),
            .I(N__39282));
    InMux I__7670 (
            .O(N__39285),
            .I(N__39279));
    Span4Mux_v I__7669 (
            .O(N__39282),
            .I(N__39276));
    LocalMux I__7668 (
            .O(N__39279),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    Odrv4 I__7667 (
            .O(N__39276),
            .I(\current_shift_inst.timer_s1.counterZ0Z_12 ));
    InMux I__7666 (
            .O(N__39271),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ));
    InMux I__7665 (
            .O(N__39268),
            .I(\current_shift_inst.timer_s1.counter_cry_24 ));
    InMux I__7664 (
            .O(N__39265),
            .I(\current_shift_inst.timer_s1.counter_cry_25 ));
    InMux I__7663 (
            .O(N__39262),
            .I(\current_shift_inst.timer_s1.counter_cry_26 ));
    InMux I__7662 (
            .O(N__39259),
            .I(\current_shift_inst.timer_s1.counter_cry_27 ));
    InMux I__7661 (
            .O(N__39256),
            .I(\current_shift_inst.timer_s1.counter_cry_28 ));
    InMux I__7660 (
            .O(N__39253),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ));
    CascadeMux I__7659 (
            .O(N__39250),
            .I(N__39246));
    CascadeMux I__7658 (
            .O(N__39249),
            .I(N__39243));
    InMux I__7657 (
            .O(N__39246),
            .I(N__39238));
    InMux I__7656 (
            .O(N__39243),
            .I(N__39238));
    LocalMux I__7655 (
            .O(N__39238),
            .I(N__39234));
    InMux I__7654 (
            .O(N__39237),
            .I(N__39231));
    Span4Mux_v I__7653 (
            .O(N__39234),
            .I(N__39228));
    LocalMux I__7652 (
            .O(N__39231),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    Odrv4 I__7651 (
            .O(N__39228),
            .I(\current_shift_inst.timer_s1.counterZ0Z_2 ));
    InMux I__7650 (
            .O(N__39223),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__7649 (
            .O(N__39220),
            .I(N__39216));
    InMux I__7648 (
            .O(N__39219),
            .I(N__39213));
    InMux I__7647 (
            .O(N__39216),
            .I(N__39210));
    LocalMux I__7646 (
            .O(N__39213),
            .I(N__39204));
    LocalMux I__7645 (
            .O(N__39210),
            .I(N__39204));
    InMux I__7644 (
            .O(N__39209),
            .I(N__39201));
    Span4Mux_v I__7643 (
            .O(N__39204),
            .I(N__39198));
    LocalMux I__7642 (
            .O(N__39201),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    Odrv4 I__7641 (
            .O(N__39198),
            .I(\current_shift_inst.timer_s1.counterZ0Z_3 ));
    InMux I__7640 (
            .O(N__39193),
            .I(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ));
    InMux I__7639 (
            .O(N__39190),
            .I(bfn_14_13_0_));
    InMux I__7638 (
            .O(N__39187),
            .I(\current_shift_inst.timer_s1.counter_cry_16 ));
    InMux I__7637 (
            .O(N__39184),
            .I(\current_shift_inst.timer_s1.counter_cry_17 ));
    InMux I__7636 (
            .O(N__39181),
            .I(\current_shift_inst.timer_s1.counter_cry_18 ));
    InMux I__7635 (
            .O(N__39178),
            .I(\current_shift_inst.timer_s1.counter_cry_19 ));
    InMux I__7634 (
            .O(N__39175),
            .I(\current_shift_inst.timer_s1.counter_cry_20 ));
    InMux I__7633 (
            .O(N__39172),
            .I(\current_shift_inst.timer_s1.counter_cry_21 ));
    InMux I__7632 (
            .O(N__39169),
            .I(\current_shift_inst.timer_s1.counter_cry_22 ));
    InMux I__7631 (
            .O(N__39166),
            .I(bfn_14_14_0_));
    InMux I__7630 (
            .O(N__39163),
            .I(\current_shift_inst.timer_s1.counter_cry_6 ));
    InMux I__7629 (
            .O(N__39160),
            .I(bfn_14_12_0_));
    InMux I__7628 (
            .O(N__39157),
            .I(\current_shift_inst.timer_s1.counter_cry_8 ));
    InMux I__7627 (
            .O(N__39154),
            .I(\current_shift_inst.timer_s1.counter_cry_9 ));
    InMux I__7626 (
            .O(N__39151),
            .I(\current_shift_inst.timer_s1.counter_cry_10 ));
    InMux I__7625 (
            .O(N__39148),
            .I(\current_shift_inst.timer_s1.counter_cry_11 ));
    InMux I__7624 (
            .O(N__39145),
            .I(\current_shift_inst.timer_s1.counter_cry_12 ));
    InMux I__7623 (
            .O(N__39142),
            .I(\current_shift_inst.timer_s1.counter_cry_13 ));
    InMux I__7622 (
            .O(N__39139),
            .I(\current_shift_inst.timer_s1.counter_cry_14 ));
    InMux I__7621 (
            .O(N__39136),
            .I(N__39131));
    InMux I__7620 (
            .O(N__39135),
            .I(N__39126));
    InMux I__7619 (
            .O(N__39134),
            .I(N__39126));
    LocalMux I__7618 (
            .O(N__39131),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ));
    LocalMux I__7617 (
            .O(N__39126),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ));
    InMux I__7616 (
            .O(N__39121),
            .I(N__39115));
    InMux I__7615 (
            .O(N__39120),
            .I(N__39115));
    LocalMux I__7614 (
            .O(N__39115),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ));
    InMux I__7613 (
            .O(N__39112),
            .I(N__39107));
    InMux I__7612 (
            .O(N__39111),
            .I(N__39102));
    InMux I__7611 (
            .O(N__39110),
            .I(N__39102));
    LocalMux I__7610 (
            .O(N__39107),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ));
    LocalMux I__7609 (
            .O(N__39102),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ));
    CascadeMux I__7608 (
            .O(N__39097),
            .I(N__39094));
    InMux I__7607 (
            .O(N__39094),
            .I(N__39091));
    LocalMux I__7606 (
            .O(N__39091),
            .I(N__39088));
    Odrv12 I__7605 (
            .O(N__39088),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ));
    CascadeMux I__7604 (
            .O(N__39085),
            .I(N__39081));
    CascadeMux I__7603 (
            .O(N__39084),
            .I(N__39078));
    InMux I__7602 (
            .O(N__39081),
            .I(N__39073));
    InMux I__7601 (
            .O(N__39078),
            .I(N__39073));
    LocalMux I__7600 (
            .O(N__39073),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ));
    InMux I__7599 (
            .O(N__39070),
            .I(bfn_14_11_0_));
    InMux I__7598 (
            .O(N__39067),
            .I(\current_shift_inst.timer_s1.counter_cry_0 ));
    InMux I__7597 (
            .O(N__39064),
            .I(\current_shift_inst.timer_s1.counter_cry_1 ));
    InMux I__7596 (
            .O(N__39061),
            .I(\current_shift_inst.timer_s1.counter_cry_2 ));
    InMux I__7595 (
            .O(N__39058),
            .I(\current_shift_inst.timer_s1.counter_cry_3 ));
    InMux I__7594 (
            .O(N__39055),
            .I(\current_shift_inst.timer_s1.counter_cry_4 ));
    InMux I__7593 (
            .O(N__39052),
            .I(\current_shift_inst.timer_s1.counter_cry_5 ));
    InMux I__7592 (
            .O(N__39049),
            .I(N__39044));
    InMux I__7591 (
            .O(N__39048),
            .I(N__39039));
    InMux I__7590 (
            .O(N__39047),
            .I(N__39039));
    LocalMux I__7589 (
            .O(N__39044),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ));
    LocalMux I__7588 (
            .O(N__39039),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ));
    InMux I__7587 (
            .O(N__39034),
            .I(N__39028));
    InMux I__7586 (
            .O(N__39033),
            .I(N__39028));
    LocalMux I__7585 (
            .O(N__39028),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ));
    CascadeMux I__7584 (
            .O(N__39025),
            .I(N__39020));
    CascadeMux I__7583 (
            .O(N__39024),
            .I(N__39017));
    InMux I__7582 (
            .O(N__39023),
            .I(N__39014));
    InMux I__7581 (
            .O(N__39020),
            .I(N__39009));
    InMux I__7580 (
            .O(N__39017),
            .I(N__39009));
    LocalMux I__7579 (
            .O(N__39014),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ));
    LocalMux I__7578 (
            .O(N__39009),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ));
    InMux I__7577 (
            .O(N__39004),
            .I(N__39001));
    LocalMux I__7576 (
            .O(N__39001),
            .I(N__38998));
    Odrv12 I__7575 (
            .O(N__38998),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ));
    InMux I__7574 (
            .O(N__38995),
            .I(N__38989));
    InMux I__7573 (
            .O(N__38994),
            .I(N__38989));
    LocalMux I__7572 (
            .O(N__38989),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ));
    InMux I__7571 (
            .O(N__38986),
            .I(N__38983));
    LocalMux I__7570 (
            .O(N__38983),
            .I(N__38980));
    Odrv4 I__7569 (
            .O(N__38980),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt24 ));
    InMux I__7568 (
            .O(N__38977),
            .I(N__38971));
    InMux I__7567 (
            .O(N__38976),
            .I(N__38971));
    LocalMux I__7566 (
            .O(N__38971),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ));
    InMux I__7565 (
            .O(N__38968),
            .I(N__38963));
    InMux I__7564 (
            .O(N__38967),
            .I(N__38958));
    InMux I__7563 (
            .O(N__38966),
            .I(N__38958));
    LocalMux I__7562 (
            .O(N__38963),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    LocalMux I__7561 (
            .O(N__38958),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ));
    CascadeMux I__7560 (
            .O(N__38953),
            .I(N__38948));
    CascadeMux I__7559 (
            .O(N__38952),
            .I(N__38945));
    InMux I__7558 (
            .O(N__38951),
            .I(N__38942));
    InMux I__7557 (
            .O(N__38948),
            .I(N__38937));
    InMux I__7556 (
            .O(N__38945),
            .I(N__38937));
    LocalMux I__7555 (
            .O(N__38942),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ));
    LocalMux I__7554 (
            .O(N__38937),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ));
    CascadeMux I__7553 (
            .O(N__38932),
            .I(N__38929));
    InMux I__7552 (
            .O(N__38929),
            .I(N__38926));
    LocalMux I__7551 (
            .O(N__38926),
            .I(N__38923));
    Odrv4 I__7550 (
            .O(N__38923),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ));
    InMux I__7549 (
            .O(N__38920),
            .I(N__38914));
    InMux I__7548 (
            .O(N__38919),
            .I(N__38914));
    LocalMux I__7547 (
            .O(N__38914),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ));
    InMux I__7546 (
            .O(N__38911),
            .I(N__38908));
    LocalMux I__7545 (
            .O(N__38908),
            .I(N__38905));
    Odrv4 I__7544 (
            .O(N__38905),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt26 ));
    InMux I__7543 (
            .O(N__38902),
            .I(N__38896));
    InMux I__7542 (
            .O(N__38901),
            .I(N__38896));
    LocalMux I__7541 (
            .O(N__38896),
            .I(N__38893));
    Span4Mux_v I__7540 (
            .O(N__38893),
            .I(N__38890));
    Odrv4 I__7539 (
            .O(N__38890),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ));
    CascadeMux I__7538 (
            .O(N__38887),
            .I(N__38883));
    InMux I__7537 (
            .O(N__38886),
            .I(N__38878));
    InMux I__7536 (
            .O(N__38883),
            .I(N__38878));
    LocalMux I__7535 (
            .O(N__38878),
            .I(N__38875));
    Odrv4 I__7534 (
            .O(N__38875),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ));
    CascadeMux I__7533 (
            .O(N__38872),
            .I(N__38867));
    InMux I__7532 (
            .O(N__38871),
            .I(N__38864));
    InMux I__7531 (
            .O(N__38870),
            .I(N__38859));
    InMux I__7530 (
            .O(N__38867),
            .I(N__38859));
    LocalMux I__7529 (
            .O(N__38864),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ));
    LocalMux I__7528 (
            .O(N__38859),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ));
    InMux I__7527 (
            .O(N__38854),
            .I(N__38849));
    InMux I__7526 (
            .O(N__38853),
            .I(N__38844));
    InMux I__7525 (
            .O(N__38852),
            .I(N__38844));
    LocalMux I__7524 (
            .O(N__38849),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ));
    LocalMux I__7523 (
            .O(N__38844),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ));
    CascadeMux I__7522 (
            .O(N__38839),
            .I(N__38836));
    InMux I__7521 (
            .O(N__38836),
            .I(N__38833));
    LocalMux I__7520 (
            .O(N__38833),
            .I(N__38830));
    Odrv4 I__7519 (
            .O(N__38830),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ));
    InMux I__7518 (
            .O(N__38827),
            .I(N__38824));
    LocalMux I__7517 (
            .O(N__38824),
            .I(elapsed_time_ns_1_RNIG23T9_0_4));
    CascadeMux I__7516 (
            .O(N__38821),
            .I(elapsed_time_ns_1_RNIG23T9_0_4_cascade_));
    InMux I__7515 (
            .O(N__38818),
            .I(N__38813));
    CascadeMux I__7514 (
            .O(N__38817),
            .I(N__38809));
    InMux I__7513 (
            .O(N__38816),
            .I(N__38804));
    LocalMux I__7512 (
            .O(N__38813),
            .I(N__38801));
    InMux I__7511 (
            .O(N__38812),
            .I(N__38798));
    InMux I__7510 (
            .O(N__38809),
            .I(N__38791));
    InMux I__7509 (
            .O(N__38808),
            .I(N__38791));
    InMux I__7508 (
            .O(N__38807),
            .I(N__38791));
    LocalMux I__7507 (
            .O(N__38804),
            .I(N__38786));
    Span4Mux_v I__7506 (
            .O(N__38801),
            .I(N__38786));
    LocalMux I__7505 (
            .O(N__38798),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    LocalMux I__7504 (
            .O(N__38791),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    Odrv4 I__7503 (
            .O(N__38786),
            .I(\phase_controller_inst1.stoper_hc.start_latchedZ0 ));
    InMux I__7502 (
            .O(N__38779),
            .I(N__38776));
    LocalMux I__7501 (
            .O(N__38776),
            .I(N__38772));
    InMux I__7500 (
            .O(N__38775),
            .I(N__38769));
    Span4Mux_v I__7499 (
            .O(N__38772),
            .I(N__38764));
    LocalMux I__7498 (
            .O(N__38769),
            .I(N__38764));
    Span4Mux_v I__7497 (
            .O(N__38764),
            .I(N__38760));
    InMux I__7496 (
            .O(N__38763),
            .I(N__38757));
    Odrv4 I__7495 (
            .O(N__38760),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ));
    LocalMux I__7494 (
            .O(N__38757),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ));
    CascadeMux I__7493 (
            .O(N__38752),
            .I(N__38748));
    InMux I__7492 (
            .O(N__38751),
            .I(N__38745));
    InMux I__7491 (
            .O(N__38748),
            .I(N__38742));
    LocalMux I__7490 (
            .O(N__38745),
            .I(\phase_controller_inst1.stoper_hc.counter ));
    LocalMux I__7489 (
            .O(N__38742),
            .I(\phase_controller_inst1.stoper_hc.counter ));
    InMux I__7488 (
            .O(N__38737),
            .I(N__38732));
    InMux I__7487 (
            .O(N__38736),
            .I(N__38727));
    InMux I__7486 (
            .O(N__38735),
            .I(N__38727));
    LocalMux I__7485 (
            .O(N__38732),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ));
    LocalMux I__7484 (
            .O(N__38727),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ));
    CascadeMux I__7483 (
            .O(N__38722),
            .I(N__38717));
    CascadeMux I__7482 (
            .O(N__38721),
            .I(N__38714));
    InMux I__7481 (
            .O(N__38720),
            .I(N__38711));
    InMux I__7480 (
            .O(N__38717),
            .I(N__38706));
    InMux I__7479 (
            .O(N__38714),
            .I(N__38706));
    LocalMux I__7478 (
            .O(N__38711),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ));
    LocalMux I__7477 (
            .O(N__38706),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ));
    CascadeMux I__7476 (
            .O(N__38701),
            .I(N__38698));
    InMux I__7475 (
            .O(N__38698),
            .I(N__38695));
    LocalMux I__7474 (
            .O(N__38695),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt20 ));
    InMux I__7473 (
            .O(N__38692),
            .I(N__38686));
    InMux I__7472 (
            .O(N__38691),
            .I(N__38686));
    LocalMux I__7471 (
            .O(N__38686),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ));
    InMux I__7470 (
            .O(N__38683),
            .I(N__38677));
    InMux I__7469 (
            .O(N__38682),
            .I(N__38677));
    LocalMux I__7468 (
            .O(N__38677),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ));
    CascadeMux I__7467 (
            .O(N__38674),
            .I(N__38671));
    InMux I__7466 (
            .O(N__38671),
            .I(N__38668));
    LocalMux I__7465 (
            .O(N__38668),
            .I(N__38665));
    Odrv12 I__7464 (
            .O(N__38665),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt22 ));
    InMux I__7463 (
            .O(N__38662),
            .I(N__38659));
    LocalMux I__7462 (
            .O(N__38659),
            .I(N__38656));
    Span4Mux_h I__7461 (
            .O(N__38656),
            .I(N__38653));
    Odrv4 I__7460 (
            .O(N__38653),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt28 ));
    CascadeMux I__7459 (
            .O(N__38650),
            .I(N__38647));
    InMux I__7458 (
            .O(N__38647),
            .I(N__38644));
    LocalMux I__7457 (
            .O(N__38644),
            .I(N__38641));
    Span12Mux_h I__7456 (
            .O(N__38641),
            .I(N__38638));
    Odrv12 I__7455 (
            .O(N__38638),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ));
    InMux I__7454 (
            .O(N__38635),
            .I(N__38632));
    LocalMux I__7453 (
            .O(N__38632),
            .I(N__38629));
    Span4Mux_h I__7452 (
            .O(N__38629),
            .I(N__38626));
    Span4Mux_h I__7451 (
            .O(N__38626),
            .I(N__38623));
    Odrv4 I__7450 (
            .O(N__38623),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt30 ));
    CascadeMux I__7449 (
            .O(N__38620),
            .I(N__38617));
    InMux I__7448 (
            .O(N__38617),
            .I(N__38614));
    LocalMux I__7447 (
            .O(N__38614),
            .I(N__38611));
    Span4Mux_v I__7446 (
            .O(N__38611),
            .I(N__38608));
    Odrv4 I__7445 (
            .O(N__38608),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ));
    InMux I__7444 (
            .O(N__38605),
            .I(bfn_14_8_0_));
    InMux I__7443 (
            .O(N__38602),
            .I(N__38599));
    LocalMux I__7442 (
            .O(N__38599),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ));
    InMux I__7441 (
            .O(N__38596),
            .I(N__38593));
    LocalMux I__7440 (
            .O(N__38593),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt16 ));
    InMux I__7439 (
            .O(N__38590),
            .I(N__38587));
    LocalMux I__7438 (
            .O(N__38587),
            .I(N__38583));
    InMux I__7437 (
            .O(N__38586),
            .I(N__38580));
    Span4Mux_v I__7436 (
            .O(N__38583),
            .I(N__38577));
    LocalMux I__7435 (
            .O(N__38580),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ));
    Odrv4 I__7434 (
            .O(N__38577),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ));
    CascadeMux I__7433 (
            .O(N__38572),
            .I(N__38569));
    InMux I__7432 (
            .O(N__38569),
            .I(N__38566));
    LocalMux I__7431 (
            .O(N__38566),
            .I(\phase_controller_inst1.stoper_hc.counter_i_10 ));
    InMux I__7430 (
            .O(N__38563),
            .I(N__38559));
    InMux I__7429 (
            .O(N__38562),
            .I(N__38556));
    LocalMux I__7428 (
            .O(N__38559),
            .I(N__38553));
    LocalMux I__7427 (
            .O(N__38556),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ));
    Odrv4 I__7426 (
            .O(N__38553),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ));
    CascadeMux I__7425 (
            .O(N__38548),
            .I(N__38545));
    InMux I__7424 (
            .O(N__38545),
            .I(N__38542));
    LocalMux I__7423 (
            .O(N__38542),
            .I(\phase_controller_inst1.stoper_hc.counter_i_11 ));
    InMux I__7422 (
            .O(N__38539),
            .I(N__38535));
    InMux I__7421 (
            .O(N__38538),
            .I(N__38532));
    LocalMux I__7420 (
            .O(N__38535),
            .I(N__38529));
    LocalMux I__7419 (
            .O(N__38532),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ));
    Odrv4 I__7418 (
            .O(N__38529),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ));
    InMux I__7417 (
            .O(N__38524),
            .I(N__38521));
    LocalMux I__7416 (
            .O(N__38521),
            .I(\phase_controller_inst1.stoper_hc.counter_i_12 ));
    InMux I__7415 (
            .O(N__38518),
            .I(N__38515));
    LocalMux I__7414 (
            .O(N__38515),
            .I(N__38511));
    InMux I__7413 (
            .O(N__38514),
            .I(N__38508));
    Span4Mux_v I__7412 (
            .O(N__38511),
            .I(N__38505));
    LocalMux I__7411 (
            .O(N__38508),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ));
    Odrv4 I__7410 (
            .O(N__38505),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ));
    CascadeMux I__7409 (
            .O(N__38500),
            .I(N__38497));
    InMux I__7408 (
            .O(N__38497),
            .I(N__38494));
    LocalMux I__7407 (
            .O(N__38494),
            .I(N__38491));
    Odrv4 I__7406 (
            .O(N__38491),
            .I(\phase_controller_inst1.stoper_hc.counter_i_13 ));
    InMux I__7405 (
            .O(N__38488),
            .I(N__38484));
    InMux I__7404 (
            .O(N__38487),
            .I(N__38481));
    LocalMux I__7403 (
            .O(N__38484),
            .I(N__38478));
    LocalMux I__7402 (
            .O(N__38481),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ));
    Odrv4 I__7401 (
            .O(N__38478),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ));
    CascadeMux I__7400 (
            .O(N__38473),
            .I(N__38470));
    InMux I__7399 (
            .O(N__38470),
            .I(N__38467));
    LocalMux I__7398 (
            .O(N__38467),
            .I(\phase_controller_inst1.stoper_hc.counter_i_14 ));
    InMux I__7397 (
            .O(N__38464),
            .I(N__38461));
    LocalMux I__7396 (
            .O(N__38461),
            .I(N__38457));
    InMux I__7395 (
            .O(N__38460),
            .I(N__38454));
    Span4Mux_h I__7394 (
            .O(N__38457),
            .I(N__38451));
    LocalMux I__7393 (
            .O(N__38454),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ));
    Odrv4 I__7392 (
            .O(N__38451),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ));
    CascadeMux I__7391 (
            .O(N__38446),
            .I(N__38443));
    InMux I__7390 (
            .O(N__38443),
            .I(N__38440));
    LocalMux I__7389 (
            .O(N__38440),
            .I(\phase_controller_inst1.stoper_hc.counter_i_15 ));
    InMux I__7388 (
            .O(N__38437),
            .I(N__38434));
    LocalMux I__7387 (
            .O(N__38434),
            .I(\phase_controller_inst1.stoper_hc.un6_running_lt18 ));
    CascadeMux I__7386 (
            .O(N__38431),
            .I(N__38428));
    InMux I__7385 (
            .O(N__38428),
            .I(N__38425));
    LocalMux I__7384 (
            .O(N__38425),
            .I(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ));
    InMux I__7383 (
            .O(N__38422),
            .I(N__38418));
    InMux I__7382 (
            .O(N__38421),
            .I(N__38415));
    LocalMux I__7381 (
            .O(N__38418),
            .I(N__38412));
    LocalMux I__7380 (
            .O(N__38415),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ));
    Odrv4 I__7379 (
            .O(N__38412),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ));
    InMux I__7378 (
            .O(N__38407),
            .I(N__38404));
    LocalMux I__7377 (
            .O(N__38404),
            .I(\phase_controller_inst1.stoper_hc.counter_i_2 ));
    InMux I__7376 (
            .O(N__38401),
            .I(N__38398));
    LocalMux I__7375 (
            .O(N__38398),
            .I(N__38394));
    InMux I__7374 (
            .O(N__38397),
            .I(N__38391));
    Span4Mux_v I__7373 (
            .O(N__38394),
            .I(N__38388));
    LocalMux I__7372 (
            .O(N__38391),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ));
    Odrv4 I__7371 (
            .O(N__38388),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ));
    CascadeMux I__7370 (
            .O(N__38383),
            .I(N__38380));
    InMux I__7369 (
            .O(N__38380),
            .I(N__38377));
    LocalMux I__7368 (
            .O(N__38377),
            .I(\phase_controller_inst1.stoper_hc.counter_i_3 ));
    InMux I__7367 (
            .O(N__38374),
            .I(N__38370));
    InMux I__7366 (
            .O(N__38373),
            .I(N__38367));
    LocalMux I__7365 (
            .O(N__38370),
            .I(N__38364));
    LocalMux I__7364 (
            .O(N__38367),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ));
    Odrv4 I__7363 (
            .O(N__38364),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ));
    InMux I__7362 (
            .O(N__38359),
            .I(N__38356));
    LocalMux I__7361 (
            .O(N__38356),
            .I(\phase_controller_inst1.stoper_hc.counter_i_4 ));
    InMux I__7360 (
            .O(N__38353),
            .I(N__38350));
    LocalMux I__7359 (
            .O(N__38350),
            .I(N__38346));
    InMux I__7358 (
            .O(N__38349),
            .I(N__38343));
    Span4Mux_h I__7357 (
            .O(N__38346),
            .I(N__38340));
    LocalMux I__7356 (
            .O(N__38343),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ));
    Odrv4 I__7355 (
            .O(N__38340),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ));
    CascadeMux I__7354 (
            .O(N__38335),
            .I(N__38332));
    InMux I__7353 (
            .O(N__38332),
            .I(N__38329));
    LocalMux I__7352 (
            .O(N__38329),
            .I(\phase_controller_inst1.stoper_hc.counter_i_5 ));
    InMux I__7351 (
            .O(N__38326),
            .I(N__38323));
    LocalMux I__7350 (
            .O(N__38323),
            .I(N__38319));
    InMux I__7349 (
            .O(N__38322),
            .I(N__38316));
    Span4Mux_v I__7348 (
            .O(N__38319),
            .I(N__38313));
    LocalMux I__7347 (
            .O(N__38316),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ));
    Odrv4 I__7346 (
            .O(N__38313),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ));
    InMux I__7345 (
            .O(N__38308),
            .I(N__38305));
    LocalMux I__7344 (
            .O(N__38305),
            .I(\phase_controller_inst1.stoper_hc.counter_i_6 ));
    InMux I__7343 (
            .O(N__38302),
            .I(N__38298));
    InMux I__7342 (
            .O(N__38301),
            .I(N__38295));
    LocalMux I__7341 (
            .O(N__38298),
            .I(N__38292));
    LocalMux I__7340 (
            .O(N__38295),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ));
    Odrv4 I__7339 (
            .O(N__38292),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ));
    CascadeMux I__7338 (
            .O(N__38287),
            .I(N__38284));
    InMux I__7337 (
            .O(N__38284),
            .I(N__38281));
    LocalMux I__7336 (
            .O(N__38281),
            .I(N__38278));
    Odrv4 I__7335 (
            .O(N__38278),
            .I(\phase_controller_inst1.stoper_hc.counter_i_7 ));
    InMux I__7334 (
            .O(N__38275),
            .I(N__38272));
    LocalMux I__7333 (
            .O(N__38272),
            .I(N__38268));
    InMux I__7332 (
            .O(N__38271),
            .I(N__38265));
    Span4Mux_h I__7331 (
            .O(N__38268),
            .I(N__38262));
    LocalMux I__7330 (
            .O(N__38265),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ));
    Odrv4 I__7329 (
            .O(N__38262),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ));
    CascadeMux I__7328 (
            .O(N__38257),
            .I(N__38254));
    InMux I__7327 (
            .O(N__38254),
            .I(N__38251));
    LocalMux I__7326 (
            .O(N__38251),
            .I(\phase_controller_inst1.stoper_hc.counter_i_8 ));
    InMux I__7325 (
            .O(N__38248),
            .I(N__38244));
    InMux I__7324 (
            .O(N__38247),
            .I(N__38241));
    LocalMux I__7323 (
            .O(N__38244),
            .I(N__38238));
    LocalMux I__7322 (
            .O(N__38241),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ));
    Odrv4 I__7321 (
            .O(N__38238),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ));
    CascadeMux I__7320 (
            .O(N__38233),
            .I(N__38230));
    InMux I__7319 (
            .O(N__38230),
            .I(N__38227));
    LocalMux I__7318 (
            .O(N__38227),
            .I(\phase_controller_inst1.stoper_hc.counter_i_9 ));
    InMux I__7317 (
            .O(N__38224),
            .I(N__38221));
    LocalMux I__7316 (
            .O(N__38221),
            .I(N__38218));
    Odrv4 I__7315 (
            .O(N__38218),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_31 ));
    InMux I__7314 (
            .O(N__38215),
            .I(N__38212));
    LocalMux I__7313 (
            .O(N__38212),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ));
    InMux I__7312 (
            .O(N__38209),
            .I(N__38206));
    LocalMux I__7311 (
            .O(N__38206),
            .I(N__38202));
    InMux I__7310 (
            .O(N__38205),
            .I(N__38199));
    Span12Mux_v I__7309 (
            .O(N__38202),
            .I(N__38196));
    LocalMux I__7308 (
            .O(N__38199),
            .I(N__38191));
    Span12Mux_h I__7307 (
            .O(N__38196),
            .I(N__38191));
    Odrv12 I__7306 (
            .O(N__38191),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_25 ));
    InMux I__7305 (
            .O(N__38188),
            .I(N__38185));
    LocalMux I__7304 (
            .O(N__38185),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ));
    InMux I__7303 (
            .O(N__38182),
            .I(N__38178));
    InMux I__7302 (
            .O(N__38181),
            .I(N__38175));
    LocalMux I__7301 (
            .O(N__38178),
            .I(N__38172));
    LocalMux I__7300 (
            .O(N__38175),
            .I(N__38169));
    Span12Mux_s10_v I__7299 (
            .O(N__38172),
            .I(N__38166));
    Odrv4 I__7298 (
            .O(N__38169),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    Odrv12 I__7297 (
            .O(N__38166),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_28 ));
    InMux I__7296 (
            .O(N__38161),
            .I(N__38158));
    LocalMux I__7295 (
            .O(N__38158),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ));
    CascadeMux I__7294 (
            .O(N__38155),
            .I(N__38151));
    InMux I__7293 (
            .O(N__38154),
            .I(N__38143));
    InMux I__7292 (
            .O(N__38151),
            .I(N__38143));
    InMux I__7291 (
            .O(N__38150),
            .I(N__38143));
    LocalMux I__7290 (
            .O(N__38143),
            .I(N__38140));
    Odrv12 I__7289 (
            .O(N__38140),
            .I(\delay_measurement_inst.stop_timer_trZ0 ));
    InMux I__7288 (
            .O(N__38137),
            .I(N__38131));
    InMux I__7287 (
            .O(N__38136),
            .I(N__38131));
    LocalMux I__7286 (
            .O(N__38131),
            .I(N__38128));
    Span4Mux_v I__7285 (
            .O(N__38128),
            .I(N__38123));
    InMux I__7284 (
            .O(N__38127),
            .I(N__38118));
    InMux I__7283 (
            .O(N__38126),
            .I(N__38118));
    Span4Mux_v I__7282 (
            .O(N__38123),
            .I(N__38115));
    LocalMux I__7281 (
            .O(N__38118),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    Odrv4 I__7280 (
            .O(N__38115),
            .I(\delay_measurement_inst.start_timer_trZ0 ));
    ClkMux I__7279 (
            .O(N__38110),
            .I(N__38107));
    GlobalMux I__7278 (
            .O(N__38107),
            .I(N__38104));
    gio2CtrlBuf I__7277 (
            .O(N__38104),
            .I(delay_tr_input_c_g));
    InMux I__7276 (
            .O(N__38101),
            .I(N__38097));
    CascadeMux I__7275 (
            .O(N__38100),
            .I(N__38092));
    LocalMux I__7274 (
            .O(N__38097),
            .I(N__38089));
    InMux I__7273 (
            .O(N__38096),
            .I(N__38084));
    InMux I__7272 (
            .O(N__38095),
            .I(N__38084));
    InMux I__7271 (
            .O(N__38092),
            .I(N__38081));
    Span12Mux_v I__7270 (
            .O(N__38089),
            .I(N__38078));
    LocalMux I__7269 (
            .O(N__38084),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    LocalMux I__7268 (
            .O(N__38081),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    Odrv12 I__7267 (
            .O(N__38078),
            .I(\phase_controller_inst1.stateZ0Z_1 ));
    IoInMux I__7266 (
            .O(N__38071),
            .I(N__38068));
    LocalMux I__7265 (
            .O(N__38068),
            .I(N__38065));
    Odrv12 I__7264 (
            .O(N__38065),
            .I(s2_phy_c));
    InMux I__7263 (
            .O(N__38062),
            .I(N__38059));
    LocalMux I__7262 (
            .O(N__38059),
            .I(N__38055));
    InMux I__7261 (
            .O(N__38058),
            .I(N__38052));
    Span4Mux_h I__7260 (
            .O(N__38055),
            .I(N__38049));
    LocalMux I__7259 (
            .O(N__38052),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ));
    Odrv4 I__7258 (
            .O(N__38049),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ));
    CascadeMux I__7257 (
            .O(N__38044),
            .I(N__38041));
    InMux I__7256 (
            .O(N__38041),
            .I(N__38038));
    LocalMux I__7255 (
            .O(N__38038),
            .I(\phase_controller_inst1.stoper_hc.counter_i_0 ));
    InMux I__7254 (
            .O(N__38035),
            .I(N__38032));
    LocalMux I__7253 (
            .O(N__38032),
            .I(N__38028));
    InMux I__7252 (
            .O(N__38031),
            .I(N__38025));
    Span4Mux_h I__7251 (
            .O(N__38028),
            .I(N__38022));
    LocalMux I__7250 (
            .O(N__38025),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ));
    Odrv4 I__7249 (
            .O(N__38022),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ));
    CascadeMux I__7248 (
            .O(N__38017),
            .I(N__38014));
    InMux I__7247 (
            .O(N__38014),
            .I(N__38011));
    LocalMux I__7246 (
            .O(N__38011),
            .I(\phase_controller_inst1.stoper_hc.counter_i_1 ));
    InMux I__7245 (
            .O(N__38008),
            .I(N__38005));
    LocalMux I__7244 (
            .O(N__38005),
            .I(N__38001));
    InMux I__7243 (
            .O(N__38004),
            .I(N__37998));
    Span4Mux_s2_h I__7242 (
            .O(N__38001),
            .I(N__37995));
    LocalMux I__7241 (
            .O(N__37998),
            .I(N__37992));
    Sp12to4 I__7240 (
            .O(N__37995),
            .I(N__37989));
    Span4Mux_v I__7239 (
            .O(N__37992),
            .I(N__37986));
    Span12Mux_s11_v I__7238 (
            .O(N__37989),
            .I(N__37983));
    Odrv4 I__7237 (
            .O(N__37986),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    Odrv12 I__7236 (
            .O(N__37983),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_22 ));
    CascadeMux I__7235 (
            .O(N__37978),
            .I(N__37975));
    InMux I__7234 (
            .O(N__37975),
            .I(N__37972));
    LocalMux I__7233 (
            .O(N__37972),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ));
    InMux I__7232 (
            .O(N__37969),
            .I(N__37966));
    LocalMux I__7231 (
            .O(N__37966),
            .I(N__37963));
    Span4Mux_v I__7230 (
            .O(N__37963),
            .I(N__37959));
    InMux I__7229 (
            .O(N__37962),
            .I(N__37956));
    Sp12to4 I__7228 (
            .O(N__37959),
            .I(N__37953));
    LocalMux I__7227 (
            .O(N__37956),
            .I(N__37948));
    Span12Mux_h I__7226 (
            .O(N__37953),
            .I(N__37948));
    Odrv12 I__7225 (
            .O(N__37948),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_23 ));
    InMux I__7224 (
            .O(N__37945),
            .I(N__37942));
    LocalMux I__7223 (
            .O(N__37942),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ));
    InMux I__7222 (
            .O(N__37939),
            .I(N__37935));
    InMux I__7221 (
            .O(N__37938),
            .I(N__37932));
    LocalMux I__7220 (
            .O(N__37935),
            .I(N__37929));
    LocalMux I__7219 (
            .O(N__37932),
            .I(N__37926));
    Span12Mux_s11_v I__7218 (
            .O(N__37929),
            .I(N__37923));
    Odrv4 I__7217 (
            .O(N__37926),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    Odrv12 I__7216 (
            .O(N__37923),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_20 ));
    InMux I__7215 (
            .O(N__37918),
            .I(N__37915));
    LocalMux I__7214 (
            .O(N__37915),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ));
    InMux I__7213 (
            .O(N__37912),
            .I(N__37909));
    LocalMux I__7212 (
            .O(N__37909),
            .I(N__37905));
    InMux I__7211 (
            .O(N__37908),
            .I(N__37902));
    Span12Mux_s6_v I__7210 (
            .O(N__37905),
            .I(N__37899));
    LocalMux I__7209 (
            .O(N__37902),
            .I(N__37896));
    Span12Mux_h I__7208 (
            .O(N__37899),
            .I(N__37893));
    Odrv4 I__7207 (
            .O(N__37896),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    Odrv12 I__7206 (
            .O(N__37893),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_21 ));
    InMux I__7205 (
            .O(N__37888),
            .I(N__37885));
    LocalMux I__7204 (
            .O(N__37885),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ));
    InMux I__7203 (
            .O(N__37882),
            .I(N__37879));
    LocalMux I__7202 (
            .O(N__37879),
            .I(N__37875));
    InMux I__7201 (
            .O(N__37878),
            .I(N__37872));
    Span12Mux_v I__7200 (
            .O(N__37875),
            .I(N__37869));
    LocalMux I__7199 (
            .O(N__37872),
            .I(N__37864));
    Span12Mux_h I__7198 (
            .O(N__37869),
            .I(N__37864));
    Odrv12 I__7197 (
            .O(N__37864),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_30 ));
    InMux I__7196 (
            .O(N__37861),
            .I(N__37858));
    LocalMux I__7195 (
            .O(N__37858),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ));
    InMux I__7194 (
            .O(N__37855),
            .I(N__37852));
    LocalMux I__7193 (
            .O(N__37852),
            .I(N__37849));
    Span4Mux_s1_h I__7192 (
            .O(N__37849),
            .I(N__37845));
    InMux I__7191 (
            .O(N__37848),
            .I(N__37842));
    Sp12to4 I__7190 (
            .O(N__37845),
            .I(N__37839));
    LocalMux I__7189 (
            .O(N__37842),
            .I(N__37836));
    Span12Mux_s10_v I__7188 (
            .O(N__37839),
            .I(N__37833));
    Odrv4 I__7187 (
            .O(N__37836),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    Odrv12 I__7186 (
            .O(N__37833),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_29 ));
    InMux I__7185 (
            .O(N__37828),
            .I(N__37825));
    LocalMux I__7184 (
            .O(N__37825),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ));
    InMux I__7183 (
            .O(N__37822),
            .I(N__37818));
    InMux I__7182 (
            .O(N__37821),
            .I(N__37815));
    LocalMux I__7181 (
            .O(N__37818),
            .I(N__37812));
    LocalMux I__7180 (
            .O(N__37815),
            .I(N__37807));
    Span12Mux_s7_v I__7179 (
            .O(N__37812),
            .I(N__37807));
    Span12Mux_h I__7178 (
            .O(N__37807),
            .I(N__37804));
    Odrv12 I__7177 (
            .O(N__37804),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_27 ));
    InMux I__7176 (
            .O(N__37801),
            .I(N__37798));
    LocalMux I__7175 (
            .O(N__37798),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ));
    InMux I__7174 (
            .O(N__37795),
            .I(N__37792));
    LocalMux I__7173 (
            .O(N__37792),
            .I(N__37789));
    Sp12to4 I__7172 (
            .O(N__37789),
            .I(N__37785));
    InMux I__7171 (
            .O(N__37788),
            .I(N__37782));
    Span12Mux_v I__7170 (
            .O(N__37785),
            .I(N__37779));
    LocalMux I__7169 (
            .O(N__37782),
            .I(N__37774));
    Span12Mux_h I__7168 (
            .O(N__37779),
            .I(N__37774));
    Odrv12 I__7167 (
            .O(N__37774),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_26 ));
    InMux I__7166 (
            .O(N__37771),
            .I(N__37768));
    LocalMux I__7165 (
            .O(N__37768),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ));
    InMux I__7164 (
            .O(N__37765),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ));
    InMux I__7163 (
            .O(N__37762),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ));
    InMux I__7162 (
            .O(N__37759),
            .I(N__37753));
    InMux I__7161 (
            .O(N__37758),
            .I(N__37753));
    LocalMux I__7160 (
            .O(N__37753),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ));
    InMux I__7159 (
            .O(N__37750),
            .I(N__37744));
    InMux I__7158 (
            .O(N__37749),
            .I(N__37744));
    LocalMux I__7157 (
            .O(N__37744),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ));
    InMux I__7156 (
            .O(N__37741),
            .I(N__37735));
    InMux I__7155 (
            .O(N__37740),
            .I(N__37735));
    LocalMux I__7154 (
            .O(N__37735),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ));
    CascadeMux I__7153 (
            .O(N__37732),
            .I(N__37728));
    InMux I__7152 (
            .O(N__37731),
            .I(N__37723));
    InMux I__7151 (
            .O(N__37728),
            .I(N__37723));
    LocalMux I__7150 (
            .O(N__37723),
            .I(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ));
    CascadeMux I__7149 (
            .O(N__37720),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ));
    InMux I__7148 (
            .O(N__37717),
            .I(N__37714));
    LocalMux I__7147 (
            .O(N__37714),
            .I(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ));
    CascadeMux I__7146 (
            .O(N__37711),
            .I(N__37708));
    InMux I__7145 (
            .O(N__37708),
            .I(N__37705));
    LocalMux I__7144 (
            .O(N__37705),
            .I(N__37700));
    CascadeMux I__7143 (
            .O(N__37704),
            .I(N__37697));
    InMux I__7142 (
            .O(N__37703),
            .I(N__37693));
    Span4Mux_h I__7141 (
            .O(N__37700),
            .I(N__37690));
    InMux I__7140 (
            .O(N__37697),
            .I(N__37687));
    InMux I__7139 (
            .O(N__37696),
            .I(N__37684));
    LocalMux I__7138 (
            .O(N__37693),
            .I(N__37681));
    Odrv4 I__7137 (
            .O(N__37690),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__7136 (
            .O(N__37687),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    LocalMux I__7135 (
            .O(N__37684),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    Odrv4 I__7134 (
            .O(N__37681),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ));
    CascadeMux I__7133 (
            .O(N__37672),
            .I(N__37668));
    InMux I__7132 (
            .O(N__37671),
            .I(N__37664));
    InMux I__7131 (
            .O(N__37668),
            .I(N__37661));
    InMux I__7130 (
            .O(N__37667),
            .I(N__37658));
    LocalMux I__7129 (
            .O(N__37664),
            .I(N__37654));
    LocalMux I__7128 (
            .O(N__37661),
            .I(N__37651));
    LocalMux I__7127 (
            .O(N__37658),
            .I(N__37648));
    InMux I__7126 (
            .O(N__37657),
            .I(N__37645));
    Span4Mux_h I__7125 (
            .O(N__37654),
            .I(N__37642));
    Odrv4 I__7124 (
            .O(N__37651),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv12 I__7123 (
            .O(N__37648),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    LocalMux I__7122 (
            .O(N__37645),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    Odrv4 I__7121 (
            .O(N__37642),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ));
    CascadeMux I__7120 (
            .O(N__37633),
            .I(N__37629));
    CascadeMux I__7119 (
            .O(N__37632),
            .I(N__37626));
    InMux I__7118 (
            .O(N__37629),
            .I(N__37623));
    InMux I__7117 (
            .O(N__37626),
            .I(N__37620));
    LocalMux I__7116 (
            .O(N__37623),
            .I(N__37616));
    LocalMux I__7115 (
            .O(N__37620),
            .I(N__37613));
    CascadeMux I__7114 (
            .O(N__37619),
            .I(N__37610));
    Span4Mux_v I__7113 (
            .O(N__37616),
            .I(N__37606));
    Span4Mux_h I__7112 (
            .O(N__37613),
            .I(N__37603));
    InMux I__7111 (
            .O(N__37610),
            .I(N__37600));
    InMux I__7110 (
            .O(N__37609),
            .I(N__37597));
    Span4Mux_h I__7109 (
            .O(N__37606),
            .I(N__37594));
    Odrv4 I__7108 (
            .O(N__37603),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__7107 (
            .O(N__37600),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    LocalMux I__7106 (
            .O(N__37597),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    Odrv4 I__7105 (
            .O(N__37594),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ));
    InMux I__7104 (
            .O(N__37585),
            .I(N__37581));
    InMux I__7103 (
            .O(N__37584),
            .I(N__37576));
    LocalMux I__7102 (
            .O(N__37581),
            .I(N__37573));
    CascadeMux I__7101 (
            .O(N__37580),
            .I(N__37570));
    CascadeMux I__7100 (
            .O(N__37579),
            .I(N__37567));
    LocalMux I__7099 (
            .O(N__37576),
            .I(N__37564));
    Span4Mux_h I__7098 (
            .O(N__37573),
            .I(N__37561));
    InMux I__7097 (
            .O(N__37570),
            .I(N__37558));
    InMux I__7096 (
            .O(N__37567),
            .I(N__37555));
    Span4Mux_h I__7095 (
            .O(N__37564),
            .I(N__37552));
    Odrv4 I__7094 (
            .O(N__37561),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__7093 (
            .O(N__37558),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    LocalMux I__7092 (
            .O(N__37555),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    Odrv4 I__7091 (
            .O(N__37552),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ));
    InMux I__7090 (
            .O(N__37543),
            .I(N__37540));
    LocalMux I__7089 (
            .O(N__37540),
            .I(N__37537));
    Span4Mux_h I__7088 (
            .O(N__37537),
            .I(N__37534));
    Odrv4 I__7087 (
            .O(N__37534),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ));
    InMux I__7086 (
            .O(N__37531),
            .I(N__37528));
    LocalMux I__7085 (
            .O(N__37528),
            .I(N__37524));
    InMux I__7084 (
            .O(N__37527),
            .I(N__37521));
    Span12Mux_v I__7083 (
            .O(N__37524),
            .I(N__37518));
    LocalMux I__7082 (
            .O(N__37521),
            .I(N__37513));
    Span12Mux_h I__7081 (
            .O(N__37518),
            .I(N__37513));
    Odrv12 I__7080 (
            .O(N__37513),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_18 ));
    InMux I__7079 (
            .O(N__37510),
            .I(N__37507));
    LocalMux I__7078 (
            .O(N__37507),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ));
    InMux I__7077 (
            .O(N__37504),
            .I(N__37501));
    LocalMux I__7076 (
            .O(N__37501),
            .I(N__37498));
    Span4Mux_s3_h I__7075 (
            .O(N__37498),
            .I(N__37494));
    InMux I__7074 (
            .O(N__37497),
            .I(N__37491));
    Span4Mux_h I__7073 (
            .O(N__37494),
            .I(N__37488));
    LocalMux I__7072 (
            .O(N__37491),
            .I(N__37483));
    Span4Mux_h I__7071 (
            .O(N__37488),
            .I(N__37483));
    Span4Mux_v I__7070 (
            .O(N__37483),
            .I(N__37480));
    Odrv4 I__7069 (
            .O(N__37480),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_24 ));
    InMux I__7068 (
            .O(N__37477),
            .I(N__37474));
    LocalMux I__7067 (
            .O(N__37474),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ));
    InMux I__7066 (
            .O(N__37471),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ));
    InMux I__7065 (
            .O(N__37468),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ));
    InMux I__7064 (
            .O(N__37465),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ));
    InMux I__7063 (
            .O(N__37462),
            .I(bfn_13_20_0_));
    InMux I__7062 (
            .O(N__37459),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ));
    InMux I__7061 (
            .O(N__37456),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ));
    InMux I__7060 (
            .O(N__37453),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ));
    InMux I__7059 (
            .O(N__37450),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ));
    InMux I__7058 (
            .O(N__37447),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ));
    InMux I__7057 (
            .O(N__37444),
            .I(N__37441));
    LocalMux I__7056 (
            .O(N__37441),
            .I(N__37438));
    Span4Mux_v I__7055 (
            .O(N__37438),
            .I(N__37435));
    Sp12to4 I__7054 (
            .O(N__37435),
            .I(N__37431));
    InMux I__7053 (
            .O(N__37434),
            .I(N__37428));
    Span12Mux_h I__7052 (
            .O(N__37431),
            .I(N__37425));
    LocalMux I__7051 (
            .O(N__37428),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    Odrv12 I__7050 (
            .O(N__37425),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_12 ));
    InMux I__7049 (
            .O(N__37420),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ));
    InMux I__7048 (
            .O(N__37417),
            .I(N__37414));
    LocalMux I__7047 (
            .O(N__37414),
            .I(N__37411));
    Span4Mux_v I__7046 (
            .O(N__37411),
            .I(N__37408));
    Sp12to4 I__7045 (
            .O(N__37408),
            .I(N__37405));
    Span12Mux_h I__7044 (
            .O(N__37405),
            .I(N__37401));
    InMux I__7043 (
            .O(N__37404),
            .I(N__37398));
    Span12Mux_v I__7042 (
            .O(N__37401),
            .I(N__37395));
    LocalMux I__7041 (
            .O(N__37398),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    Odrv12 I__7040 (
            .O(N__37395),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_13 ));
    InMux I__7039 (
            .O(N__37390),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ));
    InMux I__7038 (
            .O(N__37387),
            .I(N__37384));
    LocalMux I__7037 (
            .O(N__37384),
            .I(N__37381));
    Span4Mux_v I__7036 (
            .O(N__37381),
            .I(N__37378));
    Sp12to4 I__7035 (
            .O(N__37378),
            .I(N__37375));
    Span12Mux_s11_h I__7034 (
            .O(N__37375),
            .I(N__37371));
    InMux I__7033 (
            .O(N__37374),
            .I(N__37368));
    Span12Mux_v I__7032 (
            .O(N__37371),
            .I(N__37365));
    LocalMux I__7031 (
            .O(N__37368),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    Odrv12 I__7030 (
            .O(N__37365),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_14 ));
    InMux I__7029 (
            .O(N__37360),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ));
    InMux I__7028 (
            .O(N__37357),
            .I(N__37354));
    LocalMux I__7027 (
            .O(N__37354),
            .I(N__37351));
    Sp12to4 I__7026 (
            .O(N__37351),
            .I(N__37347));
    InMux I__7025 (
            .O(N__37350),
            .I(N__37344));
    Span12Mux_h I__7024 (
            .O(N__37347),
            .I(N__37341));
    LocalMux I__7023 (
            .O(N__37344),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    Odrv12 I__7022 (
            .O(N__37341),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_15 ));
    InMux I__7021 (
            .O(N__37336),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ));
    InMux I__7020 (
            .O(N__37333),
            .I(N__37330));
    LocalMux I__7019 (
            .O(N__37330),
            .I(N__37327));
    Sp12to4 I__7018 (
            .O(N__37327),
            .I(N__37324));
    Span12Mux_v I__7017 (
            .O(N__37324),
            .I(N__37320));
    InMux I__7016 (
            .O(N__37323),
            .I(N__37317));
    Span12Mux_h I__7015 (
            .O(N__37320),
            .I(N__37314));
    LocalMux I__7014 (
            .O(N__37317),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    Odrv12 I__7013 (
            .O(N__37314),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_16 ));
    InMux I__7012 (
            .O(N__37309),
            .I(bfn_13_19_0_));
    InMux I__7011 (
            .O(N__37306),
            .I(N__37303));
    LocalMux I__7010 (
            .O(N__37303),
            .I(N__37300));
    Span4Mux_v I__7009 (
            .O(N__37300),
            .I(N__37297));
    Sp12to4 I__7008 (
            .O(N__37297),
            .I(N__37293));
    InMux I__7007 (
            .O(N__37296),
            .I(N__37290));
    Span12Mux_h I__7006 (
            .O(N__37293),
            .I(N__37287));
    LocalMux I__7005 (
            .O(N__37290),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    Odrv12 I__7004 (
            .O(N__37287),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_17 ));
    InMux I__7003 (
            .O(N__37282),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ));
    InMux I__7002 (
            .O(N__37279),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ));
    InMux I__7001 (
            .O(N__37276),
            .I(N__37273));
    LocalMux I__7000 (
            .O(N__37273),
            .I(N__37270));
    Span4Mux_v I__6999 (
            .O(N__37270),
            .I(N__37267));
    Span4Mux_h I__6998 (
            .O(N__37267),
            .I(N__37264));
    Span4Mux_h I__6997 (
            .O(N__37264),
            .I(N__37260));
    InMux I__6996 (
            .O(N__37263),
            .I(N__37257));
    Span4Mux_h I__6995 (
            .O(N__37260),
            .I(N__37254));
    LocalMux I__6994 (
            .O(N__37257),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    Odrv4 I__6993 (
            .O(N__37254),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_19 ));
    InMux I__6992 (
            .O(N__37249),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ));
    InMux I__6991 (
            .O(N__37246),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ));
    InMux I__6990 (
            .O(N__37243),
            .I(N__37240));
    LocalMux I__6989 (
            .O(N__37240),
            .I(N__37237));
    Sp12to4 I__6988 (
            .O(N__37237),
            .I(N__37234));
    Span12Mux_v I__6987 (
            .O(N__37234),
            .I(N__37230));
    InMux I__6986 (
            .O(N__37233),
            .I(N__37227));
    Span12Mux_h I__6985 (
            .O(N__37230),
            .I(N__37224));
    LocalMux I__6984 (
            .O(N__37227),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    Odrv12 I__6983 (
            .O(N__37224),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_4 ));
    InMux I__6982 (
            .O(N__37219),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ));
    InMux I__6981 (
            .O(N__37216),
            .I(N__37213));
    LocalMux I__6980 (
            .O(N__37213),
            .I(N__37210));
    Sp12to4 I__6979 (
            .O(N__37210),
            .I(N__37207));
    Span12Mux_s9_v I__6978 (
            .O(N__37207),
            .I(N__37203));
    InMux I__6977 (
            .O(N__37206),
            .I(N__37200));
    Span12Mux_h I__6976 (
            .O(N__37203),
            .I(N__37197));
    LocalMux I__6975 (
            .O(N__37200),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    Odrv12 I__6974 (
            .O(N__37197),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_5 ));
    InMux I__6973 (
            .O(N__37192),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ));
    InMux I__6972 (
            .O(N__37189),
            .I(N__37186));
    LocalMux I__6971 (
            .O(N__37186),
            .I(N__37183));
    Sp12to4 I__6970 (
            .O(N__37183),
            .I(N__37180));
    Span12Mux_s10_v I__6969 (
            .O(N__37180),
            .I(N__37176));
    InMux I__6968 (
            .O(N__37179),
            .I(N__37173));
    Span12Mux_h I__6967 (
            .O(N__37176),
            .I(N__37170));
    LocalMux I__6966 (
            .O(N__37173),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    Odrv12 I__6965 (
            .O(N__37170),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_6 ));
    InMux I__6964 (
            .O(N__37165),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ));
    InMux I__6963 (
            .O(N__37162),
            .I(N__37159));
    LocalMux I__6962 (
            .O(N__37159),
            .I(N__37156));
    Span4Mux_v I__6961 (
            .O(N__37156),
            .I(N__37153));
    Sp12to4 I__6960 (
            .O(N__37153),
            .I(N__37149));
    InMux I__6959 (
            .O(N__37152),
            .I(N__37146));
    Span12Mux_s10_h I__6958 (
            .O(N__37149),
            .I(N__37143));
    LocalMux I__6957 (
            .O(N__37146),
            .I(N__37140));
    Span12Mux_v I__6956 (
            .O(N__37143),
            .I(N__37137));
    Odrv4 I__6955 (
            .O(N__37140),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    Odrv12 I__6954 (
            .O(N__37137),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_7 ));
    InMux I__6953 (
            .O(N__37132),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ));
    InMux I__6952 (
            .O(N__37129),
            .I(N__37126));
    LocalMux I__6951 (
            .O(N__37126),
            .I(N__37123));
    Span4Mux_v I__6950 (
            .O(N__37123),
            .I(N__37120));
    Sp12to4 I__6949 (
            .O(N__37120),
            .I(N__37116));
    InMux I__6948 (
            .O(N__37119),
            .I(N__37113));
    Span12Mux_h I__6947 (
            .O(N__37116),
            .I(N__37110));
    LocalMux I__6946 (
            .O(N__37113),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    Odrv12 I__6945 (
            .O(N__37110),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_8 ));
    InMux I__6944 (
            .O(N__37105),
            .I(bfn_13_18_0_));
    InMux I__6943 (
            .O(N__37102),
            .I(N__37099));
    LocalMux I__6942 (
            .O(N__37099),
            .I(N__37096));
    Span12Mux_s1_h I__6941 (
            .O(N__37096),
            .I(N__37092));
    InMux I__6940 (
            .O(N__37095),
            .I(N__37089));
    Span12Mux_h I__6939 (
            .O(N__37092),
            .I(N__37086));
    LocalMux I__6938 (
            .O(N__37089),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    Odrv12 I__6937 (
            .O(N__37086),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_9 ));
    InMux I__6936 (
            .O(N__37081),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ));
    InMux I__6935 (
            .O(N__37078),
            .I(N__37075));
    LocalMux I__6934 (
            .O(N__37075),
            .I(N__37072));
    Sp12to4 I__6933 (
            .O(N__37072),
            .I(N__37069));
    Span12Mux_s7_v I__6932 (
            .O(N__37069),
            .I(N__37065));
    InMux I__6931 (
            .O(N__37068),
            .I(N__37062));
    Span12Mux_h I__6930 (
            .O(N__37065),
            .I(N__37059));
    LocalMux I__6929 (
            .O(N__37062),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    Odrv12 I__6928 (
            .O(N__37059),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_10 ));
    InMux I__6927 (
            .O(N__37054),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ));
    InMux I__6926 (
            .O(N__37051),
            .I(N__37048));
    LocalMux I__6925 (
            .O(N__37048),
            .I(N__37045));
    Span4Mux_v I__6924 (
            .O(N__37045),
            .I(N__37042));
    Sp12to4 I__6923 (
            .O(N__37042),
            .I(N__37038));
    InMux I__6922 (
            .O(N__37041),
            .I(N__37035));
    Span12Mux_h I__6921 (
            .O(N__37038),
            .I(N__37032));
    LocalMux I__6920 (
            .O(N__37035),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    Odrv12 I__6919 (
            .O(N__37032),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_11 ));
    InMux I__6918 (
            .O(N__37027),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ));
    InMux I__6917 (
            .O(N__37024),
            .I(N__37021));
    LocalMux I__6916 (
            .O(N__37021),
            .I(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ));
    InMux I__6915 (
            .O(N__37018),
            .I(N__37015));
    LocalMux I__6914 (
            .O(N__37015),
            .I(N__37012));
    Span4Mux_v I__6913 (
            .O(N__37012),
            .I(N__37009));
    Sp12to4 I__6912 (
            .O(N__37009),
            .I(N__37005));
    InMux I__6911 (
            .O(N__37008),
            .I(N__37002));
    Span12Mux_h I__6910 (
            .O(N__37005),
            .I(N__36999));
    LocalMux I__6909 (
            .O(N__37002),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    Odrv12 I__6908 (
            .O(N__36999),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_1 ));
    InMux I__6907 (
            .O(N__36994),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ));
    InMux I__6906 (
            .O(N__36991),
            .I(N__36988));
    LocalMux I__6905 (
            .O(N__36988),
            .I(N__36985));
    Span12Mux_s1_h I__6904 (
            .O(N__36985),
            .I(N__36981));
    InMux I__6903 (
            .O(N__36984),
            .I(N__36978));
    Span12Mux_h I__6902 (
            .O(N__36981),
            .I(N__36975));
    LocalMux I__6901 (
            .O(N__36978),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    Odrv12 I__6900 (
            .O(N__36975),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_2 ));
    InMux I__6899 (
            .O(N__36970),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ));
    InMux I__6898 (
            .O(N__36967),
            .I(N__36964));
    LocalMux I__6897 (
            .O(N__36964),
            .I(N__36961));
    Sp12to4 I__6896 (
            .O(N__36961),
            .I(N__36958));
    Span12Mux_s7_v I__6895 (
            .O(N__36958),
            .I(N__36954));
    InMux I__6894 (
            .O(N__36957),
            .I(N__36951));
    Span12Mux_h I__6893 (
            .O(N__36954),
            .I(N__36948));
    LocalMux I__6892 (
            .O(N__36951),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    Odrv12 I__6891 (
            .O(N__36948),
            .I(\current_shift_inst.PI_CTRL.prop_term_1_3 ));
    InMux I__6890 (
            .O(N__36943),
            .I(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ));
    InMux I__6889 (
            .O(N__36940),
            .I(N__36900));
    InMux I__6888 (
            .O(N__36939),
            .I(N__36900));
    InMux I__6887 (
            .O(N__36938),
            .I(N__36900));
    InMux I__6886 (
            .O(N__36937),
            .I(N__36900));
    InMux I__6885 (
            .O(N__36936),
            .I(N__36891));
    InMux I__6884 (
            .O(N__36935),
            .I(N__36891));
    InMux I__6883 (
            .O(N__36934),
            .I(N__36891));
    InMux I__6882 (
            .O(N__36933),
            .I(N__36891));
    InMux I__6881 (
            .O(N__36932),
            .I(N__36882));
    InMux I__6880 (
            .O(N__36931),
            .I(N__36882));
    InMux I__6879 (
            .O(N__36930),
            .I(N__36882));
    InMux I__6878 (
            .O(N__36929),
            .I(N__36882));
    InMux I__6877 (
            .O(N__36928),
            .I(N__36875));
    InMux I__6876 (
            .O(N__36927),
            .I(N__36875));
    InMux I__6875 (
            .O(N__36926),
            .I(N__36875));
    InMux I__6874 (
            .O(N__36925),
            .I(N__36866));
    InMux I__6873 (
            .O(N__36924),
            .I(N__36866));
    InMux I__6872 (
            .O(N__36923),
            .I(N__36866));
    InMux I__6871 (
            .O(N__36922),
            .I(N__36866));
    InMux I__6870 (
            .O(N__36921),
            .I(N__36857));
    InMux I__6869 (
            .O(N__36920),
            .I(N__36857));
    InMux I__6868 (
            .O(N__36919),
            .I(N__36857));
    InMux I__6867 (
            .O(N__36918),
            .I(N__36857));
    InMux I__6866 (
            .O(N__36917),
            .I(N__36848));
    InMux I__6865 (
            .O(N__36916),
            .I(N__36848));
    InMux I__6864 (
            .O(N__36915),
            .I(N__36848));
    InMux I__6863 (
            .O(N__36914),
            .I(N__36848));
    InMux I__6862 (
            .O(N__36913),
            .I(N__36837));
    InMux I__6861 (
            .O(N__36912),
            .I(N__36837));
    InMux I__6860 (
            .O(N__36911),
            .I(N__36837));
    InMux I__6859 (
            .O(N__36910),
            .I(N__36837));
    InMux I__6858 (
            .O(N__36909),
            .I(N__36837));
    LocalMux I__6857 (
            .O(N__36900),
            .I(N__36820));
    LocalMux I__6856 (
            .O(N__36891),
            .I(N__36820));
    LocalMux I__6855 (
            .O(N__36882),
            .I(N__36820));
    LocalMux I__6854 (
            .O(N__36875),
            .I(N__36820));
    LocalMux I__6853 (
            .O(N__36866),
            .I(N__36820));
    LocalMux I__6852 (
            .O(N__36857),
            .I(N__36820));
    LocalMux I__6851 (
            .O(N__36848),
            .I(N__36820));
    LocalMux I__6850 (
            .O(N__36837),
            .I(N__36820));
    Odrv12 I__6849 (
            .O(N__36820),
            .I(\phase_controller_inst1.stoper_hc.start_latched_i_0 ));
    InMux I__6848 (
            .O(N__36817),
            .I(N__36807));
    InMux I__6847 (
            .O(N__36816),
            .I(N__36807));
    InMux I__6846 (
            .O(N__36815),
            .I(N__36807));
    CascadeMux I__6845 (
            .O(N__36814),
            .I(N__36804));
    LocalMux I__6844 (
            .O(N__36807),
            .I(N__36799));
    InMux I__6843 (
            .O(N__36804),
            .I(N__36794));
    InMux I__6842 (
            .O(N__36803),
            .I(N__36794));
    InMux I__6841 (
            .O(N__36802),
            .I(N__36791));
    Span4Mux_h I__6840 (
            .O(N__36799),
            .I(N__36788));
    LocalMux I__6839 (
            .O(N__36794),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    LocalMux I__6838 (
            .O(N__36791),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    Odrv4 I__6837 (
            .O(N__36788),
            .I(\phase_controller_inst1.stoper_tr.start_latchedZ0 ));
    InMux I__6836 (
            .O(N__36781),
            .I(N__36777));
    CascadeMux I__6835 (
            .O(N__36780),
            .I(N__36773));
    LocalMux I__6834 (
            .O(N__36777),
            .I(N__36767));
    InMux I__6833 (
            .O(N__36776),
            .I(N__36764));
    InMux I__6832 (
            .O(N__36773),
            .I(N__36757));
    InMux I__6831 (
            .O(N__36772),
            .I(N__36757));
    InMux I__6830 (
            .O(N__36771),
            .I(N__36757));
    InMux I__6829 (
            .O(N__36770),
            .I(N__36754));
    Span4Mux_h I__6828 (
            .O(N__36767),
            .I(N__36751));
    LocalMux I__6827 (
            .O(N__36764),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6826 (
            .O(N__36757),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    LocalMux I__6825 (
            .O(N__36754),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    Odrv4 I__6824 (
            .O(N__36751),
            .I(\phase_controller_inst1.start_timer_trZ0 ));
    CascadeMux I__6823 (
            .O(N__36742),
            .I(N__36737));
    InMux I__6822 (
            .O(N__36741),
            .I(N__36734));
    InMux I__6821 (
            .O(N__36740),
            .I(N__36731));
    InMux I__6820 (
            .O(N__36737),
            .I(N__36728));
    LocalMux I__6819 (
            .O(N__36734),
            .I(N__36725));
    LocalMux I__6818 (
            .O(N__36731),
            .I(N__36720));
    LocalMux I__6817 (
            .O(N__36728),
            .I(N__36720));
    Span4Mux_v I__6816 (
            .O(N__36725),
            .I(N__36717));
    Span4Mux_v I__6815 (
            .O(N__36720),
            .I(N__36714));
    Span4Mux_h I__6814 (
            .O(N__36717),
            .I(N__36711));
    Sp12to4 I__6813 (
            .O(N__36714),
            .I(N__36708));
    Odrv4 I__6812 (
            .O(N__36711),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ));
    Odrv12 I__6811 (
            .O(N__36708),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ));
    InMux I__6810 (
            .O(N__36703),
            .I(N__36700));
    LocalMux I__6809 (
            .O(N__36700),
            .I(N__36696));
    InMux I__6808 (
            .O(N__36699),
            .I(N__36693));
    Span4Mux_v I__6807 (
            .O(N__36696),
            .I(N__36687));
    LocalMux I__6806 (
            .O(N__36693),
            .I(N__36684));
    InMux I__6805 (
            .O(N__36692),
            .I(N__36681));
    InMux I__6804 (
            .O(N__36691),
            .I(N__36678));
    InMux I__6803 (
            .O(N__36690),
            .I(N__36674));
    Span4Mux_h I__6802 (
            .O(N__36687),
            .I(N__36669));
    Span4Mux_h I__6801 (
            .O(N__36684),
            .I(N__36669));
    LocalMux I__6800 (
            .O(N__36681),
            .I(N__36666));
    LocalMux I__6799 (
            .O(N__36678),
            .I(N__36663));
    InMux I__6798 (
            .O(N__36677),
            .I(N__36660));
    LocalMux I__6797 (
            .O(N__36674),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__6796 (
            .O(N__36669),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv12 I__6795 (
            .O(N__36666),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    Odrv4 I__6794 (
            .O(N__36663),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    LocalMux I__6793 (
            .O(N__36660),
            .I(elapsed_time_ns_1_RNI0CQBB_0_31));
    InMux I__6792 (
            .O(N__36649),
            .I(N__36646));
    LocalMux I__6791 (
            .O(N__36646),
            .I(N__36643));
    Span4Mux_h I__6790 (
            .O(N__36643),
            .I(N__36640));
    Odrv4 I__6789 (
            .O(N__36640),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ));
    CEMux I__6788 (
            .O(N__36637),
            .I(N__36633));
    CEMux I__6787 (
            .O(N__36636),
            .I(N__36630));
    LocalMux I__6786 (
            .O(N__36633),
            .I(N__36625));
    LocalMux I__6785 (
            .O(N__36630),
            .I(N__36625));
    Span4Mux_v I__6784 (
            .O(N__36625),
            .I(N__36621));
    CEMux I__6783 (
            .O(N__36624),
            .I(N__36618));
    Span4Mux_h I__6782 (
            .O(N__36621),
            .I(N__36611));
    LocalMux I__6781 (
            .O(N__36618),
            .I(N__36611));
    CEMux I__6780 (
            .O(N__36617),
            .I(N__36608));
    CEMux I__6779 (
            .O(N__36616),
            .I(N__36605));
    Span4Mux_h I__6778 (
            .O(N__36611),
            .I(N__36602));
    LocalMux I__6777 (
            .O(N__36608),
            .I(N__36599));
    LocalMux I__6776 (
            .O(N__36605),
            .I(N__36596));
    Sp12to4 I__6775 (
            .O(N__36602),
            .I(N__36588));
    Span12Mux_h I__6774 (
            .O(N__36599),
            .I(N__36588));
    Span4Mux_v I__6773 (
            .O(N__36596),
            .I(N__36585));
    CEMux I__6772 (
            .O(N__36595),
            .I(N__36582));
    CEMux I__6771 (
            .O(N__36594),
            .I(N__36579));
    CEMux I__6770 (
            .O(N__36593),
            .I(N__36576));
    Odrv12 I__6769 (
            .O(N__36588),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__6768 (
            .O(N__36585),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    LocalMux I__6767 (
            .O(N__36582),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    LocalMux I__6766 (
            .O(N__36579),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    LocalMux I__6765 (
            .O(N__36576),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ));
    CEMux I__6764 (
            .O(N__36565),
            .I(N__36561));
    CEMux I__6763 (
            .O(N__36564),
            .I(N__36558));
    LocalMux I__6762 (
            .O(N__36561),
            .I(N__36553));
    LocalMux I__6761 (
            .O(N__36558),
            .I(N__36550));
    CEMux I__6760 (
            .O(N__36557),
            .I(N__36547));
    CEMux I__6759 (
            .O(N__36556),
            .I(N__36544));
    Span4Mux_v I__6758 (
            .O(N__36553),
            .I(N__36541));
    Span4Mux_v I__6757 (
            .O(N__36550),
            .I(N__36538));
    LocalMux I__6756 (
            .O(N__36547),
            .I(N__36535));
    LocalMux I__6755 (
            .O(N__36544),
            .I(N__36532));
    Span4Mux_h I__6754 (
            .O(N__36541),
            .I(N__36529));
    Span4Mux_v I__6753 (
            .O(N__36538),
            .I(N__36526));
    Span4Mux_h I__6752 (
            .O(N__36535),
            .I(N__36523));
    Span4Mux_h I__6751 (
            .O(N__36532),
            .I(N__36520));
    Span4Mux_v I__6750 (
            .O(N__36529),
            .I(N__36515));
    Span4Mux_h I__6749 (
            .O(N__36526),
            .I(N__36515));
    Span4Mux_h I__6748 (
            .O(N__36523),
            .I(N__36512));
    Span4Mux_h I__6747 (
            .O(N__36520),
            .I(N__36509));
    Odrv4 I__6746 (
            .O(N__36515),
            .I(\delay_measurement_inst.delay_tr_timer.N_168_i ));
    Odrv4 I__6745 (
            .O(N__36512),
            .I(\delay_measurement_inst.delay_tr_timer.N_168_i ));
    Odrv4 I__6744 (
            .O(N__36509),
            .I(\delay_measurement_inst.delay_tr_timer.N_168_i ));
    InMux I__6743 (
            .O(N__36502),
            .I(N__36499));
    LocalMux I__6742 (
            .O(N__36499),
            .I(N__36493));
    InMux I__6741 (
            .O(N__36498),
            .I(N__36486));
    InMux I__6740 (
            .O(N__36497),
            .I(N__36486));
    InMux I__6739 (
            .O(N__36496),
            .I(N__36486));
    Span4Mux_h I__6738 (
            .O(N__36493),
            .I(N__36483));
    LocalMux I__6737 (
            .O(N__36486),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    Odrv4 I__6736 (
            .O(N__36483),
            .I(\delay_measurement_inst.delay_tr_timer.runningZ0 ));
    CEMux I__6735 (
            .O(N__36478),
            .I(N__36472));
    CEMux I__6734 (
            .O(N__36477),
            .I(N__36469));
    CEMux I__6733 (
            .O(N__36476),
            .I(N__36466));
    CEMux I__6732 (
            .O(N__36475),
            .I(N__36463));
    LocalMux I__6731 (
            .O(N__36472),
            .I(N__36459));
    LocalMux I__6730 (
            .O(N__36469),
            .I(N__36456));
    LocalMux I__6729 (
            .O(N__36466),
            .I(N__36453));
    LocalMux I__6728 (
            .O(N__36463),
            .I(N__36450));
    CEMux I__6727 (
            .O(N__36462),
            .I(N__36447));
    Span4Mux_v I__6726 (
            .O(N__36459),
            .I(N__36444));
    Span4Mux_h I__6725 (
            .O(N__36456),
            .I(N__36441));
    Span4Mux_v I__6724 (
            .O(N__36453),
            .I(N__36438));
    Span4Mux_v I__6723 (
            .O(N__36450),
            .I(N__36435));
    LocalMux I__6722 (
            .O(N__36447),
            .I(N__36432));
    Span4Mux_h I__6721 (
            .O(N__36444),
            .I(N__36429));
    Span4Mux_h I__6720 (
            .O(N__36441),
            .I(N__36426));
    Span4Mux_h I__6719 (
            .O(N__36438),
            .I(N__36421));
    Span4Mux_h I__6718 (
            .O(N__36435),
            .I(N__36421));
    Span4Mux_h I__6717 (
            .O(N__36432),
            .I(N__36418));
    Odrv4 I__6716 (
            .O(N__36429),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    Odrv4 I__6715 (
            .O(N__36426),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    Odrv4 I__6714 (
            .O(N__36421),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    Odrv4 I__6713 (
            .O(N__36418),
            .I(\delay_measurement_inst.delay_tr_timer.N_167_i ));
    InMux I__6712 (
            .O(N__36409),
            .I(N__36406));
    LocalMux I__6711 (
            .O(N__36406),
            .I(N__36401));
    InMux I__6710 (
            .O(N__36405),
            .I(N__36398));
    InMux I__6709 (
            .O(N__36404),
            .I(N__36395));
    Span4Mux_v I__6708 (
            .O(N__36401),
            .I(N__36388));
    LocalMux I__6707 (
            .O(N__36398),
            .I(N__36388));
    LocalMux I__6706 (
            .O(N__36395),
            .I(N__36388));
    Span4Mux_v I__6705 (
            .O(N__36388),
            .I(N__36385));
    Sp12to4 I__6704 (
            .O(N__36385),
            .I(N__36382));
    Span12Mux_h I__6703 (
            .O(N__36382),
            .I(N__36379));
    Odrv12 I__6702 (
            .O(N__36379),
            .I(il_max_comp1_c));
    InMux I__6701 (
            .O(N__36376),
            .I(N__36371));
    InMux I__6700 (
            .O(N__36375),
            .I(N__36366));
    InMux I__6699 (
            .O(N__36374),
            .I(N__36366));
    LocalMux I__6698 (
            .O(N__36371),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    LocalMux I__6697 (
            .O(N__36366),
            .I(\phase_controller_inst1.stoper_hc.runningZ0 ));
    CascadeMux I__6696 (
            .O(N__36361),
            .I(\phase_controller_inst1.stoper_hc.un4_start_0_cascade_ ));
    InMux I__6695 (
            .O(N__36358),
            .I(N__36346));
    InMux I__6694 (
            .O(N__36357),
            .I(N__36346));
    InMux I__6693 (
            .O(N__36356),
            .I(N__36346));
    InMux I__6692 (
            .O(N__36355),
            .I(N__36339));
    InMux I__6691 (
            .O(N__36354),
            .I(N__36339));
    InMux I__6690 (
            .O(N__36353),
            .I(N__36339));
    LocalMux I__6689 (
            .O(N__36346),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    LocalMux I__6688 (
            .O(N__36339),
            .I(\phase_controller_inst1.start_timer_hcZ0 ));
    InMux I__6687 (
            .O(N__36334),
            .I(N__36329));
    InMux I__6686 (
            .O(N__36333),
            .I(N__36324));
    InMux I__6685 (
            .O(N__36332),
            .I(N__36324));
    LocalMux I__6684 (
            .O(N__36329),
            .I(N__36321));
    LocalMux I__6683 (
            .O(N__36324),
            .I(N__36318));
    Span4Mux_v I__6682 (
            .O(N__36321),
            .I(N__36315));
    Span4Mux_v I__6681 (
            .O(N__36318),
            .I(N__36312));
    Sp12to4 I__6680 (
            .O(N__36315),
            .I(N__36307));
    Sp12to4 I__6679 (
            .O(N__36312),
            .I(N__36307));
    Span12Mux_h I__6678 (
            .O(N__36307),
            .I(N__36304));
    Odrv12 I__6677 (
            .O(N__36304),
            .I(il_min_comp1_c));
    CascadeMux I__6676 (
            .O(N__36301),
            .I(N__36297));
    InMux I__6675 (
            .O(N__36300),
            .I(N__36294));
    InMux I__6674 (
            .O(N__36297),
            .I(N__36289));
    LocalMux I__6673 (
            .O(N__36294),
            .I(N__36286));
    InMux I__6672 (
            .O(N__36293),
            .I(N__36281));
    InMux I__6671 (
            .O(N__36292),
            .I(N__36281));
    LocalMux I__6670 (
            .O(N__36289),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    Odrv4 I__6669 (
            .O(N__36286),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    LocalMux I__6668 (
            .O(N__36281),
            .I(\phase_controller_inst1.stateZ0Z_2 ));
    CascadeMux I__6667 (
            .O(N__36274),
            .I(N__36269));
    InMux I__6666 (
            .O(N__36273),
            .I(N__36265));
    InMux I__6665 (
            .O(N__36272),
            .I(N__36262));
    InMux I__6664 (
            .O(N__36269),
            .I(N__36257));
    InMux I__6663 (
            .O(N__36268),
            .I(N__36257));
    LocalMux I__6662 (
            .O(N__36265),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__6661 (
            .O(N__36262),
            .I(\phase_controller_inst1.hc_time_passed ));
    LocalMux I__6660 (
            .O(N__36257),
            .I(\phase_controller_inst1.hc_time_passed ));
    InMux I__6659 (
            .O(N__36250),
            .I(N__36244));
    InMux I__6658 (
            .O(N__36249),
            .I(N__36244));
    LocalMux I__6657 (
            .O(N__36244),
            .I(elapsed_time_ns_1_RNIV2EN9_0_30));
    InMux I__6656 (
            .O(N__36241),
            .I(N__36238));
    LocalMux I__6655 (
            .O(N__36238),
            .I(elapsed_time_ns_1_RNI03DN9_0_22));
    CascadeMux I__6654 (
            .O(N__36235),
            .I(elapsed_time_ns_1_RNI03DN9_0_22_cascade_));
    InMux I__6653 (
            .O(N__36232),
            .I(N__36229));
    LocalMux I__6652 (
            .O(N__36229),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29));
    CascadeMux I__6651 (
            .O(N__36226),
            .I(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_));
    InMux I__6650 (
            .O(N__36223),
            .I(N__36220));
    LocalMux I__6649 (
            .O(N__36220),
            .I(N__36217));
    Odrv4 I__6648 (
            .O(N__36217),
            .I(\phase_controller_inst1.start_timer_tr_0_sqmuxa ));
    CEMux I__6647 (
            .O(N__36214),
            .I(N__36210));
    CEMux I__6646 (
            .O(N__36213),
            .I(N__36206));
    LocalMux I__6645 (
            .O(N__36210),
            .I(N__36202));
    CEMux I__6644 (
            .O(N__36209),
            .I(N__36199));
    LocalMux I__6643 (
            .O(N__36206),
            .I(N__36196));
    CEMux I__6642 (
            .O(N__36205),
            .I(N__36193));
    Span4Mux_v I__6641 (
            .O(N__36202),
            .I(N__36190));
    LocalMux I__6640 (
            .O(N__36199),
            .I(N__36187));
    Span4Mux_v I__6639 (
            .O(N__36196),
            .I(N__36184));
    LocalMux I__6638 (
            .O(N__36193),
            .I(N__36181));
    Odrv4 I__6637 (
            .O(N__36190),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv12 I__6636 (
            .O(N__36187),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__6635 (
            .O(N__36184),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    Odrv4 I__6634 (
            .O(N__36181),
            .I(\phase_controller_inst1.stoper_hc.un2_start_0 ));
    InMux I__6633 (
            .O(N__36172),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_25 ));
    InMux I__6632 (
            .O(N__36169),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_26 ));
    InMux I__6631 (
            .O(N__36166),
            .I(N__36161));
    InMux I__6630 (
            .O(N__36165),
            .I(N__36156));
    InMux I__6629 (
            .O(N__36164),
            .I(N__36156));
    LocalMux I__6628 (
            .O(N__36161),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ));
    LocalMux I__6627 (
            .O(N__36156),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ));
    InMux I__6626 (
            .O(N__36151),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_27 ));
    InMux I__6625 (
            .O(N__36148),
            .I(N__36143));
    InMux I__6624 (
            .O(N__36147),
            .I(N__36138));
    InMux I__6623 (
            .O(N__36146),
            .I(N__36138));
    LocalMux I__6622 (
            .O(N__36143),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ));
    LocalMux I__6621 (
            .O(N__36138),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ));
    InMux I__6620 (
            .O(N__36133),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_28 ));
    InMux I__6619 (
            .O(N__36130),
            .I(N__36125));
    InMux I__6618 (
            .O(N__36129),
            .I(N__36122));
    InMux I__6617 (
            .O(N__36128),
            .I(N__36119));
    LocalMux I__6616 (
            .O(N__36125),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    LocalMux I__6615 (
            .O(N__36122),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    LocalMux I__6614 (
            .O(N__36119),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ));
    InMux I__6613 (
            .O(N__36112),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_29 ));
    InMux I__6612 (
            .O(N__36109),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_30 ));
    InMux I__6611 (
            .O(N__36106),
            .I(N__36101));
    InMux I__6610 (
            .O(N__36105),
            .I(N__36096));
    InMux I__6609 (
            .O(N__36104),
            .I(N__36096));
    LocalMux I__6608 (
            .O(N__36101),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    LocalMux I__6607 (
            .O(N__36096),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ));
    InMux I__6606 (
            .O(N__36091),
            .I(N__36088));
    LocalMux I__6605 (
            .O(N__36088),
            .I(elapsed_time_ns_1_RNI36DN9_0_25));
    CascadeMux I__6604 (
            .O(N__36085),
            .I(elapsed_time_ns_1_RNI36DN9_0_25_cascade_));
    InMux I__6603 (
            .O(N__36082),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_16 ));
    InMux I__6602 (
            .O(N__36079),
            .I(N__36072));
    InMux I__6601 (
            .O(N__36078),
            .I(N__36072));
    InMux I__6600 (
            .O(N__36077),
            .I(N__36069));
    LocalMux I__6599 (
            .O(N__36072),
            .I(N__36066));
    LocalMux I__6598 (
            .O(N__36069),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ));
    Odrv4 I__6597 (
            .O(N__36066),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ));
    InMux I__6596 (
            .O(N__36061),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_17 ));
    CascadeMux I__6595 (
            .O(N__36058),
            .I(N__36054));
    CascadeMux I__6594 (
            .O(N__36057),
            .I(N__36051));
    InMux I__6593 (
            .O(N__36054),
            .I(N__36046));
    InMux I__6592 (
            .O(N__36051),
            .I(N__36046));
    LocalMux I__6591 (
            .O(N__36046),
            .I(N__36042));
    InMux I__6590 (
            .O(N__36045),
            .I(N__36039));
    Span4Mux_h I__6589 (
            .O(N__36042),
            .I(N__36036));
    LocalMux I__6588 (
            .O(N__36039),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__6587 (
            .O(N__36036),
            .I(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ));
    InMux I__6586 (
            .O(N__36031),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_18 ));
    InMux I__6585 (
            .O(N__36028),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_19 ));
    InMux I__6584 (
            .O(N__36025),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_20 ));
    InMux I__6583 (
            .O(N__36022),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_21 ));
    InMux I__6582 (
            .O(N__36019),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_22 ));
    InMux I__6581 (
            .O(N__36016),
            .I(bfn_13_10_0_));
    InMux I__6580 (
            .O(N__36013),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_24 ));
    InMux I__6579 (
            .O(N__36010),
            .I(bfn_13_8_0_));
    InMux I__6578 (
            .O(N__36007),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_8 ));
    InMux I__6577 (
            .O(N__36004),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_9 ));
    InMux I__6576 (
            .O(N__36001),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_10 ));
    InMux I__6575 (
            .O(N__35998),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_11 ));
    InMux I__6574 (
            .O(N__35995),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_12 ));
    InMux I__6573 (
            .O(N__35992),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_13 ));
    InMux I__6572 (
            .O(N__35989),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_14 ));
    InMux I__6571 (
            .O(N__35986),
            .I(bfn_13_9_0_));
    InMux I__6570 (
            .O(N__35983),
            .I(N__35977));
    InMux I__6569 (
            .O(N__35982),
            .I(N__35977));
    LocalMux I__6568 (
            .O(N__35977),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ));
    InMux I__6567 (
            .O(N__35974),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_0 ));
    InMux I__6566 (
            .O(N__35971),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_1 ));
    InMux I__6565 (
            .O(N__35968),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_2 ));
    InMux I__6564 (
            .O(N__35965),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_3 ));
    InMux I__6563 (
            .O(N__35962),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_4 ));
    InMux I__6562 (
            .O(N__35959),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_5 ));
    InMux I__6561 (
            .O(N__35956),
            .I(\phase_controller_inst1.stoper_hc.counter_cry_6 ));
    CascadeMux I__6560 (
            .O(N__35953),
            .I(N__35949));
    CascadeMux I__6559 (
            .O(N__35952),
            .I(N__35946));
    InMux I__6558 (
            .O(N__35949),
            .I(N__35943));
    InMux I__6557 (
            .O(N__35946),
            .I(N__35939));
    LocalMux I__6556 (
            .O(N__35943),
            .I(N__35936));
    InMux I__6555 (
            .O(N__35942),
            .I(N__35933));
    LocalMux I__6554 (
            .O(N__35939),
            .I(N__35929));
    Span4Mux_v I__6553 (
            .O(N__35936),
            .I(N__35926));
    LocalMux I__6552 (
            .O(N__35933),
            .I(N__35923));
    InMux I__6551 (
            .O(N__35932),
            .I(N__35920));
    Span4Mux_v I__6550 (
            .O(N__35929),
            .I(N__35913));
    Span4Mux_h I__6549 (
            .O(N__35926),
            .I(N__35913));
    Span4Mux_v I__6548 (
            .O(N__35923),
            .I(N__35913));
    LocalMux I__6547 (
            .O(N__35920),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    Odrv4 I__6546 (
            .O(N__35913),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ));
    InMux I__6545 (
            .O(N__35908),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ));
    CascadeMux I__6544 (
            .O(N__35905),
            .I(N__35902));
    InMux I__6543 (
            .O(N__35902),
            .I(N__35899));
    LocalMux I__6542 (
            .O(N__35899),
            .I(N__35894));
    InMux I__6541 (
            .O(N__35898),
            .I(N__35890));
    InMux I__6540 (
            .O(N__35897),
            .I(N__35887));
    Span4Mux_v I__6539 (
            .O(N__35894),
            .I(N__35884));
    InMux I__6538 (
            .O(N__35893),
            .I(N__35881));
    LocalMux I__6537 (
            .O(N__35890),
            .I(N__35876));
    LocalMux I__6536 (
            .O(N__35887),
            .I(N__35876));
    Odrv4 I__6535 (
            .O(N__35884),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    LocalMux I__6534 (
            .O(N__35881),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    Odrv4 I__6533 (
            .O(N__35876),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ));
    InMux I__6532 (
            .O(N__35869),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ));
    InMux I__6531 (
            .O(N__35866),
            .I(N__35852));
    InMux I__6530 (
            .O(N__35865),
            .I(N__35845));
    InMux I__6529 (
            .O(N__35864),
            .I(N__35845));
    InMux I__6528 (
            .O(N__35863),
            .I(N__35845));
    InMux I__6527 (
            .O(N__35862),
            .I(N__35842));
    InMux I__6526 (
            .O(N__35861),
            .I(N__35833));
    InMux I__6525 (
            .O(N__35860),
            .I(N__35833));
    InMux I__6524 (
            .O(N__35859),
            .I(N__35833));
    InMux I__6523 (
            .O(N__35858),
            .I(N__35833));
    InMux I__6522 (
            .O(N__35857),
            .I(N__35830));
    InMux I__6521 (
            .O(N__35856),
            .I(N__35806));
    InMux I__6520 (
            .O(N__35855),
            .I(N__35806));
    LocalMux I__6519 (
            .O(N__35852),
            .I(N__35803));
    LocalMux I__6518 (
            .O(N__35845),
            .I(N__35800));
    LocalMux I__6517 (
            .O(N__35842),
            .I(N__35797));
    LocalMux I__6516 (
            .O(N__35833),
            .I(N__35792));
    LocalMux I__6515 (
            .O(N__35830),
            .I(N__35792));
    InMux I__6514 (
            .O(N__35829),
            .I(N__35789));
    InMux I__6513 (
            .O(N__35828),
            .I(N__35774));
    InMux I__6512 (
            .O(N__35827),
            .I(N__35774));
    InMux I__6511 (
            .O(N__35826),
            .I(N__35774));
    InMux I__6510 (
            .O(N__35825),
            .I(N__35774));
    InMux I__6509 (
            .O(N__35824),
            .I(N__35774));
    InMux I__6508 (
            .O(N__35823),
            .I(N__35774));
    InMux I__6507 (
            .O(N__35822),
            .I(N__35774));
    InMux I__6506 (
            .O(N__35821),
            .I(N__35771));
    InMux I__6505 (
            .O(N__35820),
            .I(N__35762));
    InMux I__6504 (
            .O(N__35819),
            .I(N__35762));
    InMux I__6503 (
            .O(N__35818),
            .I(N__35762));
    InMux I__6502 (
            .O(N__35817),
            .I(N__35762));
    InMux I__6501 (
            .O(N__35816),
            .I(N__35749));
    InMux I__6500 (
            .O(N__35815),
            .I(N__35749));
    InMux I__6499 (
            .O(N__35814),
            .I(N__35749));
    InMux I__6498 (
            .O(N__35813),
            .I(N__35749));
    InMux I__6497 (
            .O(N__35812),
            .I(N__35749));
    InMux I__6496 (
            .O(N__35811),
            .I(N__35749));
    LocalMux I__6495 (
            .O(N__35806),
            .I(N__35744));
    Span4Mux_h I__6494 (
            .O(N__35803),
            .I(N__35744));
    Span4Mux_v I__6493 (
            .O(N__35800),
            .I(N__35737));
    Span4Mux_h I__6492 (
            .O(N__35797),
            .I(N__35737));
    Span4Mux_h I__6491 (
            .O(N__35792),
            .I(N__35737));
    LocalMux I__6490 (
            .O(N__35789),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6489 (
            .O(N__35774),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6488 (
            .O(N__35771),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6487 (
            .O(N__35762),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    LocalMux I__6486 (
            .O(N__35749),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__6485 (
            .O(N__35744),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    Odrv4 I__6484 (
            .O(N__35737),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ));
    InMux I__6483 (
            .O(N__35722),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ));
    IoInMux I__6482 (
            .O(N__35719),
            .I(N__35716));
    LocalMux I__6481 (
            .O(N__35716),
            .I(N__35713));
    Span4Mux_s0_v I__6480 (
            .O(N__35713),
            .I(N__35710));
    Odrv4 I__6479 (
            .O(N__35710),
            .I(GB_BUFFER_reset_c_g_THRU_CO));
    InMux I__6478 (
            .O(N__35707),
            .I(N__35701));
    InMux I__6477 (
            .O(N__35706),
            .I(N__35701));
    LocalMux I__6476 (
            .O(N__35701),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ));
    InMux I__6475 (
            .O(N__35698),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ));
    CascadeMux I__6474 (
            .O(N__35695),
            .I(N__35692));
    InMux I__6473 (
            .O(N__35692),
            .I(N__35689));
    LocalMux I__6472 (
            .O(N__35689),
            .I(N__35686));
    Span4Mux_h I__6471 (
            .O(N__35686),
            .I(N__35680));
    InMux I__6470 (
            .O(N__35685),
            .I(N__35677));
    InMux I__6469 (
            .O(N__35684),
            .I(N__35672));
    InMux I__6468 (
            .O(N__35683),
            .I(N__35672));
    Odrv4 I__6467 (
            .O(N__35680),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__6466 (
            .O(N__35677),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    LocalMux I__6465 (
            .O(N__35672),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ));
    InMux I__6464 (
            .O(N__35665),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ));
    InMux I__6463 (
            .O(N__35662),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ));
    CascadeMux I__6462 (
            .O(N__35659),
            .I(N__35656));
    InMux I__6461 (
            .O(N__35656),
            .I(N__35653));
    LocalMux I__6460 (
            .O(N__35653),
            .I(N__35649));
    InMux I__6459 (
            .O(N__35652),
            .I(N__35646));
    Span4Mux_v I__6458 (
            .O(N__35649),
            .I(N__35639));
    LocalMux I__6457 (
            .O(N__35646),
            .I(N__35639));
    InMux I__6456 (
            .O(N__35645),
            .I(N__35636));
    InMux I__6455 (
            .O(N__35644),
            .I(N__35633));
    Odrv4 I__6454 (
            .O(N__35639),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__6453 (
            .O(N__35636),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    LocalMux I__6452 (
            .O(N__35633),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ));
    InMux I__6451 (
            .O(N__35626),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ));
    CascadeMux I__6450 (
            .O(N__35623),
            .I(N__35620));
    InMux I__6449 (
            .O(N__35620),
            .I(N__35617));
    LocalMux I__6448 (
            .O(N__35617),
            .I(N__35613));
    CascadeMux I__6447 (
            .O(N__35616),
            .I(N__35608));
    Span4Mux_h I__6446 (
            .O(N__35613),
            .I(N__35605));
    InMux I__6445 (
            .O(N__35612),
            .I(N__35602));
    InMux I__6444 (
            .O(N__35611),
            .I(N__35597));
    InMux I__6443 (
            .O(N__35608),
            .I(N__35597));
    Odrv4 I__6442 (
            .O(N__35605),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__6441 (
            .O(N__35602),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    LocalMux I__6440 (
            .O(N__35597),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ));
    InMux I__6439 (
            .O(N__35590),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ));
    CascadeMux I__6438 (
            .O(N__35587),
            .I(N__35584));
    InMux I__6437 (
            .O(N__35584),
            .I(N__35581));
    LocalMux I__6436 (
            .O(N__35581),
            .I(N__35578));
    Span4Mux_h I__6435 (
            .O(N__35578),
            .I(N__35572));
    InMux I__6434 (
            .O(N__35577),
            .I(N__35569));
    InMux I__6433 (
            .O(N__35576),
            .I(N__35564));
    InMux I__6432 (
            .O(N__35575),
            .I(N__35564));
    Odrv4 I__6431 (
            .O(N__35572),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__6430 (
            .O(N__35569),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    LocalMux I__6429 (
            .O(N__35564),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ));
    InMux I__6428 (
            .O(N__35557),
            .I(bfn_12_23_0_));
    CascadeMux I__6427 (
            .O(N__35554),
            .I(N__35551));
    InMux I__6426 (
            .O(N__35551),
            .I(N__35548));
    LocalMux I__6425 (
            .O(N__35548),
            .I(N__35543));
    InMux I__6424 (
            .O(N__35547),
            .I(N__35540));
    CascadeMux I__6423 (
            .O(N__35546),
            .I(N__35537));
    Span4Mux_v I__6422 (
            .O(N__35543),
            .I(N__35531));
    LocalMux I__6421 (
            .O(N__35540),
            .I(N__35531));
    InMux I__6420 (
            .O(N__35537),
            .I(N__35526));
    InMux I__6419 (
            .O(N__35536),
            .I(N__35526));
    Odrv4 I__6418 (
            .O(N__35531),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    LocalMux I__6417 (
            .O(N__35526),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ));
    InMux I__6416 (
            .O(N__35521),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ));
    CascadeMux I__6415 (
            .O(N__35518),
            .I(N__35515));
    InMux I__6414 (
            .O(N__35515),
            .I(N__35511));
    InMux I__6413 (
            .O(N__35514),
            .I(N__35508));
    LocalMux I__6412 (
            .O(N__35511),
            .I(N__35505));
    LocalMux I__6411 (
            .O(N__35508),
            .I(N__35500));
    Span4Mux_h I__6410 (
            .O(N__35505),
            .I(N__35497));
    InMux I__6409 (
            .O(N__35504),
            .I(N__35494));
    InMux I__6408 (
            .O(N__35503),
            .I(N__35491));
    Span4Mux_v I__6407 (
            .O(N__35500),
            .I(N__35488));
    Odrv4 I__6406 (
            .O(N__35497),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__6405 (
            .O(N__35494),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    LocalMux I__6404 (
            .O(N__35491),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    Odrv4 I__6403 (
            .O(N__35488),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ));
    InMux I__6402 (
            .O(N__35479),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ));
    CascadeMux I__6401 (
            .O(N__35476),
            .I(N__35473));
    InMux I__6400 (
            .O(N__35473),
            .I(N__35469));
    InMux I__6399 (
            .O(N__35472),
            .I(N__35466));
    LocalMux I__6398 (
            .O(N__35469),
            .I(N__35463));
    LocalMux I__6397 (
            .O(N__35466),
            .I(N__35458));
    Span4Mux_h I__6396 (
            .O(N__35463),
            .I(N__35455));
    InMux I__6395 (
            .O(N__35462),
            .I(N__35452));
    InMux I__6394 (
            .O(N__35461),
            .I(N__35449));
    Span4Mux_v I__6393 (
            .O(N__35458),
            .I(N__35446));
    Odrv4 I__6392 (
            .O(N__35455),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__6391 (
            .O(N__35452),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    LocalMux I__6390 (
            .O(N__35449),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    Odrv4 I__6389 (
            .O(N__35446),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ));
    InMux I__6388 (
            .O(N__35437),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ));
    InMux I__6387 (
            .O(N__35434),
            .I(N__35431));
    LocalMux I__6386 (
            .O(N__35431),
            .I(N__35428));
    Odrv4 I__6385 (
            .O(N__35428),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ));
    CascadeMux I__6384 (
            .O(N__35425),
            .I(N__35420));
    InMux I__6383 (
            .O(N__35424),
            .I(N__35417));
    CascadeMux I__6382 (
            .O(N__35423),
            .I(N__35414));
    InMux I__6381 (
            .O(N__35420),
            .I(N__35410));
    LocalMux I__6380 (
            .O(N__35417),
            .I(N__35407));
    InMux I__6379 (
            .O(N__35414),
            .I(N__35404));
    CascadeMux I__6378 (
            .O(N__35413),
            .I(N__35401));
    LocalMux I__6377 (
            .O(N__35410),
            .I(N__35394));
    Span4Mux_v I__6376 (
            .O(N__35407),
            .I(N__35394));
    LocalMux I__6375 (
            .O(N__35404),
            .I(N__35394));
    InMux I__6374 (
            .O(N__35401),
            .I(N__35391));
    Span4Mux_h I__6373 (
            .O(N__35394),
            .I(N__35388));
    LocalMux I__6372 (
            .O(N__35391),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    Odrv4 I__6371 (
            .O(N__35388),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ));
    InMux I__6370 (
            .O(N__35383),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ));
    InMux I__6369 (
            .O(N__35380),
            .I(N__35377));
    LocalMux I__6368 (
            .O(N__35377),
            .I(N__35374));
    Odrv12 I__6367 (
            .O(N__35374),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ));
    CascadeMux I__6366 (
            .O(N__35371),
            .I(N__35367));
    CascadeMux I__6365 (
            .O(N__35370),
            .I(N__35364));
    InMux I__6364 (
            .O(N__35367),
            .I(N__35359));
    InMux I__6363 (
            .O(N__35364),
            .I(N__35356));
    InMux I__6362 (
            .O(N__35363),
            .I(N__35353));
    InMux I__6361 (
            .O(N__35362),
            .I(N__35350));
    LocalMux I__6360 (
            .O(N__35359),
            .I(N__35345));
    LocalMux I__6359 (
            .O(N__35356),
            .I(N__35345));
    LocalMux I__6358 (
            .O(N__35353),
            .I(N__35342));
    LocalMux I__6357 (
            .O(N__35350),
            .I(N__35339));
    Span4Mux_h I__6356 (
            .O(N__35345),
            .I(N__35336));
    Span4Mux_h I__6355 (
            .O(N__35342),
            .I(N__35331));
    Span4Mux_h I__6354 (
            .O(N__35339),
            .I(N__35331));
    Odrv4 I__6353 (
            .O(N__35336),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    Odrv4 I__6352 (
            .O(N__35331),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ));
    InMux I__6351 (
            .O(N__35326),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ));
    InMux I__6350 (
            .O(N__35323),
            .I(N__35320));
    LocalMux I__6349 (
            .O(N__35320),
            .I(N__35317));
    Odrv4 I__6348 (
            .O(N__35317),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ));
    CascadeMux I__6347 (
            .O(N__35314),
            .I(N__35311));
    InMux I__6346 (
            .O(N__35311),
            .I(N__35308));
    LocalMux I__6345 (
            .O(N__35308),
            .I(N__35304));
    CascadeMux I__6344 (
            .O(N__35307),
            .I(N__35301));
    Span4Mux_v I__6343 (
            .O(N__35304),
            .I(N__35296));
    InMux I__6342 (
            .O(N__35301),
            .I(N__35293));
    InMux I__6341 (
            .O(N__35300),
            .I(N__35290));
    InMux I__6340 (
            .O(N__35299),
            .I(N__35287));
    Odrv4 I__6339 (
            .O(N__35296),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__6338 (
            .O(N__35293),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__6337 (
            .O(N__35290),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    LocalMux I__6336 (
            .O(N__35287),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ));
    InMux I__6335 (
            .O(N__35278),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ));
    InMux I__6334 (
            .O(N__35275),
            .I(N__35272));
    LocalMux I__6333 (
            .O(N__35272),
            .I(N__35269));
    Odrv4 I__6332 (
            .O(N__35269),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ));
    CascadeMux I__6331 (
            .O(N__35266),
            .I(N__35262));
    InMux I__6330 (
            .O(N__35265),
            .I(N__35257));
    InMux I__6329 (
            .O(N__35262),
            .I(N__35254));
    InMux I__6328 (
            .O(N__35261),
            .I(N__35251));
    InMux I__6327 (
            .O(N__35260),
            .I(N__35248));
    LocalMux I__6326 (
            .O(N__35257),
            .I(N__35245));
    LocalMux I__6325 (
            .O(N__35254),
            .I(N__35240));
    LocalMux I__6324 (
            .O(N__35251),
            .I(N__35240));
    LocalMux I__6323 (
            .O(N__35248),
            .I(N__35237));
    Span4Mux_v I__6322 (
            .O(N__35245),
            .I(N__35232));
    Span4Mux_h I__6321 (
            .O(N__35240),
            .I(N__35232));
    Span4Mux_h I__6320 (
            .O(N__35237),
            .I(N__35229));
    Odrv4 I__6319 (
            .O(N__35232),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    Odrv4 I__6318 (
            .O(N__35229),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ));
    InMux I__6317 (
            .O(N__35224),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ));
    InMux I__6316 (
            .O(N__35221),
            .I(N__35218));
    LocalMux I__6315 (
            .O(N__35218),
            .I(N__35215));
    Odrv4 I__6314 (
            .O(N__35215),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ));
    CascadeMux I__6313 (
            .O(N__35212),
            .I(N__35209));
    InMux I__6312 (
            .O(N__35209),
            .I(N__35206));
    LocalMux I__6311 (
            .O(N__35206),
            .I(N__35203));
    Span4Mux_h I__6310 (
            .O(N__35203),
            .I(N__35197));
    InMux I__6309 (
            .O(N__35202),
            .I(N__35194));
    InMux I__6308 (
            .O(N__35201),
            .I(N__35191));
    InMux I__6307 (
            .O(N__35200),
            .I(N__35188));
    Odrv4 I__6306 (
            .O(N__35197),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__6305 (
            .O(N__35194),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__6304 (
            .O(N__35191),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    LocalMux I__6303 (
            .O(N__35188),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ));
    InMux I__6302 (
            .O(N__35179),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ));
    InMux I__6301 (
            .O(N__35176),
            .I(N__35173));
    LocalMux I__6300 (
            .O(N__35173),
            .I(N__35170));
    Odrv4 I__6299 (
            .O(N__35170),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ));
    InMux I__6298 (
            .O(N__35167),
            .I(bfn_12_22_0_));
    CascadeMux I__6297 (
            .O(N__35164),
            .I(N__35161));
    InMux I__6296 (
            .O(N__35161),
            .I(N__35158));
    LocalMux I__6295 (
            .O(N__35158),
            .I(N__35154));
    CascadeMux I__6294 (
            .O(N__35157),
            .I(N__35151));
    Span4Mux_h I__6293 (
            .O(N__35154),
            .I(N__35146));
    InMux I__6292 (
            .O(N__35151),
            .I(N__35143));
    InMux I__6291 (
            .O(N__35150),
            .I(N__35140));
    InMux I__6290 (
            .O(N__35149),
            .I(N__35137));
    Odrv4 I__6289 (
            .O(N__35146),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__6288 (
            .O(N__35143),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__6287 (
            .O(N__35140),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    LocalMux I__6286 (
            .O(N__35137),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ));
    InMux I__6285 (
            .O(N__35128),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ));
    InMux I__6284 (
            .O(N__35125),
            .I(N__35122));
    LocalMux I__6283 (
            .O(N__35122),
            .I(N__35119));
    Span4Mux_v I__6282 (
            .O(N__35119),
            .I(N__35116));
    Odrv4 I__6281 (
            .O(N__35116),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ));
    InMux I__6280 (
            .O(N__35113),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ));
    InMux I__6279 (
            .O(N__35110),
            .I(N__35107));
    LocalMux I__6278 (
            .O(N__35107),
            .I(N__35104));
    Odrv4 I__6277 (
            .O(N__35104),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ));
    CascadeMux I__6276 (
            .O(N__35101),
            .I(N__35098));
    InMux I__6275 (
            .O(N__35098),
            .I(N__35095));
    LocalMux I__6274 (
            .O(N__35095),
            .I(N__35091));
    InMux I__6273 (
            .O(N__35094),
            .I(N__35086));
    Span4Mux_h I__6272 (
            .O(N__35091),
            .I(N__35083));
    InMux I__6271 (
            .O(N__35090),
            .I(N__35080));
    InMux I__6270 (
            .O(N__35089),
            .I(N__35077));
    LocalMux I__6269 (
            .O(N__35086),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    Odrv4 I__6268 (
            .O(N__35083),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__6267 (
            .O(N__35080),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    LocalMux I__6266 (
            .O(N__35077),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ));
    InMux I__6265 (
            .O(N__35068),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ));
    InMux I__6264 (
            .O(N__35065),
            .I(N__35062));
    LocalMux I__6263 (
            .O(N__35062),
            .I(N__35059));
    Odrv12 I__6262 (
            .O(N__35059),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ));
    CascadeMux I__6261 (
            .O(N__35056),
            .I(N__35053));
    InMux I__6260 (
            .O(N__35053),
            .I(N__35048));
    InMux I__6259 (
            .O(N__35052),
            .I(N__35045));
    CascadeMux I__6258 (
            .O(N__35051),
            .I(N__35042));
    LocalMux I__6257 (
            .O(N__35048),
            .I(N__35038));
    LocalMux I__6256 (
            .O(N__35045),
            .I(N__35035));
    InMux I__6255 (
            .O(N__35042),
            .I(N__35032));
    InMux I__6254 (
            .O(N__35041),
            .I(N__35029));
    Span4Mux_h I__6253 (
            .O(N__35038),
            .I(N__35026));
    Span4Mux_h I__6252 (
            .O(N__35035),
            .I(N__35023));
    LocalMux I__6251 (
            .O(N__35032),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    LocalMux I__6250 (
            .O(N__35029),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__6249 (
            .O(N__35026),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    Odrv4 I__6248 (
            .O(N__35023),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ));
    InMux I__6247 (
            .O(N__35014),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ));
    InMux I__6246 (
            .O(N__35011),
            .I(N__35008));
    LocalMux I__6245 (
            .O(N__35008),
            .I(N__35005));
    Odrv4 I__6244 (
            .O(N__35005),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ));
    CascadeMux I__6243 (
            .O(N__35002),
            .I(N__34999));
    InMux I__6242 (
            .O(N__34999),
            .I(N__34994));
    InMux I__6241 (
            .O(N__34998),
            .I(N__34991));
    InMux I__6240 (
            .O(N__34997),
            .I(N__34987));
    LocalMux I__6239 (
            .O(N__34994),
            .I(N__34984));
    LocalMux I__6238 (
            .O(N__34991),
            .I(N__34981));
    InMux I__6237 (
            .O(N__34990),
            .I(N__34978));
    LocalMux I__6236 (
            .O(N__34987),
            .I(N__34971));
    Span4Mux_v I__6235 (
            .O(N__34984),
            .I(N__34971));
    Span4Mux_v I__6234 (
            .O(N__34981),
            .I(N__34971));
    LocalMux I__6233 (
            .O(N__34978),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    Odrv4 I__6232 (
            .O(N__34971),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ));
    InMux I__6231 (
            .O(N__34966),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ));
    InMux I__6230 (
            .O(N__34963),
            .I(N__34960));
    LocalMux I__6229 (
            .O(N__34960),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ));
    CascadeMux I__6228 (
            .O(N__34957),
            .I(N__34954));
    InMux I__6227 (
            .O(N__34954),
            .I(N__34951));
    LocalMux I__6226 (
            .O(N__34951),
            .I(N__34947));
    InMux I__6225 (
            .O(N__34950),
            .I(N__34942));
    Span4Mux_h I__6224 (
            .O(N__34947),
            .I(N__34939));
    InMux I__6223 (
            .O(N__34946),
            .I(N__34936));
    InMux I__6222 (
            .O(N__34945),
            .I(N__34933));
    LocalMux I__6221 (
            .O(N__34942),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    Odrv4 I__6220 (
            .O(N__34939),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__6219 (
            .O(N__34936),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    LocalMux I__6218 (
            .O(N__34933),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ));
    InMux I__6217 (
            .O(N__34924),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ));
    InMux I__6216 (
            .O(N__34921),
            .I(N__34917));
    CascadeMux I__6215 (
            .O(N__34920),
            .I(N__34914));
    LocalMux I__6214 (
            .O(N__34917),
            .I(N__34910));
    InMux I__6213 (
            .O(N__34914),
            .I(N__34906));
    InMux I__6212 (
            .O(N__34913),
            .I(N__34903));
    Span4Mux_v I__6211 (
            .O(N__34910),
            .I(N__34900));
    InMux I__6210 (
            .O(N__34909),
            .I(N__34897));
    LocalMux I__6209 (
            .O(N__34906),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__6208 (
            .O(N__34903),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    Odrv4 I__6207 (
            .O(N__34900),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    LocalMux I__6206 (
            .O(N__34897),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ));
    CascadeMux I__6205 (
            .O(N__34888),
            .I(N__34885));
    InMux I__6204 (
            .O(N__34885),
            .I(N__34882));
    LocalMux I__6203 (
            .O(N__34882),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ));
    InMux I__6202 (
            .O(N__34879),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ));
    InMux I__6201 (
            .O(N__34876),
            .I(N__34873));
    LocalMux I__6200 (
            .O(N__34873),
            .I(N__34870));
    Odrv4 I__6199 (
            .O(N__34870),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ));
    CascadeMux I__6198 (
            .O(N__34867),
            .I(N__34864));
    InMux I__6197 (
            .O(N__34864),
            .I(N__34861));
    LocalMux I__6196 (
            .O(N__34861),
            .I(N__34856));
    CascadeMux I__6195 (
            .O(N__34860),
            .I(N__34852));
    InMux I__6194 (
            .O(N__34859),
            .I(N__34849));
    Span4Mux_h I__6193 (
            .O(N__34856),
            .I(N__34846));
    InMux I__6192 (
            .O(N__34855),
            .I(N__34843));
    InMux I__6191 (
            .O(N__34852),
            .I(N__34840));
    LocalMux I__6190 (
            .O(N__34849),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    Odrv4 I__6189 (
            .O(N__34846),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__6188 (
            .O(N__34843),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    LocalMux I__6187 (
            .O(N__34840),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ));
    InMux I__6186 (
            .O(N__34831),
            .I(bfn_12_21_0_));
    InMux I__6185 (
            .O(N__34828),
            .I(N__34825));
    LocalMux I__6184 (
            .O(N__34825),
            .I(N__34819));
    InMux I__6183 (
            .O(N__34824),
            .I(N__34816));
    InMux I__6182 (
            .O(N__34823),
            .I(N__34813));
    InMux I__6181 (
            .O(N__34822),
            .I(N__34810));
    Span4Mux_h I__6180 (
            .O(N__34819),
            .I(N__34803));
    LocalMux I__6179 (
            .O(N__34816),
            .I(N__34803));
    LocalMux I__6178 (
            .O(N__34813),
            .I(N__34803));
    LocalMux I__6177 (
            .O(N__34810),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    Odrv4 I__6176 (
            .O(N__34803),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ));
    CascadeMux I__6175 (
            .O(N__34798),
            .I(N__34795));
    InMux I__6174 (
            .O(N__34795),
            .I(N__34792));
    LocalMux I__6173 (
            .O(N__34792),
            .I(N__34789));
    Odrv12 I__6172 (
            .O(N__34789),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ));
    InMux I__6171 (
            .O(N__34786),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ));
    InMux I__6170 (
            .O(N__34783),
            .I(N__34780));
    LocalMux I__6169 (
            .O(N__34780),
            .I(N__34777));
    Odrv4 I__6168 (
            .O(N__34777),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ));
    CascadeMux I__6167 (
            .O(N__34774),
            .I(N__34771));
    InMux I__6166 (
            .O(N__34771),
            .I(N__34767));
    InMux I__6165 (
            .O(N__34770),
            .I(N__34763));
    LocalMux I__6164 (
            .O(N__34767),
            .I(N__34760));
    InMux I__6163 (
            .O(N__34766),
            .I(N__34756));
    LocalMux I__6162 (
            .O(N__34763),
            .I(N__34753));
    Span4Mux_h I__6161 (
            .O(N__34760),
            .I(N__34750));
    InMux I__6160 (
            .O(N__34759),
            .I(N__34747));
    LocalMux I__6159 (
            .O(N__34756),
            .I(N__34744));
    Span4Mux_h I__6158 (
            .O(N__34753),
            .I(N__34741));
    Odrv4 I__6157 (
            .O(N__34750),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    LocalMux I__6156 (
            .O(N__34747),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__6155 (
            .O(N__34744),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    Odrv4 I__6154 (
            .O(N__34741),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ));
    InMux I__6153 (
            .O(N__34732),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ));
    InMux I__6152 (
            .O(N__34729),
            .I(N__34726));
    LocalMux I__6151 (
            .O(N__34726),
            .I(N__34722));
    InMux I__6150 (
            .O(N__34725),
            .I(N__34719));
    Span4Mux_h I__6149 (
            .O(N__34722),
            .I(N__34716));
    LocalMux I__6148 (
            .O(N__34719),
            .I(N__34713));
    Odrv4 I__6147 (
            .O(N__34716),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    Odrv4 I__6146 (
            .O(N__34713),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ));
    CascadeMux I__6145 (
            .O(N__34708),
            .I(N__34705));
    InMux I__6144 (
            .O(N__34705),
            .I(N__34702));
    LocalMux I__6143 (
            .O(N__34702),
            .I(N__34698));
    CascadeMux I__6142 (
            .O(N__34701),
            .I(N__34694));
    Span4Mux_h I__6141 (
            .O(N__34698),
            .I(N__34690));
    InMux I__6140 (
            .O(N__34697),
            .I(N__34685));
    InMux I__6139 (
            .O(N__34694),
            .I(N__34685));
    InMux I__6138 (
            .O(N__34693),
            .I(N__34682));
    Odrv4 I__6137 (
            .O(N__34690),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__6136 (
            .O(N__34685),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    LocalMux I__6135 (
            .O(N__34682),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ));
    InMux I__6134 (
            .O(N__34675),
            .I(N__34672));
    LocalMux I__6133 (
            .O(N__34672),
            .I(N__34669));
    Odrv4 I__6132 (
            .O(N__34669),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ));
    CascadeMux I__6131 (
            .O(N__34666),
            .I(N__34663));
    InMux I__6130 (
            .O(N__34663),
            .I(N__34660));
    LocalMux I__6129 (
            .O(N__34660),
            .I(N__34657));
    Span4Mux_h I__6128 (
            .O(N__34657),
            .I(N__34652));
    InMux I__6127 (
            .O(N__34656),
            .I(N__34649));
    InMux I__6126 (
            .O(N__34655),
            .I(N__34646));
    Odrv4 I__6125 (
            .O(N__34652),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__6124 (
            .O(N__34649),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    LocalMux I__6123 (
            .O(N__34646),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ));
    InMux I__6122 (
            .O(N__34639),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ));
    InMux I__6121 (
            .O(N__34636),
            .I(N__34633));
    LocalMux I__6120 (
            .O(N__34633),
            .I(N__34630));
    Span4Mux_v I__6119 (
            .O(N__34630),
            .I(N__34624));
    InMux I__6118 (
            .O(N__34629),
            .I(N__34621));
    InMux I__6117 (
            .O(N__34628),
            .I(N__34618));
    InMux I__6116 (
            .O(N__34627),
            .I(N__34615));
    Odrv4 I__6115 (
            .O(N__34624),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__6114 (
            .O(N__34621),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__6113 (
            .O(N__34618),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    LocalMux I__6112 (
            .O(N__34615),
            .I(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ));
    CascadeMux I__6111 (
            .O(N__34606),
            .I(N__34603));
    InMux I__6110 (
            .O(N__34603),
            .I(N__34600));
    LocalMux I__6109 (
            .O(N__34600),
            .I(N__34597));
    Odrv4 I__6108 (
            .O(N__34597),
            .I(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ));
    InMux I__6107 (
            .O(N__34594),
            .I(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ));
    InMux I__6106 (
            .O(N__34591),
            .I(N__34588));
    LocalMux I__6105 (
            .O(N__34588),
            .I(N__34585));
    Odrv4 I__6104 (
            .O(N__34585),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt28 ));
    InMux I__6103 (
            .O(N__34582),
            .I(N__34578));
    InMux I__6102 (
            .O(N__34581),
            .I(N__34575));
    LocalMux I__6101 (
            .O(N__34578),
            .I(N__34572));
    LocalMux I__6100 (
            .O(N__34575),
            .I(N__34569));
    Span4Mux_v I__6099 (
            .O(N__34572),
            .I(N__34566));
    Span4Mux_h I__6098 (
            .O(N__34569),
            .I(N__34563));
    Odrv4 I__6097 (
            .O(N__34566),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_28));
    Odrv4 I__6096 (
            .O(N__34563),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_28));
    InMux I__6095 (
            .O(N__34558),
            .I(N__34553));
    InMux I__6094 (
            .O(N__34557),
            .I(N__34548));
    InMux I__6093 (
            .O(N__34556),
            .I(N__34548));
    LocalMux I__6092 (
            .O(N__34553),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    LocalMux I__6091 (
            .O(N__34548),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ));
    InMux I__6090 (
            .O(N__34543),
            .I(N__34538));
    InMux I__6089 (
            .O(N__34542),
            .I(N__34533));
    InMux I__6088 (
            .O(N__34541),
            .I(N__34533));
    LocalMux I__6087 (
            .O(N__34538),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ));
    LocalMux I__6086 (
            .O(N__34533),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ));
    CascadeMux I__6085 (
            .O(N__34528),
            .I(N__34525));
    InMux I__6084 (
            .O(N__34525),
            .I(N__34522));
    LocalMux I__6083 (
            .O(N__34522),
            .I(N__34519));
    Odrv4 I__6082 (
            .O(N__34519),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ));
    CascadeMux I__6081 (
            .O(N__34516),
            .I(N__34513));
    InMux I__6080 (
            .O(N__34513),
            .I(N__34510));
    LocalMux I__6079 (
            .O(N__34510),
            .I(N__34507));
    Odrv12 I__6078 (
            .O(N__34507),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ));
    InMux I__6077 (
            .O(N__34504),
            .I(N__34499));
    InMux I__6076 (
            .O(N__34503),
            .I(N__34494));
    InMux I__6075 (
            .O(N__34502),
            .I(N__34494));
    LocalMux I__6074 (
            .O(N__34499),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    LocalMux I__6073 (
            .O(N__34494),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ));
    CascadeMux I__6072 (
            .O(N__34489),
            .I(N__34486));
    InMux I__6071 (
            .O(N__34486),
            .I(N__34474));
    InMux I__6070 (
            .O(N__34485),
            .I(N__34474));
    InMux I__6069 (
            .O(N__34484),
            .I(N__34474));
    InMux I__6068 (
            .O(N__34483),
            .I(N__34474));
    LocalMux I__6067 (
            .O(N__34474),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ));
    InMux I__6066 (
            .O(N__34471),
            .I(N__34466));
    InMux I__6065 (
            .O(N__34470),
            .I(N__34461));
    InMux I__6064 (
            .O(N__34469),
            .I(N__34461));
    LocalMux I__6063 (
            .O(N__34466),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    LocalMux I__6062 (
            .O(N__34461),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ));
    InMux I__6061 (
            .O(N__34456),
            .I(N__34453));
    LocalMux I__6060 (
            .O(N__34453),
            .I(N__34450));
    Odrv4 I__6059 (
            .O(N__34450),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt30 ));
    InMux I__6058 (
            .O(N__34447),
            .I(N__34444));
    LocalMux I__6057 (
            .O(N__34444),
            .I(N__34441));
    Span4Mux_v I__6056 (
            .O(N__34441),
            .I(N__34437));
    InMux I__6055 (
            .O(N__34440),
            .I(N__34431));
    Span4Mux_v I__6054 (
            .O(N__34437),
            .I(N__34427));
    InMux I__6053 (
            .O(N__34436),
            .I(N__34422));
    InMux I__6052 (
            .O(N__34435),
            .I(N__34422));
    InMux I__6051 (
            .O(N__34434),
            .I(N__34419));
    LocalMux I__6050 (
            .O(N__34431),
            .I(N__34416));
    InMux I__6049 (
            .O(N__34430),
            .I(N__34413));
    Span4Mux_h I__6048 (
            .O(N__34427),
            .I(N__34410));
    LocalMux I__6047 (
            .O(N__34422),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__6046 (
            .O(N__34419),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__6045 (
            .O(N__34416),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    LocalMux I__6044 (
            .O(N__34413),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    Odrv4 I__6043 (
            .O(N__34410),
            .I(\phase_controller_inst2.start_timer_hcZ0 ));
    InMux I__6042 (
            .O(N__34399),
            .I(N__34392));
    InMux I__6041 (
            .O(N__34398),
            .I(N__34387));
    InMux I__6040 (
            .O(N__34397),
            .I(N__34387));
    CascadeMux I__6039 (
            .O(N__34396),
            .I(N__34383));
    InMux I__6038 (
            .O(N__34395),
            .I(N__34380));
    LocalMux I__6037 (
            .O(N__34392),
            .I(N__34377));
    LocalMux I__6036 (
            .O(N__34387),
            .I(N__34374));
    InMux I__6035 (
            .O(N__34386),
            .I(N__34371));
    InMux I__6034 (
            .O(N__34383),
            .I(N__34368));
    LocalMux I__6033 (
            .O(N__34380),
            .I(N__34363));
    Span12Mux_h I__6032 (
            .O(N__34377),
            .I(N__34363));
    Span4Mux_h I__6031 (
            .O(N__34374),
            .I(N__34360));
    LocalMux I__6030 (
            .O(N__34371),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    LocalMux I__6029 (
            .O(N__34368),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv12 I__6028 (
            .O(N__34363),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    Odrv4 I__6027 (
            .O(N__34360),
            .I(\phase_controller_inst2.stoper_hc.start_latchedZ0 ));
    InMux I__6026 (
            .O(N__34351),
            .I(N__34348));
    LocalMux I__6025 (
            .O(N__34348),
            .I(N__34345));
    Sp12to4 I__6024 (
            .O(N__34345),
            .I(N__34342));
    Span12Mux_v I__6023 (
            .O(N__34342),
            .I(N__34339));
    Odrv12 I__6022 (
            .O(N__34339),
            .I(\phase_controller_inst2.stoper_hc.un4_start_0 ));
    InMux I__6021 (
            .O(N__34336),
            .I(N__34330));
    InMux I__6020 (
            .O(N__34335),
            .I(N__34330));
    LocalMux I__6019 (
            .O(N__34330),
            .I(N__34327));
    Span4Mux_h I__6018 (
            .O(N__34327),
            .I(N__34323));
    InMux I__6017 (
            .O(N__34326),
            .I(N__34320));
    Odrv4 I__6016 (
            .O(N__34323),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ));
    LocalMux I__6015 (
            .O(N__34320),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ));
    InMux I__6014 (
            .O(N__34315),
            .I(N__34312));
    LocalMux I__6013 (
            .O(N__34312),
            .I(N__34307));
    InMux I__6012 (
            .O(N__34311),
            .I(N__34304));
    InMux I__6011 (
            .O(N__34310),
            .I(N__34301));
    Span4Mux_h I__6010 (
            .O(N__34307),
            .I(N__34298));
    LocalMux I__6009 (
            .O(N__34304),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    LocalMux I__6008 (
            .O(N__34301),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    Odrv4 I__6007 (
            .O(N__34298),
            .I(\phase_controller_inst1.stoper_tr.runningZ0 ));
    InMux I__6006 (
            .O(N__34291),
            .I(N__34288));
    LocalMux I__6005 (
            .O(N__34288),
            .I(N__34285));
    Span4Mux_h I__6004 (
            .O(N__34285),
            .I(N__34282));
    Span4Mux_h I__6003 (
            .O(N__34282),
            .I(N__34278));
    InMux I__6002 (
            .O(N__34281),
            .I(N__34275));
    Odrv4 I__6001 (
            .O(N__34278),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_14));
    LocalMux I__6000 (
            .O(N__34275),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_14));
    InMux I__5999 (
            .O(N__34270),
            .I(N__34267));
    LocalMux I__5998 (
            .O(N__34267),
            .I(N__34264));
    Odrv4 I__5997 (
            .O(N__34264),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ));
    InMux I__5996 (
            .O(N__34261),
            .I(N__34258));
    LocalMux I__5995 (
            .O(N__34258),
            .I(N__34255));
    Span4Mux_v I__5994 (
            .O(N__34255),
            .I(N__34251));
    InMux I__5993 (
            .O(N__34254),
            .I(N__34248));
    Odrv4 I__5992 (
            .O(N__34251),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_12));
    LocalMux I__5991 (
            .O(N__34248),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_12));
    InMux I__5990 (
            .O(N__34243),
            .I(N__34240));
    LocalMux I__5989 (
            .O(N__34240),
            .I(N__34237));
    Odrv4 I__5988 (
            .O(N__34237),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ));
    InMux I__5987 (
            .O(N__34234),
            .I(N__34231));
    LocalMux I__5986 (
            .O(N__34231),
            .I(N__34228));
    Span4Mux_v I__5985 (
            .O(N__34228),
            .I(N__34224));
    InMux I__5984 (
            .O(N__34227),
            .I(N__34221));
    Span4Mux_h I__5983 (
            .O(N__34224),
            .I(N__34218));
    LocalMux I__5982 (
            .O(N__34221),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_15));
    Odrv4 I__5981 (
            .O(N__34218),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_15));
    InMux I__5980 (
            .O(N__34213),
            .I(N__34210));
    LocalMux I__5979 (
            .O(N__34210),
            .I(N__34207));
    Span4Mux_h I__5978 (
            .O(N__34207),
            .I(N__34204));
    Odrv4 I__5977 (
            .O(N__34204),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ));
    InMux I__5976 (
            .O(N__34201),
            .I(N__34198));
    LocalMux I__5975 (
            .O(N__34198),
            .I(N__34195));
    Span4Mux_h I__5974 (
            .O(N__34195),
            .I(N__34191));
    InMux I__5973 (
            .O(N__34194),
            .I(N__34188));
    Odrv4 I__5972 (
            .O(N__34191),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_11));
    LocalMux I__5971 (
            .O(N__34188),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_11));
    InMux I__5970 (
            .O(N__34183),
            .I(N__34180));
    LocalMux I__5969 (
            .O(N__34180),
            .I(N__34177));
    Odrv4 I__5968 (
            .O(N__34177),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ));
    InMux I__5967 (
            .O(N__34174),
            .I(N__34171));
    LocalMux I__5966 (
            .O(N__34171),
            .I(N__34168));
    Span4Mux_v I__5965 (
            .O(N__34168),
            .I(N__34164));
    InMux I__5964 (
            .O(N__34167),
            .I(N__34161));
    Odrv4 I__5963 (
            .O(N__34164),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_8));
    LocalMux I__5962 (
            .O(N__34161),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_8));
    CascadeMux I__5961 (
            .O(N__34156),
            .I(N__34153));
    InMux I__5960 (
            .O(N__34153),
            .I(N__34150));
    LocalMux I__5959 (
            .O(N__34150),
            .I(N__34147));
    Span4Mux_h I__5958 (
            .O(N__34147),
            .I(N__34144));
    Odrv4 I__5957 (
            .O(N__34144),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ));
    InMux I__5956 (
            .O(N__34141),
            .I(N__34138));
    LocalMux I__5955 (
            .O(N__34138),
            .I(N__34134));
    InMux I__5954 (
            .O(N__34137),
            .I(N__34131));
    Span4Mux_v I__5953 (
            .O(N__34134),
            .I(N__34128));
    LocalMux I__5952 (
            .O(N__34131),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_9));
    Odrv4 I__5951 (
            .O(N__34128),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_9));
    InMux I__5950 (
            .O(N__34123),
            .I(N__34120));
    LocalMux I__5949 (
            .O(N__34120),
            .I(N__34117));
    Odrv4 I__5948 (
            .O(N__34117),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ));
    InMux I__5947 (
            .O(N__34114),
            .I(N__34111));
    LocalMux I__5946 (
            .O(N__34111),
            .I(N__34108));
    Span4Mux_h I__5945 (
            .O(N__34108),
            .I(N__34104));
    InMux I__5944 (
            .O(N__34107),
            .I(N__34101));
    Odrv4 I__5943 (
            .O(N__34104),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_10));
    LocalMux I__5942 (
            .O(N__34101),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_10));
    CascadeMux I__5941 (
            .O(N__34096),
            .I(N__34093));
    InMux I__5940 (
            .O(N__34093),
            .I(N__34090));
    LocalMux I__5939 (
            .O(N__34090),
            .I(N__34087));
    Odrv4 I__5938 (
            .O(N__34087),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ));
    InMux I__5937 (
            .O(N__34084),
            .I(N__34081));
    LocalMux I__5936 (
            .O(N__34081),
            .I(N__34078));
    Span12Mux_v I__5935 (
            .O(N__34078),
            .I(N__34073));
    InMux I__5934 (
            .O(N__34077),
            .I(N__34068));
    InMux I__5933 (
            .O(N__34076),
            .I(N__34068));
    Odrv12 I__5932 (
            .O(N__34073),
            .I(\phase_controller_inst2.start_flagZ0 ));
    LocalMux I__5931 (
            .O(N__34068),
            .I(\phase_controller_inst2.start_flagZ0 ));
    InMux I__5930 (
            .O(N__34063),
            .I(N__34059));
    CascadeMux I__5929 (
            .O(N__34062),
            .I(N__34056));
    LocalMux I__5928 (
            .O(N__34059),
            .I(N__34052));
    InMux I__5927 (
            .O(N__34056),
            .I(N__34047));
    InMux I__5926 (
            .O(N__34055),
            .I(N__34047));
    Span4Mux_v I__5925 (
            .O(N__34052),
            .I(N__34044));
    LocalMux I__5924 (
            .O(N__34047),
            .I(N__34039));
    Span4Mux_v I__5923 (
            .O(N__34044),
            .I(N__34039));
    Odrv4 I__5922 (
            .O(N__34039),
            .I(\phase_controller_inst2.stateZ0Z_4 ));
    InMux I__5921 (
            .O(N__34036),
            .I(N__34029));
    InMux I__5920 (
            .O(N__34035),
            .I(N__34020));
    InMux I__5919 (
            .O(N__34034),
            .I(N__34020));
    InMux I__5918 (
            .O(N__34033),
            .I(N__34020));
    InMux I__5917 (
            .O(N__34032),
            .I(N__34020));
    LocalMux I__5916 (
            .O(N__34029),
            .I(N__34017));
    LocalMux I__5915 (
            .O(N__34020),
            .I(N__34014));
    Span4Mux_v I__5914 (
            .O(N__34017),
            .I(N__34009));
    Span4Mux_v I__5913 (
            .O(N__34014),
            .I(N__34009));
    Span4Mux_v I__5912 (
            .O(N__34009),
            .I(N__34005));
    InMux I__5911 (
            .O(N__34008),
            .I(N__34002));
    Sp12to4 I__5910 (
            .O(N__34005),
            .I(N__33997));
    LocalMux I__5909 (
            .O(N__34002),
            .I(N__33997));
    Span12Mux_h I__5908 (
            .O(N__33997),
            .I(N__33994));
    Odrv12 I__5907 (
            .O(N__33994),
            .I(start_stop_c));
    InMux I__5906 (
            .O(N__33991),
            .I(N__33986));
    InMux I__5905 (
            .O(N__33990),
            .I(N__33981));
    InMux I__5904 (
            .O(N__33989),
            .I(N__33981));
    LocalMux I__5903 (
            .O(N__33986),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    LocalMux I__5902 (
            .O(N__33981),
            .I(\phase_controller_inst1.stateZ0Z_4 ));
    CascadeMux I__5901 (
            .O(N__33976),
            .I(\phase_controller_inst1.state_ns_0_0_1_cascade_ ));
    CascadeMux I__5900 (
            .O(N__33973),
            .I(N__33969));
    InMux I__5899 (
            .O(N__33972),
            .I(N__33965));
    InMux I__5898 (
            .O(N__33969),
            .I(N__33960));
    InMux I__5897 (
            .O(N__33968),
            .I(N__33960));
    LocalMux I__5896 (
            .O(N__33965),
            .I(\phase_controller_inst1.start_flagZ0 ));
    LocalMux I__5895 (
            .O(N__33960),
            .I(\phase_controller_inst1.start_flagZ0 ));
    CascadeMux I__5894 (
            .O(N__33955),
            .I(\phase_controller_inst1.stoper_tr.un4_start_0_cascade_ ));
    CascadeMux I__5893 (
            .O(N__33952),
            .I(N__33947));
    CascadeMux I__5892 (
            .O(N__33951),
            .I(N__33944));
    InMux I__5891 (
            .O(N__33950),
            .I(N__33937));
    InMux I__5890 (
            .O(N__33947),
            .I(N__33937));
    InMux I__5889 (
            .O(N__33944),
            .I(N__33937));
    LocalMux I__5888 (
            .O(N__33937),
            .I(\phase_controller_inst1.tr_time_passed ));
    InMux I__5887 (
            .O(N__33934),
            .I(N__33928));
    InMux I__5886 (
            .O(N__33933),
            .I(N__33928));
    LocalMux I__5885 (
            .O(N__33928),
            .I(\phase_controller_inst1.stateZ0Z_0 ));
    InMux I__5884 (
            .O(N__33925),
            .I(N__33922));
    LocalMux I__5883 (
            .O(N__33922),
            .I(N__33919));
    Span4Mux_h I__5882 (
            .O(N__33919),
            .I(N__33916));
    Odrv4 I__5881 (
            .O(N__33916),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ));
    InMux I__5880 (
            .O(N__33913),
            .I(N__33901));
    InMux I__5879 (
            .O(N__33912),
            .I(N__33901));
    InMux I__5878 (
            .O(N__33911),
            .I(N__33901));
    InMux I__5877 (
            .O(N__33910),
            .I(N__33901));
    LocalMux I__5876 (
            .O(N__33901),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ));
    InMux I__5875 (
            .O(N__33898),
            .I(N__33893));
    InMux I__5874 (
            .O(N__33897),
            .I(N__33888));
    InMux I__5873 (
            .O(N__33896),
            .I(N__33888));
    LocalMux I__5872 (
            .O(N__33893),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    LocalMux I__5871 (
            .O(N__33888),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ));
    InMux I__5870 (
            .O(N__33883),
            .I(N__33878));
    InMux I__5869 (
            .O(N__33882),
            .I(N__33875));
    InMux I__5868 (
            .O(N__33881),
            .I(N__33872));
    LocalMux I__5867 (
            .O(N__33878),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    LocalMux I__5866 (
            .O(N__33875),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    LocalMux I__5865 (
            .O(N__33872),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ));
    CascadeMux I__5864 (
            .O(N__33865),
            .I(N__33862));
    InMux I__5863 (
            .O(N__33862),
            .I(N__33859));
    LocalMux I__5862 (
            .O(N__33859),
            .I(N__33856));
    Span4Mux_h I__5861 (
            .O(N__33856),
            .I(N__33853));
    Odrv4 I__5860 (
            .O(N__33853),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt30 ));
    InMux I__5859 (
            .O(N__33850),
            .I(N__33847));
    LocalMux I__5858 (
            .O(N__33847),
            .I(N__33844));
    Span4Mux_h I__5857 (
            .O(N__33844),
            .I(N__33840));
    InMux I__5856 (
            .O(N__33843),
            .I(N__33837));
    Odrv4 I__5855 (
            .O(N__33840),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    LocalMux I__5854 (
            .O(N__33837),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ));
    InMux I__5853 (
            .O(N__33832),
            .I(N__33829));
    LocalMux I__5852 (
            .O(N__33829),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13));
    CascadeMux I__5851 (
            .O(N__33826),
            .I(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_));
    InMux I__5850 (
            .O(N__33823),
            .I(N__33820));
    LocalMux I__5849 (
            .O(N__33820),
            .I(N__33817));
    Odrv4 I__5848 (
            .O(N__33817),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ));
    InMux I__5847 (
            .O(N__33814),
            .I(N__33811));
    LocalMux I__5846 (
            .O(N__33811),
            .I(N__33808));
    Span4Mux_h I__5845 (
            .O(N__33808),
            .I(N__33804));
    InMux I__5844 (
            .O(N__33807),
            .I(N__33801));
    Odrv4 I__5843 (
            .O(N__33804),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    LocalMux I__5842 (
            .O(N__33801),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ));
    InMux I__5841 (
            .O(N__33796),
            .I(N__33793));
    LocalMux I__5840 (
            .O(N__33793),
            .I(N__33789));
    InMux I__5839 (
            .O(N__33792),
            .I(N__33786));
    Span12Mux_v I__5838 (
            .O(N__33789),
            .I(N__33783));
    LocalMux I__5837 (
            .O(N__33786),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    Odrv12 I__5836 (
            .O(N__33783),
            .I(elapsed_time_ns_1_RNIV9PBB_0_21));
    InMux I__5835 (
            .O(N__33778),
            .I(N__33773));
    InMux I__5834 (
            .O(N__33777),
            .I(N__33762));
    InMux I__5833 (
            .O(N__33776),
            .I(N__33762));
    LocalMux I__5832 (
            .O(N__33773),
            .I(N__33759));
    InMux I__5831 (
            .O(N__33772),
            .I(N__33754));
    InMux I__5830 (
            .O(N__33771),
            .I(N__33754));
    InMux I__5829 (
            .O(N__33770),
            .I(N__33744));
    InMux I__5828 (
            .O(N__33769),
            .I(N__33744));
    InMux I__5827 (
            .O(N__33768),
            .I(N__33741));
    InMux I__5826 (
            .O(N__33767),
            .I(N__33738));
    LocalMux I__5825 (
            .O(N__33762),
            .I(N__33735));
    Span4Mux_h I__5824 (
            .O(N__33759),
            .I(N__33730));
    LocalMux I__5823 (
            .O(N__33754),
            .I(N__33730));
    InMux I__5822 (
            .O(N__33753),
            .I(N__33714));
    InMux I__5821 (
            .O(N__33752),
            .I(N__33714));
    InMux I__5820 (
            .O(N__33751),
            .I(N__33714));
    InMux I__5819 (
            .O(N__33750),
            .I(N__33714));
    InMux I__5818 (
            .O(N__33749),
            .I(N__33711));
    LocalMux I__5817 (
            .O(N__33744),
            .I(N__33704));
    LocalMux I__5816 (
            .O(N__33741),
            .I(N__33704));
    LocalMux I__5815 (
            .O(N__33738),
            .I(N__33699));
    Span4Mux_v I__5814 (
            .O(N__33735),
            .I(N__33699));
    Span4Mux_v I__5813 (
            .O(N__33730),
            .I(N__33696));
    InMux I__5812 (
            .O(N__33729),
            .I(N__33686));
    InMux I__5811 (
            .O(N__33728),
            .I(N__33686));
    CascadeMux I__5810 (
            .O(N__33727),
            .I(N__33683));
    InMux I__5809 (
            .O(N__33726),
            .I(N__33672));
    InMux I__5808 (
            .O(N__33725),
            .I(N__33672));
    InMux I__5807 (
            .O(N__33724),
            .I(N__33672));
    InMux I__5806 (
            .O(N__33723),
            .I(N__33672));
    LocalMux I__5805 (
            .O(N__33714),
            .I(N__33667));
    LocalMux I__5804 (
            .O(N__33711),
            .I(N__33667));
    InMux I__5803 (
            .O(N__33710),
            .I(N__33662));
    InMux I__5802 (
            .O(N__33709),
            .I(N__33662));
    Span4Mux_v I__5801 (
            .O(N__33704),
            .I(N__33659));
    Sp12to4 I__5800 (
            .O(N__33699),
            .I(N__33654));
    Sp12to4 I__5799 (
            .O(N__33696),
            .I(N__33654));
    InMux I__5798 (
            .O(N__33695),
            .I(N__33649));
    InMux I__5797 (
            .O(N__33694),
            .I(N__33649));
    InMux I__5796 (
            .O(N__33693),
            .I(N__33642));
    InMux I__5795 (
            .O(N__33692),
            .I(N__33642));
    InMux I__5794 (
            .O(N__33691),
            .I(N__33642));
    LocalMux I__5793 (
            .O(N__33686),
            .I(N__33639));
    InMux I__5792 (
            .O(N__33683),
            .I(N__33632));
    InMux I__5791 (
            .O(N__33682),
            .I(N__33632));
    InMux I__5790 (
            .O(N__33681),
            .I(N__33632));
    LocalMux I__5789 (
            .O(N__33672),
            .I(N__33627));
    Span4Mux_h I__5788 (
            .O(N__33667),
            .I(N__33627));
    LocalMux I__5787 (
            .O(N__33662),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5786 (
            .O(N__33659),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__5785 (
            .O(N__33654),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5784 (
            .O(N__33649),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5783 (
            .O(N__33642),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv12 I__5782 (
            .O(N__33639),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    LocalMux I__5781 (
            .O(N__33632),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    Odrv4 I__5780 (
            .O(N__33627),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3 ));
    InMux I__5779 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__5778 (
            .O(N__33607),
            .I(N__33604));
    Span4Mux_v I__5777 (
            .O(N__33604),
            .I(N__33600));
    InMux I__5776 (
            .O(N__33603),
            .I(N__33597));
    Odrv4 I__5775 (
            .O(N__33600),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    LocalMux I__5774 (
            .O(N__33597),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ));
    InMux I__5773 (
            .O(N__33592),
            .I(N__33589));
    LocalMux I__5772 (
            .O(N__33589),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30));
    CascadeMux I__5771 (
            .O(N__33586),
            .I(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_));
    InMux I__5770 (
            .O(N__33583),
            .I(N__33580));
    LocalMux I__5769 (
            .O(N__33580),
            .I(N__33577));
    Span4Mux_h I__5768 (
            .O(N__33577),
            .I(N__33574));
    Odrv4 I__5767 (
            .O(N__33574),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ));
    InMux I__5766 (
            .O(N__33571),
            .I(N__33565));
    InMux I__5765 (
            .O(N__33570),
            .I(N__33565));
    LocalMux I__5764 (
            .O(N__33565),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ));
    InMux I__5763 (
            .O(N__33562),
            .I(N__33555));
    InMux I__5762 (
            .O(N__33561),
            .I(N__33555));
    InMux I__5761 (
            .O(N__33560),
            .I(N__33552));
    LocalMux I__5760 (
            .O(N__33555),
            .I(N__33549));
    LocalMux I__5759 (
            .O(N__33552),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ));
    Odrv4 I__5758 (
            .O(N__33549),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ));
    CascadeMux I__5757 (
            .O(N__33544),
            .I(N__33540));
    CascadeMux I__5756 (
            .O(N__33543),
            .I(N__33537));
    InMux I__5755 (
            .O(N__33540),
            .I(N__33532));
    InMux I__5754 (
            .O(N__33537),
            .I(N__33532));
    LocalMux I__5753 (
            .O(N__33532),
            .I(N__33529));
    Span4Mux_h I__5752 (
            .O(N__33529),
            .I(N__33526));
    Odrv4 I__5751 (
            .O(N__33526),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ));
    InMux I__5750 (
            .O(N__33523),
            .I(N__33516));
    InMux I__5749 (
            .O(N__33522),
            .I(N__33516));
    InMux I__5748 (
            .O(N__33521),
            .I(N__33513));
    LocalMux I__5747 (
            .O(N__33516),
            .I(N__33510));
    LocalMux I__5746 (
            .O(N__33513),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ));
    Odrv4 I__5745 (
            .O(N__33510),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ));
    CascadeMux I__5744 (
            .O(N__33505),
            .I(N__33502));
    InMux I__5743 (
            .O(N__33502),
            .I(N__33499));
    LocalMux I__5742 (
            .O(N__33499),
            .I(N__33496));
    Odrv4 I__5741 (
            .O(N__33496),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ));
    InMux I__5740 (
            .O(N__33493),
            .I(N__33490));
    LocalMux I__5739 (
            .O(N__33490),
            .I(N__33487));
    Odrv4 I__5738 (
            .O(N__33487),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt26 ));
    InMux I__5737 (
            .O(N__33484),
            .I(N__33478));
    InMux I__5736 (
            .O(N__33483),
            .I(N__33478));
    LocalMux I__5735 (
            .O(N__33478),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ));
    InMux I__5734 (
            .O(N__33475),
            .I(N__33468));
    InMux I__5733 (
            .O(N__33474),
            .I(N__33468));
    InMux I__5732 (
            .O(N__33473),
            .I(N__33465));
    LocalMux I__5731 (
            .O(N__33468),
            .I(N__33462));
    LocalMux I__5730 (
            .O(N__33465),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ));
    Odrv4 I__5729 (
            .O(N__33462),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ));
    CascadeMux I__5728 (
            .O(N__33457),
            .I(N__33453));
    CascadeMux I__5727 (
            .O(N__33456),
            .I(N__33450));
    InMux I__5726 (
            .O(N__33453),
            .I(N__33445));
    InMux I__5725 (
            .O(N__33450),
            .I(N__33445));
    LocalMux I__5724 (
            .O(N__33445),
            .I(N__33441));
    InMux I__5723 (
            .O(N__33444),
            .I(N__33438));
    Span4Mux_v I__5722 (
            .O(N__33441),
            .I(N__33435));
    LocalMux I__5721 (
            .O(N__33438),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ));
    Odrv4 I__5720 (
            .O(N__33435),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ));
    CascadeMux I__5719 (
            .O(N__33430),
            .I(N__33427));
    InMux I__5718 (
            .O(N__33427),
            .I(N__33424));
    LocalMux I__5717 (
            .O(N__33424),
            .I(N__33421));
    Span4Mux_h I__5716 (
            .O(N__33421),
            .I(N__33418));
    Odrv4 I__5715 (
            .O(N__33418),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ));
    InMux I__5714 (
            .O(N__33415),
            .I(N__33409));
    InMux I__5713 (
            .O(N__33414),
            .I(N__33409));
    LocalMux I__5712 (
            .O(N__33409),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ));
    InMux I__5711 (
            .O(N__33406),
            .I(N__33403));
    LocalMux I__5710 (
            .O(N__33403),
            .I(N__33400));
    Span4Mux_h I__5709 (
            .O(N__33400),
            .I(N__33397));
    Odrv4 I__5708 (
            .O(N__33397),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt28 ));
    InMux I__5707 (
            .O(N__33394),
            .I(N__33389));
    InMux I__5706 (
            .O(N__33393),
            .I(N__33384));
    InMux I__5705 (
            .O(N__33392),
            .I(N__33384));
    LocalMux I__5704 (
            .O(N__33389),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ));
    LocalMux I__5703 (
            .O(N__33384),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ));
    InMux I__5702 (
            .O(N__33379),
            .I(N__33374));
    InMux I__5701 (
            .O(N__33378),
            .I(N__33369));
    InMux I__5700 (
            .O(N__33377),
            .I(N__33369));
    LocalMux I__5699 (
            .O(N__33374),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ));
    LocalMux I__5698 (
            .O(N__33369),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ));
    CascadeMux I__5697 (
            .O(N__33364),
            .I(N__33361));
    InMux I__5696 (
            .O(N__33361),
            .I(N__33358));
    LocalMux I__5695 (
            .O(N__33358),
            .I(N__33355));
    Span4Mux_v I__5694 (
            .O(N__33355),
            .I(N__33352));
    Odrv4 I__5693 (
            .O(N__33352),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ));
    InMux I__5692 (
            .O(N__33349),
            .I(N__33343));
    InMux I__5691 (
            .O(N__33348),
            .I(N__33343));
    LocalMux I__5690 (
            .O(N__33343),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ));
    InMux I__5689 (
            .O(N__33340),
            .I(N__33334));
    InMux I__5688 (
            .O(N__33339),
            .I(N__33334));
    LocalMux I__5687 (
            .O(N__33334),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ));
    InMux I__5686 (
            .O(N__33331),
            .I(N__33325));
    InMux I__5685 (
            .O(N__33330),
            .I(N__33325));
    LocalMux I__5684 (
            .O(N__33325),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ));
    InMux I__5683 (
            .O(N__33322),
            .I(N__33310));
    InMux I__5682 (
            .O(N__33321),
            .I(N__33310));
    InMux I__5681 (
            .O(N__33320),
            .I(N__33310));
    InMux I__5680 (
            .O(N__33319),
            .I(N__33310));
    LocalMux I__5679 (
            .O(N__33310),
            .I(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ));
    InMux I__5678 (
            .O(N__33307),
            .I(N__33304));
    LocalMux I__5677 (
            .O(N__33304),
            .I(N__33301));
    Odrv4 I__5676 (
            .O(N__33301),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt24 ));
    InMux I__5675 (
            .O(N__33298),
            .I(N__33295));
    LocalMux I__5674 (
            .O(N__33295),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ));
    InMux I__5673 (
            .O(N__33292),
            .I(N__33289));
    LocalMux I__5672 (
            .O(N__33289),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ));
    InMux I__5671 (
            .O(N__33286),
            .I(N__33283));
    LocalMux I__5670 (
            .O(N__33283),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt16 ));
    InMux I__5669 (
            .O(N__33280),
            .I(N__33274));
    InMux I__5668 (
            .O(N__33279),
            .I(N__33274));
    LocalMux I__5667 (
            .O(N__33274),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ));
    InMux I__5666 (
            .O(N__33271),
            .I(N__33265));
    InMux I__5665 (
            .O(N__33270),
            .I(N__33265));
    LocalMux I__5664 (
            .O(N__33265),
            .I(N__33261));
    InMux I__5663 (
            .O(N__33264),
            .I(N__33258));
    Span4Mux_h I__5662 (
            .O(N__33261),
            .I(N__33255));
    LocalMux I__5661 (
            .O(N__33258),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ));
    Odrv4 I__5660 (
            .O(N__33255),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ));
    CascadeMux I__5659 (
            .O(N__33250),
            .I(N__33246));
    CascadeMux I__5658 (
            .O(N__33249),
            .I(N__33243));
    InMux I__5657 (
            .O(N__33246),
            .I(N__33238));
    InMux I__5656 (
            .O(N__33243),
            .I(N__33238));
    LocalMux I__5655 (
            .O(N__33238),
            .I(N__33234));
    InMux I__5654 (
            .O(N__33237),
            .I(N__33231));
    Span4Mux_h I__5653 (
            .O(N__33234),
            .I(N__33228));
    LocalMux I__5652 (
            .O(N__33231),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ));
    Odrv4 I__5651 (
            .O(N__33228),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ));
    CascadeMux I__5650 (
            .O(N__33223),
            .I(N__33220));
    InMux I__5649 (
            .O(N__33220),
            .I(N__33217));
    LocalMux I__5648 (
            .O(N__33217),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ));
    InMux I__5647 (
            .O(N__33214),
            .I(N__33208));
    InMux I__5646 (
            .O(N__33213),
            .I(N__33208));
    LocalMux I__5645 (
            .O(N__33208),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ));
    InMux I__5644 (
            .O(N__33205),
            .I(N__33201));
    InMux I__5643 (
            .O(N__33204),
            .I(N__33198));
    LocalMux I__5642 (
            .O(N__33201),
            .I(N__33195));
    LocalMux I__5641 (
            .O(N__33198),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ));
    Odrv4 I__5640 (
            .O(N__33195),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ));
    InMux I__5639 (
            .O(N__33190),
            .I(N__33186));
    InMux I__5638 (
            .O(N__33189),
            .I(N__33182));
    LocalMux I__5637 (
            .O(N__33186),
            .I(N__33179));
    InMux I__5636 (
            .O(N__33185),
            .I(N__33176));
    LocalMux I__5635 (
            .O(N__33182),
            .I(N__33171));
    Span4Mux_h I__5634 (
            .O(N__33179),
            .I(N__33171));
    LocalMux I__5633 (
            .O(N__33176),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    Odrv4 I__5632 (
            .O(N__33171),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ));
    CascadeMux I__5631 (
            .O(N__33166),
            .I(N__33162));
    CascadeMux I__5630 (
            .O(N__33165),
            .I(N__33159));
    InMux I__5629 (
            .O(N__33162),
            .I(N__33156));
    InMux I__5628 (
            .O(N__33159),
            .I(N__33153));
    LocalMux I__5627 (
            .O(N__33156),
            .I(N__33149));
    LocalMux I__5626 (
            .O(N__33153),
            .I(N__33146));
    InMux I__5625 (
            .O(N__33152),
            .I(N__33143));
    Span4Mux_h I__5624 (
            .O(N__33149),
            .I(N__33140));
    Span4Mux_h I__5623 (
            .O(N__33146),
            .I(N__33137));
    LocalMux I__5622 (
            .O(N__33143),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    Odrv4 I__5621 (
            .O(N__33140),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    Odrv4 I__5620 (
            .O(N__33137),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ));
    CascadeMux I__5619 (
            .O(N__33130),
            .I(N__33127));
    InMux I__5618 (
            .O(N__33127),
            .I(N__33124));
    LocalMux I__5617 (
            .O(N__33124),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ));
    InMux I__5616 (
            .O(N__33121),
            .I(N__33117));
    InMux I__5615 (
            .O(N__33120),
            .I(N__33114));
    LocalMux I__5614 (
            .O(N__33117),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ));
    LocalMux I__5613 (
            .O(N__33114),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ));
    InMux I__5612 (
            .O(N__33109),
            .I(N__33103));
    InMux I__5611 (
            .O(N__33108),
            .I(N__33103));
    LocalMux I__5610 (
            .O(N__33103),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ));
    InMux I__5609 (
            .O(N__33100),
            .I(N__33097));
    LocalMux I__5608 (
            .O(N__33097),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ));
    InMux I__5607 (
            .O(N__33094),
            .I(N__33091));
    LocalMux I__5606 (
            .O(N__33091),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ));
    InMux I__5605 (
            .O(N__33088),
            .I(N__33085));
    LocalMux I__5604 (
            .O(N__33085),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ));
    InMux I__5603 (
            .O(N__33082),
            .I(N__33079));
    LocalMux I__5602 (
            .O(N__33079),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ));
    CascadeMux I__5601 (
            .O(N__33076),
            .I(N__33073));
    InMux I__5600 (
            .O(N__33073),
            .I(N__33070));
    LocalMux I__5599 (
            .O(N__33070),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ));
    InMux I__5598 (
            .O(N__33067),
            .I(N__33064));
    LocalMux I__5597 (
            .O(N__33064),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ));
    InMux I__5596 (
            .O(N__33061),
            .I(N__33058));
    LocalMux I__5595 (
            .O(N__33058),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ));
    InMux I__5594 (
            .O(N__33055),
            .I(N__33052));
    LocalMux I__5593 (
            .O(N__33052),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ));
    InMux I__5592 (
            .O(N__33049),
            .I(N__33046));
    LocalMux I__5591 (
            .O(N__33046),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ));
    CascadeMux I__5590 (
            .O(N__33043),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ));
    InMux I__5589 (
            .O(N__33040),
            .I(N__33037));
    LocalMux I__5588 (
            .O(N__33037),
            .I(N__33034));
    Odrv4 I__5587 (
            .O(N__33034),
            .I(\current_shift_inst.PI_CTRL.N_46_21 ));
    InMux I__5586 (
            .O(N__33031),
            .I(N__33028));
    LocalMux I__5585 (
            .O(N__33028),
            .I(N__33025));
    Odrv4 I__5584 (
            .O(N__33025),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ));
    InMux I__5583 (
            .O(N__33022),
            .I(N__33019));
    LocalMux I__5582 (
            .O(N__33019),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ));
    InMux I__5581 (
            .O(N__33016),
            .I(N__33013));
    LocalMux I__5580 (
            .O(N__33013),
            .I(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ));
    InMux I__5579 (
            .O(N__33010),
            .I(N__33007));
    LocalMux I__5578 (
            .O(N__33007),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ));
    InMux I__5577 (
            .O(N__33004),
            .I(N__33001));
    LocalMux I__5576 (
            .O(N__33001),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ));
    InMux I__5575 (
            .O(N__32998),
            .I(N__32995));
    LocalMux I__5574 (
            .O(N__32995),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ));
    InMux I__5573 (
            .O(N__32992),
            .I(N__32989));
    LocalMux I__5572 (
            .O(N__32989),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ));
    CascadeMux I__5571 (
            .O(N__32986),
            .I(N__32983));
    InMux I__5570 (
            .O(N__32983),
            .I(N__32980));
    LocalMux I__5569 (
            .O(N__32980),
            .I(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ));
    InMux I__5568 (
            .O(N__32977),
            .I(N__32974));
    LocalMux I__5567 (
            .O(N__32974),
            .I(N__32971));
    Span4Mux_h I__5566 (
            .O(N__32971),
            .I(N__32968));
    Odrv4 I__5565 (
            .O(N__32968),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ));
    CascadeMux I__5564 (
            .O(N__32965),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ));
    InMux I__5563 (
            .O(N__32962),
            .I(N__32959));
    LocalMux I__5562 (
            .O(N__32959),
            .I(\current_shift_inst.PI_CTRL.N_47 ));
    CascadeMux I__5561 (
            .O(N__32956),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ));
    InMux I__5560 (
            .O(N__32953),
            .I(N__32950));
    LocalMux I__5559 (
            .O(N__32950),
            .I(\current_shift_inst.PI_CTRL.N_77 ));
    InMux I__5558 (
            .O(N__32947),
            .I(N__32944));
    LocalMux I__5557 (
            .O(N__32944),
            .I(\current_shift_inst.PI_CTRL.N_43 ));
    CascadeMux I__5556 (
            .O(N__32941),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ));
    InMux I__5555 (
            .O(N__32938),
            .I(N__32935));
    LocalMux I__5554 (
            .O(N__32935),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ));
    InMux I__5553 (
            .O(N__32932),
            .I(N__32929));
    LocalMux I__5552 (
            .O(N__32929),
            .I(\current_shift_inst.PI_CTRL.N_46_16 ));
    InMux I__5551 (
            .O(N__32926),
            .I(N__32919));
    InMux I__5550 (
            .O(N__32925),
            .I(N__32919));
    CEMux I__5549 (
            .O(N__32924),
            .I(N__32895));
    LocalMux I__5548 (
            .O(N__32919),
            .I(N__32892));
    InMux I__5547 (
            .O(N__32918),
            .I(N__32883));
    InMux I__5546 (
            .O(N__32917),
            .I(N__32883));
    InMux I__5545 (
            .O(N__32916),
            .I(N__32883));
    InMux I__5544 (
            .O(N__32915),
            .I(N__32883));
    InMux I__5543 (
            .O(N__32914),
            .I(N__32874));
    InMux I__5542 (
            .O(N__32913),
            .I(N__32871));
    InMux I__5541 (
            .O(N__32912),
            .I(N__32858));
    InMux I__5540 (
            .O(N__32911),
            .I(N__32858));
    InMux I__5539 (
            .O(N__32910),
            .I(N__32858));
    InMux I__5538 (
            .O(N__32909),
            .I(N__32858));
    InMux I__5537 (
            .O(N__32908),
            .I(N__32858));
    InMux I__5536 (
            .O(N__32907),
            .I(N__32858));
    InMux I__5535 (
            .O(N__32906),
            .I(N__32843));
    InMux I__5534 (
            .O(N__32905),
            .I(N__32843));
    InMux I__5533 (
            .O(N__32904),
            .I(N__32843));
    InMux I__5532 (
            .O(N__32903),
            .I(N__32843));
    InMux I__5531 (
            .O(N__32902),
            .I(N__32843));
    InMux I__5530 (
            .O(N__32901),
            .I(N__32843));
    InMux I__5529 (
            .O(N__32900),
            .I(N__32843));
    InMux I__5528 (
            .O(N__32899),
            .I(N__32838));
    InMux I__5527 (
            .O(N__32898),
            .I(N__32838));
    LocalMux I__5526 (
            .O(N__32895),
            .I(N__32835));
    Span4Mux_v I__5525 (
            .O(N__32892),
            .I(N__32830));
    LocalMux I__5524 (
            .O(N__32883),
            .I(N__32830));
    InMux I__5523 (
            .O(N__32882),
            .I(N__32825));
    InMux I__5522 (
            .O(N__32881),
            .I(N__32825));
    InMux I__5521 (
            .O(N__32880),
            .I(N__32822));
    InMux I__5520 (
            .O(N__32879),
            .I(N__32819));
    InMux I__5519 (
            .O(N__32878),
            .I(N__32814));
    InMux I__5518 (
            .O(N__32877),
            .I(N__32814));
    LocalMux I__5517 (
            .O(N__32874),
            .I(N__32811));
    LocalMux I__5516 (
            .O(N__32871),
            .I(N__32808));
    LocalMux I__5515 (
            .O(N__32858),
            .I(N__32803));
    LocalMux I__5514 (
            .O(N__32843),
            .I(N__32803));
    LocalMux I__5513 (
            .O(N__32838),
            .I(N__32796));
    Span4Mux_v I__5512 (
            .O(N__32835),
            .I(N__32796));
    Span4Mux_v I__5511 (
            .O(N__32830),
            .I(N__32796));
    LocalMux I__5510 (
            .O(N__32825),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__5509 (
            .O(N__32822),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__5508 (
            .O(N__32819),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    LocalMux I__5507 (
            .O(N__32814),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv12 I__5506 (
            .O(N__32811),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__5505 (
            .O(N__32808),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__5504 (
            .O(N__32803),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    Odrv4 I__5503 (
            .O(N__32796),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0 ));
    InMux I__5502 (
            .O(N__32779),
            .I(N__32776));
    LocalMux I__5501 (
            .O(N__32776),
            .I(N__32773));
    Odrv4 I__5500 (
            .O(N__32773),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ));
    CascadeMux I__5499 (
            .O(N__32770),
            .I(N__32767));
    InMux I__5498 (
            .O(N__32767),
            .I(N__32764));
    LocalMux I__5497 (
            .O(N__32764),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt22 ));
    InMux I__5496 (
            .O(N__32761),
            .I(N__32758));
    LocalMux I__5495 (
            .O(N__32758),
            .I(N__32755));
    Span4Mux_h I__5494 (
            .O(N__32755),
            .I(N__32751));
    InMux I__5493 (
            .O(N__32754),
            .I(N__32748));
    Odrv4 I__5492 (
            .O(N__32751),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_22));
    LocalMux I__5491 (
            .O(N__32748),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_22));
    InMux I__5490 (
            .O(N__32743),
            .I(N__32736));
    InMux I__5489 (
            .O(N__32742),
            .I(N__32736));
    InMux I__5488 (
            .O(N__32741),
            .I(N__32733));
    LocalMux I__5487 (
            .O(N__32736),
            .I(N__32730));
    LocalMux I__5486 (
            .O(N__32733),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    Odrv4 I__5485 (
            .O(N__32730),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ));
    InMux I__5484 (
            .O(N__32725),
            .I(N__32719));
    InMux I__5483 (
            .O(N__32724),
            .I(N__32719));
    LocalMux I__5482 (
            .O(N__32719),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ));
    CascadeMux I__5481 (
            .O(N__32716),
            .I(N__32712));
    CascadeMux I__5480 (
            .O(N__32715),
            .I(N__32709));
    InMux I__5479 (
            .O(N__32712),
            .I(N__32703));
    InMux I__5478 (
            .O(N__32709),
            .I(N__32703));
    InMux I__5477 (
            .O(N__32708),
            .I(N__32700));
    LocalMux I__5476 (
            .O(N__32703),
            .I(N__32697));
    LocalMux I__5475 (
            .O(N__32700),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    Odrv4 I__5474 (
            .O(N__32697),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ));
    InMux I__5473 (
            .O(N__32692),
            .I(N__32689));
    LocalMux I__5472 (
            .O(N__32689),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ));
    InMux I__5471 (
            .O(N__32686),
            .I(N__32683));
    LocalMux I__5470 (
            .O(N__32683),
            .I(N__32680));
    Span4Mux_h I__5469 (
            .O(N__32680),
            .I(N__32676));
    InMux I__5468 (
            .O(N__32679),
            .I(N__32673));
    Odrv4 I__5467 (
            .O(N__32676),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_23));
    LocalMux I__5466 (
            .O(N__32673),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_23));
    InMux I__5465 (
            .O(N__32668),
            .I(N__32662));
    InMux I__5464 (
            .O(N__32667),
            .I(N__32662));
    LocalMux I__5463 (
            .O(N__32662),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ));
    InMux I__5462 (
            .O(N__32659),
            .I(N__32647));
    InMux I__5461 (
            .O(N__32658),
            .I(N__32647));
    InMux I__5460 (
            .O(N__32657),
            .I(N__32647));
    InMux I__5459 (
            .O(N__32656),
            .I(N__32647));
    LocalMux I__5458 (
            .O(N__32647),
            .I(N__32644));
    Span4Mux_h I__5457 (
            .O(N__32644),
            .I(N__32641));
    Odrv4 I__5456 (
            .O(N__32641),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ));
    CEMux I__5455 (
            .O(N__32638),
            .I(N__32632));
    CEMux I__5454 (
            .O(N__32637),
            .I(N__32629));
    CEMux I__5453 (
            .O(N__32636),
            .I(N__32626));
    CEMux I__5452 (
            .O(N__32635),
            .I(N__32623));
    LocalMux I__5451 (
            .O(N__32632),
            .I(N__32620));
    LocalMux I__5450 (
            .O(N__32629),
            .I(N__32616));
    LocalMux I__5449 (
            .O(N__32626),
            .I(N__32612));
    LocalMux I__5448 (
            .O(N__32623),
            .I(N__32609));
    Span4Mux_v I__5447 (
            .O(N__32620),
            .I(N__32606));
    CEMux I__5446 (
            .O(N__32619),
            .I(N__32603));
    Span4Mux_v I__5445 (
            .O(N__32616),
            .I(N__32600));
    CEMux I__5444 (
            .O(N__32615),
            .I(N__32597));
    Span4Mux_h I__5443 (
            .O(N__32612),
            .I(N__32593));
    Span4Mux_h I__5442 (
            .O(N__32609),
            .I(N__32582));
    Span4Mux_h I__5441 (
            .O(N__32606),
            .I(N__32582));
    LocalMux I__5440 (
            .O(N__32603),
            .I(N__32582));
    Span4Mux_v I__5439 (
            .O(N__32600),
            .I(N__32582));
    LocalMux I__5438 (
            .O(N__32597),
            .I(N__32582));
    CEMux I__5437 (
            .O(N__32596),
            .I(N__32579));
    Span4Mux_v I__5436 (
            .O(N__32593),
            .I(N__32576));
    Span4Mux_v I__5435 (
            .O(N__32582),
            .I(N__32571));
    LocalMux I__5434 (
            .O(N__32579),
            .I(N__32571));
    Span4Mux_v I__5433 (
            .O(N__32576),
            .I(N__32568));
    Span4Mux_v I__5432 (
            .O(N__32571),
            .I(N__32565));
    Odrv4 I__5431 (
            .O(N__32568),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    Odrv4 I__5430 (
            .O(N__32565),
            .I(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ));
    InMux I__5429 (
            .O(N__32560),
            .I(N__32557));
    LocalMux I__5428 (
            .O(N__32557),
            .I(N__32552));
    InMux I__5427 (
            .O(N__32556),
            .I(N__32549));
    CascadeMux I__5426 (
            .O(N__32555),
            .I(N__32546));
    Span4Mux_v I__5425 (
            .O(N__32552),
            .I(N__32541));
    LocalMux I__5424 (
            .O(N__32549),
            .I(N__32538));
    InMux I__5423 (
            .O(N__32546),
            .I(N__32530));
    InMux I__5422 (
            .O(N__32545),
            .I(N__32530));
    InMux I__5421 (
            .O(N__32544),
            .I(N__32530));
    Span4Mux_h I__5420 (
            .O(N__32541),
            .I(N__32525));
    Span4Mux_v I__5419 (
            .O(N__32538),
            .I(N__32525));
    InMux I__5418 (
            .O(N__32537),
            .I(N__32522));
    LocalMux I__5417 (
            .O(N__32530),
            .I(N__32519));
    Sp12to4 I__5416 (
            .O(N__32525),
            .I(N__32516));
    LocalMux I__5415 (
            .O(N__32522),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv4 I__5414 (
            .O(N__32519),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    Odrv12 I__5413 (
            .O(N__32516),
            .I(\phase_controller_inst2.stoper_tr.start_latchedZ0 ));
    InMux I__5412 (
            .O(N__32509),
            .I(N__32471));
    InMux I__5411 (
            .O(N__32508),
            .I(N__32471));
    InMux I__5410 (
            .O(N__32507),
            .I(N__32471));
    InMux I__5409 (
            .O(N__32506),
            .I(N__32462));
    InMux I__5408 (
            .O(N__32505),
            .I(N__32462));
    InMux I__5407 (
            .O(N__32504),
            .I(N__32462));
    InMux I__5406 (
            .O(N__32503),
            .I(N__32462));
    InMux I__5405 (
            .O(N__32502),
            .I(N__32453));
    InMux I__5404 (
            .O(N__32501),
            .I(N__32453));
    InMux I__5403 (
            .O(N__32500),
            .I(N__32453));
    InMux I__5402 (
            .O(N__32499),
            .I(N__32453));
    InMux I__5401 (
            .O(N__32498),
            .I(N__32442));
    InMux I__5400 (
            .O(N__32497),
            .I(N__32442));
    InMux I__5399 (
            .O(N__32496),
            .I(N__32442));
    InMux I__5398 (
            .O(N__32495),
            .I(N__32442));
    InMux I__5397 (
            .O(N__32494),
            .I(N__32442));
    InMux I__5396 (
            .O(N__32493),
            .I(N__32433));
    InMux I__5395 (
            .O(N__32492),
            .I(N__32433));
    InMux I__5394 (
            .O(N__32491),
            .I(N__32433));
    InMux I__5393 (
            .O(N__32490),
            .I(N__32433));
    InMux I__5392 (
            .O(N__32489),
            .I(N__32424));
    InMux I__5391 (
            .O(N__32488),
            .I(N__32424));
    InMux I__5390 (
            .O(N__32487),
            .I(N__32424));
    InMux I__5389 (
            .O(N__32486),
            .I(N__32424));
    InMux I__5388 (
            .O(N__32485),
            .I(N__32415));
    InMux I__5387 (
            .O(N__32484),
            .I(N__32415));
    InMux I__5386 (
            .O(N__32483),
            .I(N__32415));
    InMux I__5385 (
            .O(N__32482),
            .I(N__32415));
    InMux I__5384 (
            .O(N__32481),
            .I(N__32406));
    InMux I__5383 (
            .O(N__32480),
            .I(N__32406));
    InMux I__5382 (
            .O(N__32479),
            .I(N__32406));
    InMux I__5381 (
            .O(N__32478),
            .I(N__32406));
    LocalMux I__5380 (
            .O(N__32471),
            .I(N__32403));
    LocalMux I__5379 (
            .O(N__32462),
            .I(N__32398));
    LocalMux I__5378 (
            .O(N__32453),
            .I(N__32398));
    LocalMux I__5377 (
            .O(N__32442),
            .I(N__32395));
    LocalMux I__5376 (
            .O(N__32433),
            .I(N__32390));
    LocalMux I__5375 (
            .O(N__32424),
            .I(N__32390));
    LocalMux I__5374 (
            .O(N__32415),
            .I(N__32381));
    LocalMux I__5373 (
            .O(N__32406),
            .I(N__32381));
    Span4Mux_v I__5372 (
            .O(N__32403),
            .I(N__32381));
    Span4Mux_v I__5371 (
            .O(N__32398),
            .I(N__32381));
    Span4Mux_v I__5370 (
            .O(N__32395),
            .I(N__32374));
    Span4Mux_v I__5369 (
            .O(N__32390),
            .I(N__32374));
    Span4Mux_h I__5368 (
            .O(N__32381),
            .I(N__32374));
    Odrv4 I__5367 (
            .O(N__32374),
            .I(\phase_controller_inst2.stoper_tr.start_latched_i_0 ));
    CascadeMux I__5366 (
            .O(N__32371),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ));
    InMux I__5365 (
            .O(N__32368),
            .I(N__32362));
    InMux I__5364 (
            .O(N__32367),
            .I(N__32362));
    LocalMux I__5363 (
            .O(N__32362),
            .I(N__32358));
    InMux I__5362 (
            .O(N__32361),
            .I(N__32355));
    Span4Mux_h I__5361 (
            .O(N__32358),
            .I(N__32352));
    LocalMux I__5360 (
            .O(N__32355),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    Odrv4 I__5359 (
            .O(N__32352),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ));
    InMux I__5358 (
            .O(N__32347),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_26 ));
    InMux I__5357 (
            .O(N__32344),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_27 ));
    InMux I__5356 (
            .O(N__32341),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_28 ));
    InMux I__5355 (
            .O(N__32338),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_29 ));
    InMux I__5354 (
            .O(N__32335),
            .I(N__32303));
    InMux I__5353 (
            .O(N__32334),
            .I(N__32303));
    InMux I__5352 (
            .O(N__32333),
            .I(N__32303));
    InMux I__5351 (
            .O(N__32332),
            .I(N__32303));
    InMux I__5350 (
            .O(N__32331),
            .I(N__32294));
    InMux I__5349 (
            .O(N__32330),
            .I(N__32294));
    InMux I__5348 (
            .O(N__32329),
            .I(N__32294));
    InMux I__5347 (
            .O(N__32328),
            .I(N__32294));
    InMux I__5346 (
            .O(N__32327),
            .I(N__32285));
    InMux I__5345 (
            .O(N__32326),
            .I(N__32285));
    InMux I__5344 (
            .O(N__32325),
            .I(N__32285));
    InMux I__5343 (
            .O(N__32324),
            .I(N__32285));
    InMux I__5342 (
            .O(N__32323),
            .I(N__32276));
    InMux I__5341 (
            .O(N__32322),
            .I(N__32276));
    InMux I__5340 (
            .O(N__32321),
            .I(N__32276));
    InMux I__5339 (
            .O(N__32320),
            .I(N__32276));
    InMux I__5338 (
            .O(N__32319),
            .I(N__32259));
    InMux I__5337 (
            .O(N__32318),
            .I(N__32259));
    InMux I__5336 (
            .O(N__32317),
            .I(N__32259));
    InMux I__5335 (
            .O(N__32316),
            .I(N__32259));
    InMux I__5334 (
            .O(N__32315),
            .I(N__32250));
    InMux I__5333 (
            .O(N__32314),
            .I(N__32250));
    InMux I__5332 (
            .O(N__32313),
            .I(N__32250));
    InMux I__5331 (
            .O(N__32312),
            .I(N__32250));
    LocalMux I__5330 (
            .O(N__32303),
            .I(N__32247));
    LocalMux I__5329 (
            .O(N__32294),
            .I(N__32244));
    LocalMux I__5328 (
            .O(N__32285),
            .I(N__32241));
    LocalMux I__5327 (
            .O(N__32276),
            .I(N__32238));
    InMux I__5326 (
            .O(N__32275),
            .I(N__32229));
    InMux I__5325 (
            .O(N__32274),
            .I(N__32229));
    InMux I__5324 (
            .O(N__32273),
            .I(N__32229));
    InMux I__5323 (
            .O(N__32272),
            .I(N__32229));
    InMux I__5322 (
            .O(N__32271),
            .I(N__32220));
    InMux I__5321 (
            .O(N__32270),
            .I(N__32220));
    InMux I__5320 (
            .O(N__32269),
            .I(N__32220));
    InMux I__5319 (
            .O(N__32268),
            .I(N__32220));
    LocalMux I__5318 (
            .O(N__32259),
            .I(N__32215));
    LocalMux I__5317 (
            .O(N__32250),
            .I(N__32215));
    Span4Mux_h I__5316 (
            .O(N__32247),
            .I(N__32210));
    Span4Mux_h I__5315 (
            .O(N__32244),
            .I(N__32210));
    Span4Mux_h I__5314 (
            .O(N__32241),
            .I(N__32205));
    Span4Mux_h I__5313 (
            .O(N__32238),
            .I(N__32205));
    LocalMux I__5312 (
            .O(N__32229),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    LocalMux I__5311 (
            .O(N__32220),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    Odrv4 I__5310 (
            .O(N__32215),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    Odrv4 I__5309 (
            .O(N__32210),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    Odrv4 I__5308 (
            .O(N__32205),
            .I(\phase_controller_inst1.stoper_tr.start_latched_i_0 ));
    InMux I__5307 (
            .O(N__32194),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_30 ));
    CEMux I__5306 (
            .O(N__32191),
            .I(N__32179));
    CEMux I__5305 (
            .O(N__32190),
            .I(N__32179));
    CEMux I__5304 (
            .O(N__32189),
            .I(N__32179));
    CEMux I__5303 (
            .O(N__32188),
            .I(N__32179));
    GlobalMux I__5302 (
            .O(N__32179),
            .I(N__32176));
    gio2CtrlBuf I__5301 (
            .O(N__32176),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0_g ));
    CascadeMux I__5300 (
            .O(N__32173),
            .I(N__32170));
    InMux I__5299 (
            .O(N__32170),
            .I(N__32167));
    LocalMux I__5298 (
            .O(N__32167),
            .I(N__32164));
    Odrv4 I__5297 (
            .O(N__32164),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt20 ));
    InMux I__5296 (
            .O(N__32161),
            .I(N__32158));
    LocalMux I__5295 (
            .O(N__32158),
            .I(N__32155));
    Span4Mux_h I__5294 (
            .O(N__32155),
            .I(N__32151));
    InMux I__5293 (
            .O(N__32154),
            .I(N__32148));
    Odrv4 I__5292 (
            .O(N__32151),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_20));
    LocalMux I__5291 (
            .O(N__32148),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_20));
    InMux I__5290 (
            .O(N__32143),
            .I(N__32137));
    InMux I__5289 (
            .O(N__32142),
            .I(N__32137));
    LocalMux I__5288 (
            .O(N__32137),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ));
    InMux I__5287 (
            .O(N__32134),
            .I(N__32128));
    InMux I__5286 (
            .O(N__32133),
            .I(N__32128));
    LocalMux I__5285 (
            .O(N__32128),
            .I(N__32125));
    Odrv12 I__5284 (
            .O(N__32125),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ));
    CascadeMux I__5283 (
            .O(N__32122),
            .I(N__32118));
    CascadeMux I__5282 (
            .O(N__32121),
            .I(N__32115));
    InMux I__5281 (
            .O(N__32118),
            .I(N__32109));
    InMux I__5280 (
            .O(N__32115),
            .I(N__32109));
    InMux I__5279 (
            .O(N__32114),
            .I(N__32106));
    LocalMux I__5278 (
            .O(N__32109),
            .I(N__32103));
    LocalMux I__5277 (
            .O(N__32106),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    Odrv4 I__5276 (
            .O(N__32103),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ));
    InMux I__5275 (
            .O(N__32098),
            .I(N__32091));
    InMux I__5274 (
            .O(N__32097),
            .I(N__32091));
    InMux I__5273 (
            .O(N__32096),
            .I(N__32088));
    LocalMux I__5272 (
            .O(N__32091),
            .I(N__32085));
    LocalMux I__5271 (
            .O(N__32088),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    Odrv4 I__5270 (
            .O(N__32085),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ));
    InMux I__5269 (
            .O(N__32080),
            .I(N__32077));
    LocalMux I__5268 (
            .O(N__32077),
            .I(N__32074));
    Span4Mux_h I__5267 (
            .O(N__32074),
            .I(N__32071));
    Odrv4 I__5266 (
            .O(N__32071),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ));
    InMux I__5265 (
            .O(N__32068),
            .I(N__32061));
    InMux I__5264 (
            .O(N__32067),
            .I(N__32061));
    InMux I__5263 (
            .O(N__32066),
            .I(N__32058));
    LocalMux I__5262 (
            .O(N__32061),
            .I(N__32055));
    LocalMux I__5261 (
            .O(N__32058),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ));
    Odrv12 I__5260 (
            .O(N__32055),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ));
    InMux I__5259 (
            .O(N__32050),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_17 ));
    InMux I__5258 (
            .O(N__32047),
            .I(N__32040));
    InMux I__5257 (
            .O(N__32046),
            .I(N__32040));
    InMux I__5256 (
            .O(N__32045),
            .I(N__32037));
    LocalMux I__5255 (
            .O(N__32040),
            .I(N__32034));
    LocalMux I__5254 (
            .O(N__32037),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ));
    Odrv12 I__5253 (
            .O(N__32034),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ));
    InMux I__5252 (
            .O(N__32029),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_18 ));
    InMux I__5251 (
            .O(N__32026),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_19 ));
    InMux I__5250 (
            .O(N__32023),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_20 ));
    InMux I__5249 (
            .O(N__32020),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_21 ));
    InMux I__5248 (
            .O(N__32017),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_22 ));
    InMux I__5247 (
            .O(N__32014),
            .I(N__32008));
    InMux I__5246 (
            .O(N__32013),
            .I(N__32008));
    LocalMux I__5245 (
            .O(N__32008),
            .I(N__32004));
    InMux I__5244 (
            .O(N__32007),
            .I(N__32001));
    Span4Mux_h I__5243 (
            .O(N__32004),
            .I(N__31998));
    LocalMux I__5242 (
            .O(N__32001),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    Odrv4 I__5241 (
            .O(N__31998),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ));
    InMux I__5240 (
            .O(N__31993),
            .I(bfn_11_16_0_));
    InMux I__5239 (
            .O(N__31990),
            .I(N__31984));
    InMux I__5238 (
            .O(N__31989),
            .I(N__31984));
    LocalMux I__5237 (
            .O(N__31984),
            .I(N__31980));
    InMux I__5236 (
            .O(N__31983),
            .I(N__31977));
    Span4Mux_h I__5235 (
            .O(N__31980),
            .I(N__31974));
    LocalMux I__5234 (
            .O(N__31977),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    Odrv4 I__5233 (
            .O(N__31974),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ));
    InMux I__5232 (
            .O(N__31969),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_24 ));
    CascadeMux I__5231 (
            .O(N__31966),
            .I(N__31962));
    CascadeMux I__5230 (
            .O(N__31965),
            .I(N__31959));
    InMux I__5229 (
            .O(N__31962),
            .I(N__31954));
    InMux I__5228 (
            .O(N__31959),
            .I(N__31954));
    LocalMux I__5227 (
            .O(N__31954),
            .I(N__31950));
    InMux I__5226 (
            .O(N__31953),
            .I(N__31947));
    Span4Mux_h I__5225 (
            .O(N__31950),
            .I(N__31944));
    LocalMux I__5224 (
            .O(N__31947),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ));
    Odrv4 I__5223 (
            .O(N__31944),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ));
    InMux I__5222 (
            .O(N__31939),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_25 ));
    InMux I__5221 (
            .O(N__31936),
            .I(N__31933));
    LocalMux I__5220 (
            .O(N__31933),
            .I(N__31929));
    InMux I__5219 (
            .O(N__31932),
            .I(N__31926));
    Span4Mux_h I__5218 (
            .O(N__31929),
            .I(N__31923));
    LocalMux I__5217 (
            .O(N__31926),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ));
    Odrv4 I__5216 (
            .O(N__31923),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ));
    InMux I__5215 (
            .O(N__31918),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_9 ));
    InMux I__5214 (
            .O(N__31915),
            .I(N__31911));
    InMux I__5213 (
            .O(N__31914),
            .I(N__31908));
    LocalMux I__5212 (
            .O(N__31911),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ));
    LocalMux I__5211 (
            .O(N__31908),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ));
    InMux I__5210 (
            .O(N__31903),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_10 ));
    InMux I__5209 (
            .O(N__31900),
            .I(N__31896));
    InMux I__5208 (
            .O(N__31899),
            .I(N__31893));
    LocalMux I__5207 (
            .O(N__31896),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ));
    LocalMux I__5206 (
            .O(N__31893),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ));
    InMux I__5205 (
            .O(N__31888),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_11 ));
    InMux I__5204 (
            .O(N__31885),
            .I(N__31881));
    InMux I__5203 (
            .O(N__31884),
            .I(N__31878));
    LocalMux I__5202 (
            .O(N__31881),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ));
    LocalMux I__5201 (
            .O(N__31878),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ));
    InMux I__5200 (
            .O(N__31873),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_12 ));
    InMux I__5199 (
            .O(N__31870),
            .I(N__31866));
    InMux I__5198 (
            .O(N__31869),
            .I(N__31863));
    LocalMux I__5197 (
            .O(N__31866),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ));
    LocalMux I__5196 (
            .O(N__31863),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ));
    InMux I__5195 (
            .O(N__31858),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_13 ));
    InMux I__5194 (
            .O(N__31855),
            .I(N__31851));
    InMux I__5193 (
            .O(N__31854),
            .I(N__31848));
    LocalMux I__5192 (
            .O(N__31851),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ));
    LocalMux I__5191 (
            .O(N__31848),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ));
    InMux I__5190 (
            .O(N__31843),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_14 ));
    CascadeMux I__5189 (
            .O(N__31840),
            .I(N__31836));
    CascadeMux I__5188 (
            .O(N__31839),
            .I(N__31833));
    InMux I__5187 (
            .O(N__31836),
            .I(N__31828));
    InMux I__5186 (
            .O(N__31833),
            .I(N__31828));
    LocalMux I__5185 (
            .O(N__31828),
            .I(N__31824));
    InMux I__5184 (
            .O(N__31827),
            .I(N__31821));
    Span4Mux_h I__5183 (
            .O(N__31824),
            .I(N__31818));
    LocalMux I__5182 (
            .O(N__31821),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    Odrv4 I__5181 (
            .O(N__31818),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ));
    InMux I__5180 (
            .O(N__31813),
            .I(bfn_11_15_0_));
    InMux I__5179 (
            .O(N__31810),
            .I(N__31804));
    InMux I__5178 (
            .O(N__31809),
            .I(N__31804));
    LocalMux I__5177 (
            .O(N__31804),
            .I(N__31800));
    InMux I__5176 (
            .O(N__31803),
            .I(N__31797));
    Span4Mux_h I__5175 (
            .O(N__31800),
            .I(N__31794));
    LocalMux I__5174 (
            .O(N__31797),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    Odrv4 I__5173 (
            .O(N__31794),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ));
    InMux I__5172 (
            .O(N__31789),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_16 ));
    InMux I__5171 (
            .O(N__31786),
            .I(N__31782));
    InMux I__5170 (
            .O(N__31785),
            .I(N__31779));
    LocalMux I__5169 (
            .O(N__31782),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ));
    LocalMux I__5168 (
            .O(N__31779),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ));
    InMux I__5167 (
            .O(N__31774),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_0 ));
    InMux I__5166 (
            .O(N__31771),
            .I(N__31767));
    InMux I__5165 (
            .O(N__31770),
            .I(N__31764));
    LocalMux I__5164 (
            .O(N__31767),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ));
    LocalMux I__5163 (
            .O(N__31764),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ));
    InMux I__5162 (
            .O(N__31759),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_1 ));
    InMux I__5161 (
            .O(N__31756),
            .I(N__31752));
    InMux I__5160 (
            .O(N__31755),
            .I(N__31749));
    LocalMux I__5159 (
            .O(N__31752),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ));
    LocalMux I__5158 (
            .O(N__31749),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ));
    InMux I__5157 (
            .O(N__31744),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_2 ));
    InMux I__5156 (
            .O(N__31741),
            .I(N__31737));
    InMux I__5155 (
            .O(N__31740),
            .I(N__31734));
    LocalMux I__5154 (
            .O(N__31737),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ));
    LocalMux I__5153 (
            .O(N__31734),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ));
    InMux I__5152 (
            .O(N__31729),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_3 ));
    InMux I__5151 (
            .O(N__31726),
            .I(N__31722));
    InMux I__5150 (
            .O(N__31725),
            .I(N__31719));
    LocalMux I__5149 (
            .O(N__31722),
            .I(N__31716));
    LocalMux I__5148 (
            .O(N__31719),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ));
    Odrv4 I__5147 (
            .O(N__31716),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ));
    InMux I__5146 (
            .O(N__31711),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_4 ));
    InMux I__5145 (
            .O(N__31708),
            .I(N__31704));
    InMux I__5144 (
            .O(N__31707),
            .I(N__31701));
    LocalMux I__5143 (
            .O(N__31704),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ));
    LocalMux I__5142 (
            .O(N__31701),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ));
    InMux I__5141 (
            .O(N__31696),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_5 ));
    InMux I__5140 (
            .O(N__31693),
            .I(N__31689));
    InMux I__5139 (
            .O(N__31692),
            .I(N__31686));
    LocalMux I__5138 (
            .O(N__31689),
            .I(N__31683));
    LocalMux I__5137 (
            .O(N__31686),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ));
    Odrv4 I__5136 (
            .O(N__31683),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ));
    InMux I__5135 (
            .O(N__31678),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_6 ));
    InMux I__5134 (
            .O(N__31675),
            .I(N__31671));
    InMux I__5133 (
            .O(N__31674),
            .I(N__31668));
    LocalMux I__5132 (
            .O(N__31671),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ));
    LocalMux I__5131 (
            .O(N__31668),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ));
    InMux I__5130 (
            .O(N__31663),
            .I(bfn_11_14_0_));
    InMux I__5129 (
            .O(N__31660),
            .I(N__31656));
    InMux I__5128 (
            .O(N__31659),
            .I(N__31653));
    LocalMux I__5127 (
            .O(N__31656),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ));
    LocalMux I__5126 (
            .O(N__31653),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ));
    InMux I__5125 (
            .O(N__31648),
            .I(\phase_controller_inst1.stoper_tr.counter_cry_8 ));
    InMux I__5124 (
            .O(N__31645),
            .I(bfn_11_12_0_));
    InMux I__5123 (
            .O(N__31642),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_24 ));
    InMux I__5122 (
            .O(N__31639),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_25 ));
    InMux I__5121 (
            .O(N__31636),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_26 ));
    InMux I__5120 (
            .O(N__31633),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_27 ));
    InMux I__5119 (
            .O(N__31630),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_28 ));
    InMux I__5118 (
            .O(N__31627),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_29 ));
    InMux I__5117 (
            .O(N__31624),
            .I(N__31590));
    InMux I__5116 (
            .O(N__31623),
            .I(N__31590));
    InMux I__5115 (
            .O(N__31622),
            .I(N__31590));
    InMux I__5114 (
            .O(N__31621),
            .I(N__31579));
    InMux I__5113 (
            .O(N__31620),
            .I(N__31579));
    InMux I__5112 (
            .O(N__31619),
            .I(N__31579));
    InMux I__5111 (
            .O(N__31618),
            .I(N__31579));
    InMux I__5110 (
            .O(N__31617),
            .I(N__31579));
    InMux I__5109 (
            .O(N__31616),
            .I(N__31566));
    InMux I__5108 (
            .O(N__31615),
            .I(N__31566));
    InMux I__5107 (
            .O(N__31614),
            .I(N__31566));
    InMux I__5106 (
            .O(N__31613),
            .I(N__31566));
    InMux I__5105 (
            .O(N__31612),
            .I(N__31557));
    InMux I__5104 (
            .O(N__31611),
            .I(N__31557));
    InMux I__5103 (
            .O(N__31610),
            .I(N__31557));
    InMux I__5102 (
            .O(N__31609),
            .I(N__31557));
    InMux I__5101 (
            .O(N__31608),
            .I(N__31548));
    InMux I__5100 (
            .O(N__31607),
            .I(N__31548));
    InMux I__5099 (
            .O(N__31606),
            .I(N__31548));
    InMux I__5098 (
            .O(N__31605),
            .I(N__31548));
    InMux I__5097 (
            .O(N__31604),
            .I(N__31539));
    InMux I__5096 (
            .O(N__31603),
            .I(N__31539));
    InMux I__5095 (
            .O(N__31602),
            .I(N__31539));
    InMux I__5094 (
            .O(N__31601),
            .I(N__31539));
    InMux I__5093 (
            .O(N__31600),
            .I(N__31530));
    InMux I__5092 (
            .O(N__31599),
            .I(N__31530));
    InMux I__5091 (
            .O(N__31598),
            .I(N__31530));
    InMux I__5090 (
            .O(N__31597),
            .I(N__31530));
    LocalMux I__5089 (
            .O(N__31590),
            .I(N__31527));
    LocalMux I__5088 (
            .O(N__31579),
            .I(N__31524));
    InMux I__5087 (
            .O(N__31578),
            .I(N__31515));
    InMux I__5086 (
            .O(N__31577),
            .I(N__31515));
    InMux I__5085 (
            .O(N__31576),
            .I(N__31515));
    InMux I__5084 (
            .O(N__31575),
            .I(N__31515));
    LocalMux I__5083 (
            .O(N__31566),
            .I(N__31500));
    LocalMux I__5082 (
            .O(N__31557),
            .I(N__31500));
    LocalMux I__5081 (
            .O(N__31548),
            .I(N__31500));
    LocalMux I__5080 (
            .O(N__31539),
            .I(N__31500));
    LocalMux I__5079 (
            .O(N__31530),
            .I(N__31500));
    Span4Mux_v I__5078 (
            .O(N__31527),
            .I(N__31500));
    Span4Mux_v I__5077 (
            .O(N__31524),
            .I(N__31500));
    LocalMux I__5076 (
            .O(N__31515),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    Odrv4 I__5075 (
            .O(N__31500),
            .I(\phase_controller_inst2.stoper_hc.start_latched_i_0 ));
    InMux I__5074 (
            .O(N__31495),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_30 ));
    CEMux I__5073 (
            .O(N__31492),
            .I(N__31486));
    CEMux I__5072 (
            .O(N__31491),
            .I(N__31483));
    CEMux I__5071 (
            .O(N__31490),
            .I(N__31480));
    CEMux I__5070 (
            .O(N__31489),
            .I(N__31477));
    LocalMux I__5069 (
            .O(N__31486),
            .I(N__31474));
    LocalMux I__5068 (
            .O(N__31483),
            .I(N__31469));
    LocalMux I__5067 (
            .O(N__31480),
            .I(N__31469));
    LocalMux I__5066 (
            .O(N__31477),
            .I(N__31466));
    Span4Mux_v I__5065 (
            .O(N__31474),
            .I(N__31463));
    Span4Mux_v I__5064 (
            .O(N__31469),
            .I(N__31460));
    Span4Mux_h I__5063 (
            .O(N__31466),
            .I(N__31457));
    Span4Mux_h I__5062 (
            .O(N__31463),
            .I(N__31452));
    Span4Mux_h I__5061 (
            .O(N__31460),
            .I(N__31452));
    Odrv4 I__5060 (
            .O(N__31457),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    Odrv4 I__5059 (
            .O(N__31452),
            .I(\phase_controller_inst2.stoper_hc.un2_start_0 ));
    CascadeMux I__5058 (
            .O(N__31447),
            .I(N__31443));
    InMux I__5057 (
            .O(N__31446),
            .I(N__31440));
    InMux I__5056 (
            .O(N__31443),
            .I(N__31437));
    LocalMux I__5055 (
            .O(N__31440),
            .I(N__31432));
    LocalMux I__5054 (
            .O(N__31437),
            .I(N__31432));
    Span4Mux_v I__5053 (
            .O(N__31432),
            .I(N__31429));
    Odrv4 I__5052 (
            .O(N__31429),
            .I(\phase_controller_inst1.stoper_tr.counter ));
    InMux I__5051 (
            .O(N__31426),
            .I(N__31422));
    InMux I__5050 (
            .O(N__31425),
            .I(N__31419));
    LocalMux I__5049 (
            .O(N__31422),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ));
    LocalMux I__5048 (
            .O(N__31419),
            .I(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ));
    InMux I__5047 (
            .O(N__31414),
            .I(bfn_11_11_0_));
    InMux I__5046 (
            .O(N__31411),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_16 ));
    InMux I__5045 (
            .O(N__31408),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_17 ));
    InMux I__5044 (
            .O(N__31405),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_18 ));
    InMux I__5043 (
            .O(N__31402),
            .I(N__31395));
    InMux I__5042 (
            .O(N__31401),
            .I(N__31395));
    InMux I__5041 (
            .O(N__31400),
            .I(N__31392));
    LocalMux I__5040 (
            .O(N__31395),
            .I(N__31389));
    LocalMux I__5039 (
            .O(N__31392),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ));
    Odrv4 I__5038 (
            .O(N__31389),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ));
    InMux I__5037 (
            .O(N__31384),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_19 ));
    CascadeMux I__5036 (
            .O(N__31381),
            .I(N__31377));
    CascadeMux I__5035 (
            .O(N__31380),
            .I(N__31374));
    InMux I__5034 (
            .O(N__31377),
            .I(N__31368));
    InMux I__5033 (
            .O(N__31374),
            .I(N__31368));
    InMux I__5032 (
            .O(N__31373),
            .I(N__31365));
    LocalMux I__5031 (
            .O(N__31368),
            .I(N__31362));
    LocalMux I__5030 (
            .O(N__31365),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ));
    Odrv4 I__5029 (
            .O(N__31362),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ));
    InMux I__5028 (
            .O(N__31357),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_20 ));
    CascadeMux I__5027 (
            .O(N__31354),
            .I(N__31350));
    InMux I__5026 (
            .O(N__31353),
            .I(N__31345));
    InMux I__5025 (
            .O(N__31350),
            .I(N__31345));
    LocalMux I__5024 (
            .O(N__31345),
            .I(N__31341));
    InMux I__5023 (
            .O(N__31344),
            .I(N__31338));
    Span4Mux_h I__5022 (
            .O(N__31341),
            .I(N__31335));
    LocalMux I__5021 (
            .O(N__31338),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ));
    Odrv4 I__5020 (
            .O(N__31335),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ));
    InMux I__5019 (
            .O(N__31330),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_21 ));
    CascadeMux I__5018 (
            .O(N__31327),
            .I(N__31323));
    InMux I__5017 (
            .O(N__31326),
            .I(N__31318));
    InMux I__5016 (
            .O(N__31323),
            .I(N__31318));
    LocalMux I__5015 (
            .O(N__31318),
            .I(N__31314));
    InMux I__5014 (
            .O(N__31317),
            .I(N__31311));
    Span4Mux_h I__5013 (
            .O(N__31314),
            .I(N__31308));
    LocalMux I__5012 (
            .O(N__31311),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ));
    Odrv4 I__5011 (
            .O(N__31308),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ));
    InMux I__5010 (
            .O(N__31303),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_22 ));
    InMux I__5009 (
            .O(N__31300),
            .I(N__31297));
    LocalMux I__5008 (
            .O(N__31297),
            .I(N__31293));
    InMux I__5007 (
            .O(N__31296),
            .I(N__31290));
    Span4Mux_v I__5006 (
            .O(N__31293),
            .I(N__31287));
    LocalMux I__5005 (
            .O(N__31290),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ));
    Odrv4 I__5004 (
            .O(N__31287),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ));
    InMux I__5003 (
            .O(N__31282),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_6 ));
    InMux I__5002 (
            .O(N__31279),
            .I(N__31276));
    LocalMux I__5001 (
            .O(N__31276),
            .I(N__31272));
    InMux I__5000 (
            .O(N__31275),
            .I(N__31269));
    Span4Mux_v I__4999 (
            .O(N__31272),
            .I(N__31266));
    LocalMux I__4998 (
            .O(N__31269),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ));
    Odrv4 I__4997 (
            .O(N__31266),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ));
    InMux I__4996 (
            .O(N__31261),
            .I(bfn_11_10_0_));
    InMux I__4995 (
            .O(N__31258),
            .I(N__31254));
    InMux I__4994 (
            .O(N__31257),
            .I(N__31251));
    LocalMux I__4993 (
            .O(N__31254),
            .I(N__31248));
    LocalMux I__4992 (
            .O(N__31251),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ));
    Odrv12 I__4991 (
            .O(N__31248),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ));
    InMux I__4990 (
            .O(N__31243),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_8 ));
    InMux I__4989 (
            .O(N__31240),
            .I(N__31236));
    InMux I__4988 (
            .O(N__31239),
            .I(N__31233));
    LocalMux I__4987 (
            .O(N__31236),
            .I(N__31230));
    LocalMux I__4986 (
            .O(N__31233),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ));
    Odrv12 I__4985 (
            .O(N__31230),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ));
    InMux I__4984 (
            .O(N__31225),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_9 ));
    InMux I__4983 (
            .O(N__31222),
            .I(N__31218));
    InMux I__4982 (
            .O(N__31221),
            .I(N__31215));
    LocalMux I__4981 (
            .O(N__31218),
            .I(N__31212));
    LocalMux I__4980 (
            .O(N__31215),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ));
    Odrv12 I__4979 (
            .O(N__31212),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ));
    InMux I__4978 (
            .O(N__31207),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_10 ));
    InMux I__4977 (
            .O(N__31204),
            .I(N__31200));
    InMux I__4976 (
            .O(N__31203),
            .I(N__31197));
    LocalMux I__4975 (
            .O(N__31200),
            .I(N__31194));
    LocalMux I__4974 (
            .O(N__31197),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ));
    Odrv12 I__4973 (
            .O(N__31194),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ));
    InMux I__4972 (
            .O(N__31189),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_11 ));
    InMux I__4971 (
            .O(N__31186),
            .I(N__31183));
    LocalMux I__4970 (
            .O(N__31183),
            .I(N__31179));
    InMux I__4969 (
            .O(N__31182),
            .I(N__31176));
    Span4Mux_v I__4968 (
            .O(N__31179),
            .I(N__31173));
    LocalMux I__4967 (
            .O(N__31176),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ));
    Odrv4 I__4966 (
            .O(N__31173),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ));
    InMux I__4965 (
            .O(N__31168),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_12 ));
    InMux I__4964 (
            .O(N__31165),
            .I(N__31161));
    InMux I__4963 (
            .O(N__31164),
            .I(N__31158));
    LocalMux I__4962 (
            .O(N__31161),
            .I(N__31155));
    LocalMux I__4961 (
            .O(N__31158),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ));
    Odrv12 I__4960 (
            .O(N__31155),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ));
    InMux I__4959 (
            .O(N__31150),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_13 ));
    InMux I__4958 (
            .O(N__31147),
            .I(N__31144));
    LocalMux I__4957 (
            .O(N__31144),
            .I(N__31140));
    InMux I__4956 (
            .O(N__31143),
            .I(N__31137));
    Span4Mux_v I__4955 (
            .O(N__31140),
            .I(N__31134));
    LocalMux I__4954 (
            .O(N__31137),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ));
    Odrv4 I__4953 (
            .O(N__31134),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ));
    InMux I__4952 (
            .O(N__31129),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_14 ));
    CascadeMux I__4951 (
            .O(N__31126),
            .I(N__31123));
    InMux I__4950 (
            .O(N__31123),
            .I(N__31120));
    LocalMux I__4949 (
            .O(N__31120),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ));
    CascadeMux I__4948 (
            .O(N__31117),
            .I(N__31113));
    InMux I__4947 (
            .O(N__31116),
            .I(N__31110));
    InMux I__4946 (
            .O(N__31113),
            .I(N__31107));
    LocalMux I__4945 (
            .O(N__31110),
            .I(\phase_controller_inst2.stoper_hc.counter ));
    LocalMux I__4944 (
            .O(N__31107),
            .I(\phase_controller_inst2.stoper_hc.counter ));
    InMux I__4943 (
            .O(N__31102),
            .I(N__31098));
    InMux I__4942 (
            .O(N__31101),
            .I(N__31095));
    LocalMux I__4941 (
            .O(N__31098),
            .I(N__31092));
    LocalMux I__4940 (
            .O(N__31095),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ));
    Odrv12 I__4939 (
            .O(N__31092),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ));
    InMux I__4938 (
            .O(N__31087),
            .I(N__31084));
    LocalMux I__4937 (
            .O(N__31084),
            .I(N__31080));
    InMux I__4936 (
            .O(N__31083),
            .I(N__31077));
    Span4Mux_v I__4935 (
            .O(N__31080),
            .I(N__31074));
    LocalMux I__4934 (
            .O(N__31077),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ));
    Odrv4 I__4933 (
            .O(N__31074),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ));
    InMux I__4932 (
            .O(N__31069),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_0 ));
    InMux I__4931 (
            .O(N__31066),
            .I(N__31062));
    InMux I__4930 (
            .O(N__31065),
            .I(N__31059));
    LocalMux I__4929 (
            .O(N__31062),
            .I(N__31056));
    LocalMux I__4928 (
            .O(N__31059),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ));
    Odrv12 I__4927 (
            .O(N__31056),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ));
    InMux I__4926 (
            .O(N__31051),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_1 ));
    InMux I__4925 (
            .O(N__31048),
            .I(N__31044));
    CascadeMux I__4924 (
            .O(N__31047),
            .I(N__31041));
    LocalMux I__4923 (
            .O(N__31044),
            .I(N__31038));
    InMux I__4922 (
            .O(N__31041),
            .I(N__31035));
    Span4Mux_h I__4921 (
            .O(N__31038),
            .I(N__31032));
    LocalMux I__4920 (
            .O(N__31035),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ));
    Odrv4 I__4919 (
            .O(N__31032),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ));
    InMux I__4918 (
            .O(N__31027),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_2 ));
    InMux I__4917 (
            .O(N__31024),
            .I(N__31020));
    InMux I__4916 (
            .O(N__31023),
            .I(N__31017));
    LocalMux I__4915 (
            .O(N__31020),
            .I(N__31014));
    LocalMux I__4914 (
            .O(N__31017),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ));
    Odrv12 I__4913 (
            .O(N__31014),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ));
    InMux I__4912 (
            .O(N__31009),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_3 ));
    InMux I__4911 (
            .O(N__31006),
            .I(N__31002));
    InMux I__4910 (
            .O(N__31005),
            .I(N__30999));
    LocalMux I__4909 (
            .O(N__31002),
            .I(N__30996));
    LocalMux I__4908 (
            .O(N__30999),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ));
    Odrv12 I__4907 (
            .O(N__30996),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ));
    InMux I__4906 (
            .O(N__30991),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_4 ));
    InMux I__4905 (
            .O(N__30988),
            .I(N__30984));
    InMux I__4904 (
            .O(N__30987),
            .I(N__30981));
    LocalMux I__4903 (
            .O(N__30984),
            .I(N__30978));
    LocalMux I__4902 (
            .O(N__30981),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ));
    Odrv12 I__4901 (
            .O(N__30978),
            .I(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ));
    InMux I__4900 (
            .O(N__30973),
            .I(\phase_controller_inst2.stoper_hc.counter_cry_5 ));
    InMux I__4899 (
            .O(N__30970),
            .I(bfn_11_8_0_));
    InMux I__4898 (
            .O(N__30967),
            .I(N__30964));
    LocalMux I__4897 (
            .O(N__30964),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt20 ));
    InMux I__4896 (
            .O(N__30961),
            .I(N__30958));
    LocalMux I__4895 (
            .O(N__30958),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt18 ));
    CascadeMux I__4894 (
            .O(N__30955),
            .I(N__30951));
    CascadeMux I__4893 (
            .O(N__30954),
            .I(N__30948));
    InMux I__4892 (
            .O(N__30951),
            .I(N__30945));
    InMux I__4891 (
            .O(N__30948),
            .I(N__30942));
    LocalMux I__4890 (
            .O(N__30945),
            .I(N__30939));
    LocalMux I__4889 (
            .O(N__30942),
            .I(N__30935));
    Span4Mux_v I__4888 (
            .O(N__30939),
            .I(N__30932));
    InMux I__4887 (
            .O(N__30938),
            .I(N__30929));
    Odrv4 I__4886 (
            .O(N__30935),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    Odrv4 I__4885 (
            .O(N__30932),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    LocalMux I__4884 (
            .O(N__30929),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ));
    CascadeMux I__4883 (
            .O(N__30922),
            .I(N__30919));
    InMux I__4882 (
            .O(N__30919),
            .I(N__30916));
    LocalMux I__4881 (
            .O(N__30916),
            .I(\phase_controller_inst2.stoper_hc.un6_running_lt22 ));
    InMux I__4880 (
            .O(N__30913),
            .I(N__30910));
    LocalMux I__4879 (
            .O(N__30910),
            .I(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ));
    CascadeMux I__4878 (
            .O(N__30907),
            .I(N__30904));
    InMux I__4877 (
            .O(N__30904),
            .I(N__30901));
    LocalMux I__4876 (
            .O(N__30901),
            .I(\phase_controller_inst2.stoper_hc.counter_i_13 ));
    CascadeMux I__4875 (
            .O(N__30898),
            .I(N__30895));
    InMux I__4874 (
            .O(N__30895),
            .I(N__30892));
    LocalMux I__4873 (
            .O(N__30892),
            .I(N__30889));
    Odrv4 I__4872 (
            .O(N__30889),
            .I(\phase_controller_inst2.stoper_hc.counter_i_14 ));
    CascadeMux I__4871 (
            .O(N__30886),
            .I(N__30883));
    InMux I__4870 (
            .O(N__30883),
            .I(N__30880));
    LocalMux I__4869 (
            .O(N__30880),
            .I(\phase_controller_inst2.stoper_hc.counter_i_15 ));
    CascadeMux I__4868 (
            .O(N__30877),
            .I(N__30874));
    InMux I__4867 (
            .O(N__30874),
            .I(N__30871));
    LocalMux I__4866 (
            .O(N__30871),
            .I(\phase_controller_inst2.stoper_hc.counter_i_5 ));
    CascadeMux I__4865 (
            .O(N__30868),
            .I(N__30865));
    InMux I__4864 (
            .O(N__30865),
            .I(N__30862));
    LocalMux I__4863 (
            .O(N__30862),
            .I(\phase_controller_inst2.stoper_hc.counter_i_6 ));
    CascadeMux I__4862 (
            .O(N__30859),
            .I(N__30856));
    InMux I__4861 (
            .O(N__30856),
            .I(N__30853));
    LocalMux I__4860 (
            .O(N__30853),
            .I(\phase_controller_inst2.stoper_hc.counter_i_7 ));
    InMux I__4859 (
            .O(N__30850),
            .I(N__30847));
    LocalMux I__4858 (
            .O(N__30847),
            .I(\phase_controller_inst2.stoper_hc.counter_i_8 ));
    CascadeMux I__4857 (
            .O(N__30844),
            .I(N__30841));
    InMux I__4856 (
            .O(N__30841),
            .I(N__30838));
    LocalMux I__4855 (
            .O(N__30838),
            .I(\phase_controller_inst2.stoper_hc.counter_i_9 ));
    CascadeMux I__4854 (
            .O(N__30835),
            .I(N__30832));
    InMux I__4853 (
            .O(N__30832),
            .I(N__30829));
    LocalMux I__4852 (
            .O(N__30829),
            .I(\phase_controller_inst2.stoper_hc.counter_i_10 ));
    InMux I__4851 (
            .O(N__30826),
            .I(N__30823));
    LocalMux I__4850 (
            .O(N__30823),
            .I(\phase_controller_inst2.stoper_hc.counter_i_11 ));
    CascadeMux I__4849 (
            .O(N__30820),
            .I(N__30817));
    InMux I__4848 (
            .O(N__30817),
            .I(N__30814));
    LocalMux I__4847 (
            .O(N__30814),
            .I(N__30811));
    Odrv4 I__4846 (
            .O(N__30811),
            .I(\phase_controller_inst2.stoper_hc.counter_i_12 ));
    InMux I__4845 (
            .O(N__30808),
            .I(N__30805));
    LocalMux I__4844 (
            .O(N__30805),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ));
    InMux I__4843 (
            .O(N__30802),
            .I(N__30799));
    LocalMux I__4842 (
            .O(N__30799),
            .I(N__30796));
    Odrv4 I__4841 (
            .O(N__30796),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ));
    InMux I__4840 (
            .O(N__30793),
            .I(N__30790));
    LocalMux I__4839 (
            .O(N__30790),
            .I(N__30787));
    Span4Mux_h I__4838 (
            .O(N__30787),
            .I(N__30784));
    Sp12to4 I__4837 (
            .O(N__30784),
            .I(N__30781));
    Span12Mux_s6_v I__4836 (
            .O(N__30781),
            .I(N__30778));
    Odrv12 I__4835 (
            .O(N__30778),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_15 ));
    InMux I__4834 (
            .O(N__30775),
            .I(N__30761));
    CascadeMux I__4833 (
            .O(N__30774),
            .I(N__30758));
    CascadeMux I__4832 (
            .O(N__30773),
            .I(N__30755));
    CascadeMux I__4831 (
            .O(N__30772),
            .I(N__30752));
    CascadeMux I__4830 (
            .O(N__30771),
            .I(N__30749));
    CascadeMux I__4829 (
            .O(N__30770),
            .I(N__30746));
    CascadeMux I__4828 (
            .O(N__30769),
            .I(N__30743));
    CascadeMux I__4827 (
            .O(N__30768),
            .I(N__30740));
    CascadeMux I__4826 (
            .O(N__30767),
            .I(N__30737));
    CascadeMux I__4825 (
            .O(N__30766),
            .I(N__30734));
    CascadeMux I__4824 (
            .O(N__30765),
            .I(N__30731));
    CascadeMux I__4823 (
            .O(N__30764),
            .I(N__30728));
    LocalMux I__4822 (
            .O(N__30761),
            .I(N__30725));
    InMux I__4821 (
            .O(N__30758),
            .I(N__30718));
    InMux I__4820 (
            .O(N__30755),
            .I(N__30718));
    InMux I__4819 (
            .O(N__30752),
            .I(N__30718));
    InMux I__4818 (
            .O(N__30749),
            .I(N__30709));
    InMux I__4817 (
            .O(N__30746),
            .I(N__30709));
    InMux I__4816 (
            .O(N__30743),
            .I(N__30709));
    InMux I__4815 (
            .O(N__30740),
            .I(N__30709));
    InMux I__4814 (
            .O(N__30737),
            .I(N__30704));
    InMux I__4813 (
            .O(N__30734),
            .I(N__30704));
    InMux I__4812 (
            .O(N__30731),
            .I(N__30699));
    InMux I__4811 (
            .O(N__30728),
            .I(N__30699));
    Span4Mux_v I__4810 (
            .O(N__30725),
            .I(N__30696));
    LocalMux I__4809 (
            .O(N__30718),
            .I(N__30687));
    LocalMux I__4808 (
            .O(N__30709),
            .I(N__30687));
    LocalMux I__4807 (
            .O(N__30704),
            .I(N__30687));
    LocalMux I__4806 (
            .O(N__30699),
            .I(N__30687));
    Span4Mux_v I__4805 (
            .O(N__30696),
            .I(N__30684));
    Span4Mux_v I__4804 (
            .O(N__30687),
            .I(N__30681));
    Sp12to4 I__4803 (
            .O(N__30684),
            .I(N__30676));
    Sp12to4 I__4802 (
            .O(N__30681),
            .I(N__30676));
    Span12Mux_h I__4801 (
            .O(N__30676),
            .I(N__30673));
    Odrv12 I__4800 (
            .O(N__30673),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_19 ));
    CascadeMux I__4799 (
            .O(N__30670),
            .I(N__30667));
    InMux I__4798 (
            .O(N__30667),
            .I(N__30664));
    LocalMux I__4797 (
            .O(N__30664),
            .I(N__30661));
    Odrv4 I__4796 (
            .O(N__30661),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30 ));
    CascadeMux I__4795 (
            .O(N__30658),
            .I(N__30655));
    InMux I__4794 (
            .O(N__30655),
            .I(N__30652));
    LocalMux I__4793 (
            .O(N__30652),
            .I(\phase_controller_inst2.stoper_hc.counter_i_0 ));
    CascadeMux I__4792 (
            .O(N__30649),
            .I(N__30646));
    InMux I__4791 (
            .O(N__30646),
            .I(N__30643));
    LocalMux I__4790 (
            .O(N__30643),
            .I(\phase_controller_inst2.stoper_hc.counter_i_1 ));
    CascadeMux I__4789 (
            .O(N__30640),
            .I(N__30637));
    InMux I__4788 (
            .O(N__30637),
            .I(N__30634));
    LocalMux I__4787 (
            .O(N__30634),
            .I(N__30631));
    Odrv4 I__4786 (
            .O(N__30631),
            .I(\phase_controller_inst2.stoper_hc.counter_i_2 ));
    CascadeMux I__4785 (
            .O(N__30628),
            .I(N__30625));
    InMux I__4784 (
            .O(N__30625),
            .I(N__30622));
    LocalMux I__4783 (
            .O(N__30622),
            .I(\phase_controller_inst2.stoper_hc.counter_i_3 ));
    CascadeMux I__4782 (
            .O(N__30619),
            .I(N__30616));
    InMux I__4781 (
            .O(N__30616),
            .I(N__30613));
    LocalMux I__4780 (
            .O(N__30613),
            .I(N__30610));
    Odrv4 I__4779 (
            .O(N__30610),
            .I(\phase_controller_inst2.stoper_hc.counter_i_4 ));
    InMux I__4778 (
            .O(N__30607),
            .I(N__30604));
    LocalMux I__4777 (
            .O(N__30604),
            .I(N__30601));
    Odrv4 I__4776 (
            .O(N__30601),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ));
    InMux I__4775 (
            .O(N__30598),
            .I(N__30595));
    LocalMux I__4774 (
            .O(N__30595),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ));
    InMux I__4773 (
            .O(N__30592),
            .I(N__30589));
    LocalMux I__4772 (
            .O(N__30589),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ));
    InMux I__4771 (
            .O(N__30586),
            .I(N__30583));
    LocalMux I__4770 (
            .O(N__30583),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ));
    InMux I__4769 (
            .O(N__30580),
            .I(N__30577));
    LocalMux I__4768 (
            .O(N__30577),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ));
    InMux I__4767 (
            .O(N__30574),
            .I(N__30571));
    LocalMux I__4766 (
            .O(N__30571),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ));
    InMux I__4765 (
            .O(N__30568),
            .I(N__30565));
    LocalMux I__4764 (
            .O(N__30565),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ));
    InMux I__4763 (
            .O(N__30562),
            .I(N__30559));
    LocalMux I__4762 (
            .O(N__30559),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ));
    InMux I__4761 (
            .O(N__30556),
            .I(N__30553));
    LocalMux I__4760 (
            .O(N__30553),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ));
    InMux I__4759 (
            .O(N__30550),
            .I(N__30547));
    LocalMux I__4758 (
            .O(N__30547),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ));
    InMux I__4757 (
            .O(N__30544),
            .I(N__30541));
    LocalMux I__4756 (
            .O(N__30541),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ));
    InMux I__4755 (
            .O(N__30538),
            .I(N__30535));
    LocalMux I__4754 (
            .O(N__30535),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ));
    InMux I__4753 (
            .O(N__30532),
            .I(N__30529));
    LocalMux I__4752 (
            .O(N__30529),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ));
    InMux I__4751 (
            .O(N__30526),
            .I(N__30523));
    LocalMux I__4750 (
            .O(N__30523),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ));
    InMux I__4749 (
            .O(N__30520),
            .I(N__30517));
    LocalMux I__4748 (
            .O(N__30517),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ));
    InMux I__4747 (
            .O(N__30514),
            .I(N__30511));
    LocalMux I__4746 (
            .O(N__30511),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ));
    InMux I__4745 (
            .O(N__30508),
            .I(N__30505));
    LocalMux I__4744 (
            .O(N__30505),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ));
    InMux I__4743 (
            .O(N__30502),
            .I(bfn_10_17_0_));
    IoInMux I__4742 (
            .O(N__30499),
            .I(N__30496));
    LocalMux I__4741 (
            .O(N__30496),
            .I(N__30493));
    Span4Mux_s2_v I__4740 (
            .O(N__30493),
            .I(N__30490));
    Span4Mux_h I__4739 (
            .O(N__30490),
            .I(N__30487));
    Span4Mux_v I__4738 (
            .O(N__30487),
            .I(N__30484));
    Span4Mux_v I__4737 (
            .O(N__30484),
            .I(N__30481));
    Odrv4 I__4736 (
            .O(N__30481),
            .I(\phase_controller_inst1.stoper_tr.un2_start_0 ));
    InMux I__4735 (
            .O(N__30478),
            .I(N__30475));
    LocalMux I__4734 (
            .O(N__30475),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ));
    InMux I__4733 (
            .O(N__30472),
            .I(N__30469));
    LocalMux I__4732 (
            .O(N__30469),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ));
    CascadeMux I__4731 (
            .O(N__30466),
            .I(\current_shift_inst.PI_CTRL.N_44_cascade_ ));
    InMux I__4730 (
            .O(N__30463),
            .I(N__30460));
    LocalMux I__4729 (
            .O(N__30460),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ));
    CascadeMux I__4728 (
            .O(N__30457),
            .I(\current_shift_inst.PI_CTRL.un3_enable_0_cascade_ ));
    InMux I__4727 (
            .O(N__30454),
            .I(N__30451));
    LocalMux I__4726 (
            .O(N__30451),
            .I(N__30448));
    Span4Mux_h I__4725 (
            .O(N__30448),
            .I(N__30445));
    Span4Mux_h I__4724 (
            .O(N__30445),
            .I(N__30442));
    Odrv4 I__4723 (
            .O(N__30442),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ));
    CascadeMux I__4722 (
            .O(N__30439),
            .I(N__30436));
    InMux I__4721 (
            .O(N__30436),
            .I(N__30433));
    LocalMux I__4720 (
            .O(N__30433),
            .I(N__30430));
    Span4Mux_h I__4719 (
            .O(N__30430),
            .I(N__30427));
    Span4Mux_h I__4718 (
            .O(N__30427),
            .I(N__30424));
    Odrv4 I__4717 (
            .O(N__30424),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt16 ));
    InMux I__4716 (
            .O(N__30421),
            .I(N__30418));
    LocalMux I__4715 (
            .O(N__30418),
            .I(N__30415));
    Span4Mux_h I__4714 (
            .O(N__30415),
            .I(N__30412));
    Span4Mux_h I__4713 (
            .O(N__30412),
            .I(N__30409));
    Odrv4 I__4712 (
            .O(N__30409),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ));
    CascadeMux I__4711 (
            .O(N__30406),
            .I(N__30403));
    InMux I__4710 (
            .O(N__30403),
            .I(N__30400));
    LocalMux I__4709 (
            .O(N__30400),
            .I(N__30397));
    Span4Mux_v I__4708 (
            .O(N__30397),
            .I(N__30394));
    Span4Mux_h I__4707 (
            .O(N__30394),
            .I(N__30391));
    Odrv4 I__4706 (
            .O(N__30391),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt18 ));
    InMux I__4705 (
            .O(N__30388),
            .I(N__30385));
    LocalMux I__4704 (
            .O(N__30385),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ));
    CascadeMux I__4703 (
            .O(N__30382),
            .I(N__30379));
    InMux I__4702 (
            .O(N__30379),
            .I(N__30376));
    LocalMux I__4701 (
            .O(N__30376),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt24 ));
    InMux I__4700 (
            .O(N__30373),
            .I(N__30370));
    LocalMux I__4699 (
            .O(N__30370),
            .I(\phase_controller_inst1.stoper_tr.un6_running_lt26 ));
    CascadeMux I__4698 (
            .O(N__30367),
            .I(N__30364));
    InMux I__4697 (
            .O(N__30364),
            .I(N__30361));
    LocalMux I__4696 (
            .O(N__30361),
            .I(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ));
    InMux I__4695 (
            .O(N__30358),
            .I(N__30355));
    LocalMux I__4694 (
            .O(N__30355),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ));
    CascadeMux I__4693 (
            .O(N__30352),
            .I(N__30349));
    InMux I__4692 (
            .O(N__30349),
            .I(N__30346));
    LocalMux I__4691 (
            .O(N__30346),
            .I(N__30343));
    Odrv4 I__4690 (
            .O(N__30343),
            .I(\phase_controller_inst1.stoper_tr.counter_i_7 ));
    InMux I__4689 (
            .O(N__30340),
            .I(N__30337));
    LocalMux I__4688 (
            .O(N__30337),
            .I(\phase_controller_inst1.stoper_tr.counter_i_8 ));
    CascadeMux I__4687 (
            .O(N__30334),
            .I(N__30331));
    InMux I__4686 (
            .O(N__30331),
            .I(N__30328));
    LocalMux I__4685 (
            .O(N__30328),
            .I(\phase_controller_inst1.stoper_tr.counter_i_9 ));
    InMux I__4684 (
            .O(N__30325),
            .I(N__30322));
    LocalMux I__4683 (
            .O(N__30322),
            .I(\phase_controller_inst1.stoper_tr.counter_i_10 ));
    CascadeMux I__4682 (
            .O(N__30319),
            .I(N__30316));
    InMux I__4681 (
            .O(N__30316),
            .I(N__30313));
    LocalMux I__4680 (
            .O(N__30313),
            .I(\phase_controller_inst1.stoper_tr.counter_i_11 ));
    CascadeMux I__4679 (
            .O(N__30310),
            .I(N__30307));
    InMux I__4678 (
            .O(N__30307),
            .I(N__30304));
    LocalMux I__4677 (
            .O(N__30304),
            .I(\phase_controller_inst1.stoper_tr.counter_i_12 ));
    InMux I__4676 (
            .O(N__30301),
            .I(N__30298));
    LocalMux I__4675 (
            .O(N__30298),
            .I(N__30295));
    Odrv12 I__4674 (
            .O(N__30295),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ));
    CascadeMux I__4673 (
            .O(N__30292),
            .I(N__30289));
    InMux I__4672 (
            .O(N__30289),
            .I(N__30286));
    LocalMux I__4671 (
            .O(N__30286),
            .I(\phase_controller_inst1.stoper_tr.counter_i_13 ));
    CascadeMux I__4670 (
            .O(N__30283),
            .I(N__30280));
    InMux I__4669 (
            .O(N__30280),
            .I(N__30277));
    LocalMux I__4668 (
            .O(N__30277),
            .I(\phase_controller_inst1.stoper_tr.counter_i_14 ));
    CascadeMux I__4667 (
            .O(N__30274),
            .I(N__30271));
    InMux I__4666 (
            .O(N__30271),
            .I(N__30268));
    LocalMux I__4665 (
            .O(N__30268),
            .I(\phase_controller_inst1.stoper_tr.counter_i_15 ));
    InMux I__4664 (
            .O(N__30265),
            .I(N__30261));
    InMux I__4663 (
            .O(N__30264),
            .I(N__30258));
    LocalMux I__4662 (
            .O(N__30261),
            .I(N__30255));
    LocalMux I__4661 (
            .O(N__30258),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_3));
    Odrv4 I__4660 (
            .O(N__30255),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_3));
    CascadeMux I__4659 (
            .O(N__30250),
            .I(N__30247));
    InMux I__4658 (
            .O(N__30247),
            .I(N__30244));
    LocalMux I__4657 (
            .O(N__30244),
            .I(\phase_controller_inst1.stoper_tr.counter_i_0 ));
    InMux I__4656 (
            .O(N__30241),
            .I(N__30238));
    LocalMux I__4655 (
            .O(N__30238),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ));
    CascadeMux I__4654 (
            .O(N__30235),
            .I(N__30232));
    InMux I__4653 (
            .O(N__30232),
            .I(N__30229));
    LocalMux I__4652 (
            .O(N__30229),
            .I(\phase_controller_inst1.stoper_tr.counter_i_1 ));
    CascadeMux I__4651 (
            .O(N__30226),
            .I(N__30223));
    InMux I__4650 (
            .O(N__30223),
            .I(N__30220));
    LocalMux I__4649 (
            .O(N__30220),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ));
    InMux I__4648 (
            .O(N__30217),
            .I(N__30214));
    LocalMux I__4647 (
            .O(N__30214),
            .I(\phase_controller_inst1.stoper_tr.counter_i_2 ));
    InMux I__4646 (
            .O(N__30211),
            .I(N__30208));
    LocalMux I__4645 (
            .O(N__30208),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ));
    CascadeMux I__4644 (
            .O(N__30205),
            .I(N__30202));
    InMux I__4643 (
            .O(N__30202),
            .I(N__30199));
    LocalMux I__4642 (
            .O(N__30199),
            .I(\phase_controller_inst1.stoper_tr.counter_i_3 ));
    InMux I__4641 (
            .O(N__30196),
            .I(N__30193));
    LocalMux I__4640 (
            .O(N__30193),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ));
    CascadeMux I__4639 (
            .O(N__30190),
            .I(N__30187));
    InMux I__4638 (
            .O(N__30187),
            .I(N__30184));
    LocalMux I__4637 (
            .O(N__30184),
            .I(\phase_controller_inst1.stoper_tr.counter_i_4 ));
    InMux I__4636 (
            .O(N__30181),
            .I(N__30178));
    LocalMux I__4635 (
            .O(N__30178),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ));
    CascadeMux I__4634 (
            .O(N__30175),
            .I(N__30172));
    InMux I__4633 (
            .O(N__30172),
            .I(N__30169));
    LocalMux I__4632 (
            .O(N__30169),
            .I(\phase_controller_inst1.stoper_tr.counter_i_5 ));
    InMux I__4631 (
            .O(N__30166),
            .I(N__30163));
    LocalMux I__4630 (
            .O(N__30163),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ));
    CascadeMux I__4629 (
            .O(N__30160),
            .I(N__30157));
    InMux I__4628 (
            .O(N__30157),
            .I(N__30154));
    LocalMux I__4627 (
            .O(N__30154),
            .I(\phase_controller_inst1.stoper_tr.counter_i_6 ));
    CascadeMux I__4626 (
            .O(N__30151),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_));
    InMux I__4625 (
            .O(N__30148),
            .I(N__30145));
    LocalMux I__4624 (
            .O(N__30145),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ));
    InMux I__4623 (
            .O(N__30142),
            .I(N__30138));
    InMux I__4622 (
            .O(N__30141),
            .I(N__30135));
    LocalMux I__4621 (
            .O(N__30138),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    LocalMux I__4620 (
            .O(N__30135),
            .I(elapsed_time_ns_1_RNI3EPBB_0_25));
    InMux I__4619 (
            .O(N__30130),
            .I(N__30127));
    LocalMux I__4618 (
            .O(N__30127),
            .I(N__30124));
    Odrv4 I__4617 (
            .O(N__30124),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ));
    InMux I__4616 (
            .O(N__30121),
            .I(N__30117));
    InMux I__4615 (
            .O(N__30120),
            .I(N__30114));
    LocalMux I__4614 (
            .O(N__30117),
            .I(N__30111));
    LocalMux I__4613 (
            .O(N__30114),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_1));
    Odrv4 I__4612 (
            .O(N__30111),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_1));
    InMux I__4611 (
            .O(N__30106),
            .I(N__30102));
    InMux I__4610 (
            .O(N__30105),
            .I(N__30099));
    LocalMux I__4609 (
            .O(N__30102),
            .I(N__30096));
    LocalMux I__4608 (
            .O(N__30099),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_6));
    Odrv4 I__4607 (
            .O(N__30096),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_6));
    InMux I__4606 (
            .O(N__30091),
            .I(N__30087));
    InMux I__4605 (
            .O(N__30090),
            .I(N__30084));
    LocalMux I__4604 (
            .O(N__30087),
            .I(N__30081));
    LocalMux I__4603 (
            .O(N__30084),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_5));
    Odrv4 I__4602 (
            .O(N__30081),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_5));
    InMux I__4601 (
            .O(N__30076),
            .I(N__30073));
    LocalMux I__4600 (
            .O(N__30073),
            .I(N__30070));
    Span4Mux_h I__4599 (
            .O(N__30070),
            .I(N__30066));
    InMux I__4598 (
            .O(N__30069),
            .I(N__30063));
    Odrv4 I__4597 (
            .O(N__30066),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_13));
    LocalMux I__4596 (
            .O(N__30063),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_13));
    InMux I__4595 (
            .O(N__30058),
            .I(N__30054));
    InMux I__4594 (
            .O(N__30057),
            .I(N__30051));
    LocalMux I__4593 (
            .O(N__30054),
            .I(N__30048));
    LocalMux I__4592 (
            .O(N__30051),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_7));
    Odrv4 I__4591 (
            .O(N__30048),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_7));
    InMux I__4590 (
            .O(N__30043),
            .I(N__30039));
    InMux I__4589 (
            .O(N__30042),
            .I(N__30036));
    LocalMux I__4588 (
            .O(N__30039),
            .I(N__30033));
    LocalMux I__4587 (
            .O(N__30036),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_4));
    Odrv4 I__4586 (
            .O(N__30033),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_4));
    InMux I__4585 (
            .O(N__30028),
            .I(N__30025));
    LocalMux I__4584 (
            .O(N__30025),
            .I(N__30021));
    InMux I__4583 (
            .O(N__30024),
            .I(N__30018));
    Span4Mux_v I__4582 (
            .O(N__30021),
            .I(N__30013));
    LocalMux I__4581 (
            .O(N__30018),
            .I(N__30013));
    Odrv4 I__4580 (
            .O(N__30013),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_2));
    InMux I__4579 (
            .O(N__30010),
            .I(N__30007));
    LocalMux I__4578 (
            .O(N__30007),
            .I(N__30004));
    Span4Mux_v I__4577 (
            .O(N__30004),
            .I(N__30000));
    InMux I__4576 (
            .O(N__30003),
            .I(N__29997));
    Odrv4 I__4575 (
            .O(N__30000),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    LocalMux I__4574 (
            .O(N__29997),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ));
    InMux I__4573 (
            .O(N__29992),
            .I(N__29989));
    LocalMux I__4572 (
            .O(N__29989),
            .I(N__29985));
    CascadeMux I__4571 (
            .O(N__29988),
            .I(N__29982));
    Span4Mux_h I__4570 (
            .O(N__29985),
            .I(N__29979));
    InMux I__4569 (
            .O(N__29982),
            .I(N__29976));
    Odrv4 I__4568 (
            .O(N__29979),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    LocalMux I__4567 (
            .O(N__29976),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ));
    InMux I__4566 (
            .O(N__29971),
            .I(N__29967));
    InMux I__4565 (
            .O(N__29970),
            .I(N__29964));
    LocalMux I__4564 (
            .O(N__29967),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    LocalMux I__4563 (
            .O(N__29964),
            .I(elapsed_time_ns_1_RNIGF91B_0_4));
    InMux I__4562 (
            .O(N__29959),
            .I(N__29956));
    LocalMux I__4561 (
            .O(N__29956),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ));
    InMux I__4560 (
            .O(N__29953),
            .I(N__29949));
    InMux I__4559 (
            .O(N__29952),
            .I(N__29946));
    LocalMux I__4558 (
            .O(N__29949),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    LocalMux I__4557 (
            .O(N__29946),
            .I(elapsed_time_ns_1_RNI2DPBB_0_24));
    InMux I__4556 (
            .O(N__29941),
            .I(N__29938));
    LocalMux I__4555 (
            .O(N__29938),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ));
    InMux I__4554 (
            .O(N__29935),
            .I(N__29931));
    InMux I__4553 (
            .O(N__29934),
            .I(N__29928));
    LocalMux I__4552 (
            .O(N__29931),
            .I(N__29923));
    LocalMux I__4551 (
            .O(N__29928),
            .I(N__29923));
    Span4Mux_v I__4550 (
            .O(N__29923),
            .I(N__29920));
    Odrv4 I__4549 (
            .O(N__29920),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ));
    InMux I__4548 (
            .O(N__29917),
            .I(N__29914));
    LocalMux I__4547 (
            .O(N__29914),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8));
    CascadeMux I__4546 (
            .O(N__29911),
            .I(elapsed_time_ns_1_RNIKJ91B_0_8_cascade_));
    InMux I__4545 (
            .O(N__29908),
            .I(N__29905));
    LocalMux I__4544 (
            .O(N__29905),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ));
    InMux I__4543 (
            .O(N__29902),
            .I(N__29898));
    InMux I__4542 (
            .O(N__29901),
            .I(N__29895));
    LocalMux I__4541 (
            .O(N__29898),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    LocalMux I__4540 (
            .O(N__29895),
            .I(elapsed_time_ns_1_RNI0BPBB_0_22));
    InMux I__4539 (
            .O(N__29890),
            .I(N__29887));
    LocalMux I__4538 (
            .O(N__29887),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ));
    InMux I__4537 (
            .O(N__29884),
            .I(N__29881));
    LocalMux I__4536 (
            .O(N__29881),
            .I(N__29877));
    CascadeMux I__4535 (
            .O(N__29880),
            .I(N__29874));
    Span4Mux_h I__4534 (
            .O(N__29877),
            .I(N__29871));
    InMux I__4533 (
            .O(N__29874),
            .I(N__29868));
    Odrv4 I__4532 (
            .O(N__29871),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    LocalMux I__4531 (
            .O(N__29868),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ));
    InMux I__4530 (
            .O(N__29863),
            .I(N__29860));
    LocalMux I__4529 (
            .O(N__29860),
            .I(elapsed_time_ns_1_RNIU8PBB_0_20));
    InMux I__4528 (
            .O(N__29857),
            .I(N__29854));
    LocalMux I__4527 (
            .O(N__29854),
            .I(N__29851));
    Span4Mux_h I__4526 (
            .O(N__29851),
            .I(N__29847));
    InMux I__4525 (
            .O(N__29850),
            .I(N__29844));
    Odrv4 I__4524 (
            .O(N__29847),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    LocalMux I__4523 (
            .O(N__29844),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ));
    InMux I__4522 (
            .O(N__29839),
            .I(N__29836));
    LocalMux I__4521 (
            .O(N__29836),
            .I(N__29832));
    CascadeMux I__4520 (
            .O(N__29835),
            .I(N__29829));
    Span4Mux_v I__4519 (
            .O(N__29832),
            .I(N__29825));
    InMux I__4518 (
            .O(N__29829),
            .I(N__29822));
    InMux I__4517 (
            .O(N__29828),
            .I(N__29819));
    Odrv4 I__4516 (
            .O(N__29825),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__4515 (
            .O(N__29822),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    LocalMux I__4514 (
            .O(N__29819),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ));
    CascadeMux I__4513 (
            .O(N__29812),
            .I(N__29809));
    InMux I__4512 (
            .O(N__29809),
            .I(N__29805));
    InMux I__4511 (
            .O(N__29808),
            .I(N__29802));
    LocalMux I__4510 (
            .O(N__29805),
            .I(N__29799));
    LocalMux I__4509 (
            .O(N__29802),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    Odrv4 I__4508 (
            .O(N__29799),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ));
    InMux I__4507 (
            .O(N__29794),
            .I(N__29791));
    LocalMux I__4506 (
            .O(N__29791),
            .I(N__29787));
    CascadeMux I__4505 (
            .O(N__29790),
            .I(N__29784));
    Span4Mux_v I__4504 (
            .O(N__29787),
            .I(N__29780));
    InMux I__4503 (
            .O(N__29784),
            .I(N__29777));
    InMux I__4502 (
            .O(N__29783),
            .I(N__29774));
    Odrv4 I__4501 (
            .O(N__29780),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__4500 (
            .O(N__29777),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    LocalMux I__4499 (
            .O(N__29774),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ));
    InMux I__4498 (
            .O(N__29767),
            .I(N__29763));
    InMux I__4497 (
            .O(N__29766),
            .I(N__29760));
    LocalMux I__4496 (
            .O(N__29763),
            .I(N__29757));
    LocalMux I__4495 (
            .O(N__29760),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    Odrv4 I__4494 (
            .O(N__29757),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ));
    InMux I__4493 (
            .O(N__29752),
            .I(N__29748));
    InMux I__4492 (
            .O(N__29751),
            .I(N__29745));
    LocalMux I__4491 (
            .O(N__29748),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    LocalMux I__4490 (
            .O(N__29745),
            .I(elapsed_time_ns_1_RNIED91B_0_2));
    InMux I__4489 (
            .O(N__29740),
            .I(N__29736));
    InMux I__4488 (
            .O(N__29739),
            .I(N__29733));
    LocalMux I__4487 (
            .O(N__29736),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    LocalMux I__4486 (
            .O(N__29733),
            .I(elapsed_time_ns_1_RNIFE91B_0_3));
    InMux I__4485 (
            .O(N__29728),
            .I(N__29725));
    LocalMux I__4484 (
            .O(N__29725),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ));
    InMux I__4483 (
            .O(N__29722),
            .I(N__29719));
    LocalMux I__4482 (
            .O(N__29719),
            .I(N__29716));
    Span4Mux_h I__4481 (
            .O(N__29716),
            .I(N__29712));
    InMux I__4480 (
            .O(N__29715),
            .I(N__29709));
    Odrv4 I__4479 (
            .O(N__29712),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    LocalMux I__4478 (
            .O(N__29709),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ));
    InMux I__4477 (
            .O(N__29704),
            .I(N__29701));
    LocalMux I__4476 (
            .O(N__29701),
            .I(N__29698));
    Span4Mux_h I__4475 (
            .O(N__29698),
            .I(N__29694));
    InMux I__4474 (
            .O(N__29697),
            .I(N__29691));
    Odrv4 I__4473 (
            .O(N__29694),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    LocalMux I__4472 (
            .O(N__29691),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ));
    InMux I__4471 (
            .O(N__29686),
            .I(N__29683));
    LocalMux I__4470 (
            .O(N__29683),
            .I(elapsed_time_ns_1_RNIIH91B_0_6));
    CascadeMux I__4469 (
            .O(N__29680),
            .I(elapsed_time_ns_1_RNIIH91B_0_6_cascade_));
    InMux I__4468 (
            .O(N__29677),
            .I(N__29674));
    LocalMux I__4467 (
            .O(N__29674),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ));
    InMux I__4466 (
            .O(N__29671),
            .I(N__29668));
    LocalMux I__4465 (
            .O(N__29668),
            .I(N__29665));
    Span4Mux_h I__4464 (
            .O(N__29665),
            .I(N__29661));
    InMux I__4463 (
            .O(N__29664),
            .I(N__29658));
    Odrv4 I__4462 (
            .O(N__29661),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    LocalMux I__4461 (
            .O(N__29658),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ));
    InMux I__4460 (
            .O(N__29653),
            .I(N__29648));
    InMux I__4459 (
            .O(N__29652),
            .I(N__29643));
    InMux I__4458 (
            .O(N__29651),
            .I(N__29643));
    LocalMux I__4457 (
            .O(N__29648),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    LocalMux I__4456 (
            .O(N__29643),
            .I(\phase_controller_inst2.stoper_tr.runningZ0 ));
    InMux I__4455 (
            .O(N__29638),
            .I(N__29635));
    LocalMux I__4454 (
            .O(N__29635),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ));
    CascadeMux I__4453 (
            .O(N__29632),
            .I(N__29629));
    InMux I__4452 (
            .O(N__29629),
            .I(N__29625));
    InMux I__4451 (
            .O(N__29628),
            .I(N__29622));
    LocalMux I__4450 (
            .O(N__29625),
            .I(N__29619));
    LocalMux I__4449 (
            .O(N__29622),
            .I(N__29616));
    Span4Mux_v I__4448 (
            .O(N__29619),
            .I(N__29613));
    Odrv4 I__4447 (
            .O(N__29616),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    Odrv4 I__4446 (
            .O(N__29613),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ));
    InMux I__4445 (
            .O(N__29608),
            .I(N__29605));
    LocalMux I__4444 (
            .O(N__29605),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ));
    InMux I__4443 (
            .O(N__29602),
            .I(N__29599));
    LocalMux I__4442 (
            .O(N__29599),
            .I(N__29595));
    InMux I__4441 (
            .O(N__29598),
            .I(N__29592));
    Span4Mux_h I__4440 (
            .O(N__29595),
            .I(N__29589));
    LocalMux I__4439 (
            .O(N__29592),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    Odrv4 I__4438 (
            .O(N__29589),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ));
    InMux I__4437 (
            .O(N__29584),
            .I(N__29581));
    LocalMux I__4436 (
            .O(N__29581),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ));
    CascadeMux I__4435 (
            .O(N__29578),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ));
    InMux I__4434 (
            .O(N__29575),
            .I(N__29572));
    LocalMux I__4433 (
            .O(N__29572),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ));
    CascadeMux I__4432 (
            .O(N__29569),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ));
    InMux I__4431 (
            .O(N__29566),
            .I(N__29562));
    InMux I__4430 (
            .O(N__29565),
            .I(N__29559));
    LocalMux I__4429 (
            .O(N__29562),
            .I(N__29556));
    LocalMux I__4428 (
            .O(N__29559),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    Odrv4 I__4427 (
            .O(N__29556),
            .I(elapsed_time_ns_1_RNIDC91B_0_1));
    InMux I__4426 (
            .O(N__29551),
            .I(N__29548));
    LocalMux I__4425 (
            .O(N__29548),
            .I(N__29545));
    Span4Mux_v I__4424 (
            .O(N__29545),
            .I(N__29542));
    Odrv4 I__4423 (
            .O(N__29542),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ));
    InMux I__4422 (
            .O(N__29539),
            .I(N__29536));
    LocalMux I__4421 (
            .O(N__29536),
            .I(N__29532));
    InMux I__4420 (
            .O(N__29535),
            .I(N__29529));
    Odrv4 I__4419 (
            .O(N__29532),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    LocalMux I__4418 (
            .O(N__29529),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ));
    InMux I__4417 (
            .O(N__29524),
            .I(N__29518));
    InMux I__4416 (
            .O(N__29523),
            .I(N__29518));
    LocalMux I__4415 (
            .O(N__29518),
            .I(elapsed_time_ns_1_RNI4EOBB_0_17));
    InMux I__4414 (
            .O(N__29515),
            .I(N__29512));
    LocalMux I__4413 (
            .O(N__29512),
            .I(N__29508));
    InMux I__4412 (
            .O(N__29511),
            .I(N__29505));
    Odrv4 I__4411 (
            .O(N__29508),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    LocalMux I__4410 (
            .O(N__29505),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ));
    InMux I__4409 (
            .O(N__29500),
            .I(N__29497));
    LocalMux I__4408 (
            .O(N__29497),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11));
    CascadeMux I__4407 (
            .O(N__29494),
            .I(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_));
    InMux I__4406 (
            .O(N__29491),
            .I(N__29488));
    LocalMux I__4405 (
            .O(N__29488),
            .I(N__29485));
    Odrv4 I__4404 (
            .O(N__29485),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ));
    IoInMux I__4403 (
            .O(N__29482),
            .I(N__29479));
    LocalMux I__4402 (
            .O(N__29479),
            .I(N__29476));
    Span4Mux_s0_v I__4401 (
            .O(N__29476),
            .I(N__29473));
    Span4Mux_v I__4400 (
            .O(N__29473),
            .I(N__29470));
    Odrv4 I__4399 (
            .O(N__29470),
            .I(s4_phy_c));
    InMux I__4398 (
            .O(N__29467),
            .I(N__29462));
    InMux I__4397 (
            .O(N__29466),
            .I(N__29459));
    InMux I__4396 (
            .O(N__29465),
            .I(N__29456));
    LocalMux I__4395 (
            .O(N__29462),
            .I(N__29451));
    LocalMux I__4394 (
            .O(N__29459),
            .I(N__29451));
    LocalMux I__4393 (
            .O(N__29456),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    Odrv4 I__4392 (
            .O(N__29451),
            .I(\phase_controller_inst2.stoper_hc.runningZ0 ));
    InMux I__4391 (
            .O(N__29446),
            .I(N__29443));
    LocalMux I__4390 (
            .O(N__29443),
            .I(N__29438));
    InMux I__4389 (
            .O(N__29442),
            .I(N__29433));
    InMux I__4388 (
            .O(N__29441),
            .I(N__29433));
    Span4Mux_v I__4387 (
            .O(N__29438),
            .I(N__29428));
    LocalMux I__4386 (
            .O(N__29433),
            .I(N__29428));
    Span4Mux_h I__4385 (
            .O(N__29428),
            .I(N__29425));
    Span4Mux_v I__4384 (
            .O(N__29425),
            .I(N__29422));
    Odrv4 I__4383 (
            .O(N__29422),
            .I(il_min_comp2_c));
    InMux I__4382 (
            .O(N__29419),
            .I(N__29416));
    LocalMux I__4381 (
            .O(N__29416),
            .I(N__29413));
    Span4Mux_v I__4380 (
            .O(N__29413),
            .I(N__29410));
    Span4Mux_v I__4379 (
            .O(N__29410),
            .I(N__29406));
    CascadeMux I__4378 (
            .O(N__29409),
            .I(N__29401));
    Span4Mux_v I__4377 (
            .O(N__29406),
            .I(N__29398));
    InMux I__4376 (
            .O(N__29405),
            .I(N__29395));
    InMux I__4375 (
            .O(N__29404),
            .I(N__29390));
    InMux I__4374 (
            .O(N__29401),
            .I(N__29390));
    Span4Mux_v I__4373 (
            .O(N__29398),
            .I(N__29387));
    LocalMux I__4372 (
            .O(N__29395),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    LocalMux I__4371 (
            .O(N__29390),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    Odrv4 I__4370 (
            .O(N__29387),
            .I(\phase_controller_inst2.stateZ0Z_1 ));
    InMux I__4369 (
            .O(N__29380),
            .I(N__29377));
    LocalMux I__4368 (
            .O(N__29377),
            .I(N__29372));
    InMux I__4367 (
            .O(N__29376),
            .I(N__29367));
    InMux I__4366 (
            .O(N__29375),
            .I(N__29367));
    Span4Mux_h I__4365 (
            .O(N__29372),
            .I(N__29362));
    LocalMux I__4364 (
            .O(N__29367),
            .I(N__29362));
    Span4Mux_v I__4363 (
            .O(N__29362),
            .I(N__29359));
    IoSpan4Mux I__4362 (
            .O(N__29359),
            .I(N__29356));
    Odrv4 I__4361 (
            .O(N__29356),
            .I(il_max_comp2_c));
    CascadeMux I__4360 (
            .O(N__29353),
            .I(N__29350));
    InMux I__4359 (
            .O(N__29350),
            .I(N__29346));
    InMux I__4358 (
            .O(N__29349),
            .I(N__29343));
    LocalMux I__4357 (
            .O(N__29346),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    LocalMux I__4356 (
            .O(N__29343),
            .I(\phase_controller_inst2.stateZ0Z_0 ));
    CascadeMux I__4355 (
            .O(N__29338),
            .I(\phase_controller_inst2.state_ns_0_0_1_cascade_ ));
    InMux I__4354 (
            .O(N__29335),
            .I(N__29332));
    LocalMux I__4353 (
            .O(N__29332),
            .I(N__29328));
    CascadeMux I__4352 (
            .O(N__29331),
            .I(N__29324));
    Sp12to4 I__4351 (
            .O(N__29328),
            .I(N__29320));
    InMux I__4350 (
            .O(N__29327),
            .I(N__29315));
    InMux I__4349 (
            .O(N__29324),
            .I(N__29315));
    InMux I__4348 (
            .O(N__29323),
            .I(N__29312));
    Span12Mux_v I__4347 (
            .O(N__29320),
            .I(N__29309));
    LocalMux I__4346 (
            .O(N__29315),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    LocalMux I__4345 (
            .O(N__29312),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    Odrv12 I__4344 (
            .O(N__29309),
            .I(\phase_controller_inst2.stateZ0Z_3 ));
    CascadeMux I__4343 (
            .O(N__29302),
            .I(\phase_controller_inst2.stoper_tr.un4_start_0_cascade_ ));
    CascadeMux I__4342 (
            .O(N__29299),
            .I(N__29294));
    InMux I__4341 (
            .O(N__29298),
            .I(N__29291));
    InMux I__4340 (
            .O(N__29297),
            .I(N__29286));
    InMux I__4339 (
            .O(N__29294),
            .I(N__29286));
    LocalMux I__4338 (
            .O(N__29291),
            .I(\phase_controller_inst2.tr_time_passed ));
    LocalMux I__4337 (
            .O(N__29286),
            .I(\phase_controller_inst2.tr_time_passed ));
    IoInMux I__4336 (
            .O(N__29281),
            .I(N__29278));
    LocalMux I__4335 (
            .O(N__29278),
            .I(N__29275));
    Span12Mux_s6_v I__4334 (
            .O(N__29275),
            .I(N__29272));
    Odrv12 I__4333 (
            .O(N__29272),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0 ));
    InMux I__4332 (
            .O(N__29269),
            .I(N__29261));
    InMux I__4331 (
            .O(N__29268),
            .I(N__29258));
    InMux I__4330 (
            .O(N__29267),
            .I(N__29255));
    InMux I__4329 (
            .O(N__29266),
            .I(N__29248));
    InMux I__4328 (
            .O(N__29265),
            .I(N__29248));
    InMux I__4327 (
            .O(N__29264),
            .I(N__29248));
    LocalMux I__4326 (
            .O(N__29261),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__4325 (
            .O(N__29258),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__4324 (
            .O(N__29255),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    LocalMux I__4323 (
            .O(N__29248),
            .I(\phase_controller_inst2.start_timer_trZ0 ));
    InMux I__4322 (
            .O(N__29239),
            .I(N__29233));
    InMux I__4321 (
            .O(N__29238),
            .I(N__29233));
    LocalMux I__4320 (
            .O(N__29233),
            .I(N__29230));
    Span4Mux_v I__4319 (
            .O(N__29230),
            .I(N__29227));
    Span4Mux_v I__4318 (
            .O(N__29227),
            .I(N__29224));
    Span4Mux_v I__4317 (
            .O(N__29224),
            .I(N__29221));
    Span4Mux_h I__4316 (
            .O(N__29221),
            .I(N__29217));
    InMux I__4315 (
            .O(N__29220),
            .I(N__29214));
    Odrv4 I__4314 (
            .O(N__29217),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    LocalMux I__4313 (
            .O(N__29214),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ));
    CascadeMux I__4312 (
            .O(N__29209),
            .I(N__29206));
    InMux I__4311 (
            .O(N__29206),
            .I(N__29203));
    LocalMux I__4310 (
            .O(N__29203),
            .I(\current_shift_inst.PI_CTRL.integrator_1_30 ));
    InMux I__4309 (
            .O(N__29200),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ));
    InMux I__4308 (
            .O(N__29197),
            .I(N__29194));
    LocalMux I__4307 (
            .O(N__29194),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ));
    InMux I__4306 (
            .O(N__29191),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ));
    InMux I__4305 (
            .O(N__29188),
            .I(N__29185));
    LocalMux I__4304 (
            .O(N__29185),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ));
    InMux I__4303 (
            .O(N__29182),
            .I(N__29179));
    LocalMux I__4302 (
            .O(N__29179),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ));
    InMux I__4301 (
            .O(N__29176),
            .I(N__29173));
    LocalMux I__4300 (
            .O(N__29173),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ));
    InMux I__4299 (
            .O(N__29170),
            .I(N__29167));
    LocalMux I__4298 (
            .O(N__29167),
            .I(N__29164));
    Odrv4 I__4297 (
            .O(N__29164),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ));
    InMux I__4296 (
            .O(N__29161),
            .I(N__29158));
    LocalMux I__4295 (
            .O(N__29158),
            .I(N__29155));
    Odrv12 I__4294 (
            .O(N__29155),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ));
    InMux I__4293 (
            .O(N__29152),
            .I(N__29149));
    LocalMux I__4292 (
            .O(N__29149),
            .I(N__29146));
    Odrv12 I__4291 (
            .O(N__29146),
            .I(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ));
    IoInMux I__4290 (
            .O(N__29143),
            .I(N__29140));
    LocalMux I__4289 (
            .O(N__29140),
            .I(N__29137));
    Span4Mux_s3_v I__4288 (
            .O(N__29137),
            .I(N__29134));
    Odrv4 I__4287 (
            .O(N__29134),
            .I(s3_phy_c));
    CascadeMux I__4286 (
            .O(N__29131),
            .I(N__29128));
    InMux I__4285 (
            .O(N__29128),
            .I(N__29125));
    LocalMux I__4284 (
            .O(N__29125),
            .I(N__29122));
    Odrv4 I__4283 (
            .O(N__29122),
            .I(\current_shift_inst.PI_CTRL.integrator_1_21 ));
    InMux I__4282 (
            .O(N__29119),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ));
    InMux I__4281 (
            .O(N__29116),
            .I(N__29113));
    LocalMux I__4280 (
            .O(N__29113),
            .I(\current_shift_inst.PI_CTRL.integrator_1_22 ));
    InMux I__4279 (
            .O(N__29110),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ));
    CascadeMux I__4278 (
            .O(N__29107),
            .I(N__29104));
    InMux I__4277 (
            .O(N__29104),
            .I(N__29101));
    LocalMux I__4276 (
            .O(N__29101),
            .I(\current_shift_inst.PI_CTRL.integrator_1_23 ));
    InMux I__4275 (
            .O(N__29098),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ));
    CascadeMux I__4274 (
            .O(N__29095),
            .I(N__29092));
    InMux I__4273 (
            .O(N__29092),
            .I(N__29089));
    LocalMux I__4272 (
            .O(N__29089),
            .I(N__29086));
    Span4Mux_h I__4271 (
            .O(N__29086),
            .I(N__29083));
    Odrv4 I__4270 (
            .O(N__29083),
            .I(\current_shift_inst.PI_CTRL.integrator_1_24 ));
    InMux I__4269 (
            .O(N__29080),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ));
    CascadeMux I__4268 (
            .O(N__29077),
            .I(N__29074));
    InMux I__4267 (
            .O(N__29074),
            .I(N__29071));
    LocalMux I__4266 (
            .O(N__29071),
            .I(\current_shift_inst.PI_CTRL.integrator_1_25 ));
    InMux I__4265 (
            .O(N__29068),
            .I(bfn_9_21_0_));
    CascadeMux I__4264 (
            .O(N__29065),
            .I(N__29062));
    InMux I__4263 (
            .O(N__29062),
            .I(N__29059));
    LocalMux I__4262 (
            .O(N__29059),
            .I(\current_shift_inst.PI_CTRL.integrator_1_26 ));
    InMux I__4261 (
            .O(N__29056),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ));
    CascadeMux I__4260 (
            .O(N__29053),
            .I(N__29050));
    InMux I__4259 (
            .O(N__29050),
            .I(N__29047));
    LocalMux I__4258 (
            .O(N__29047),
            .I(\current_shift_inst.PI_CTRL.integrator_1_27 ));
    InMux I__4257 (
            .O(N__29044),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ));
    CascadeMux I__4256 (
            .O(N__29041),
            .I(N__29038));
    InMux I__4255 (
            .O(N__29038),
            .I(N__29035));
    LocalMux I__4254 (
            .O(N__29035),
            .I(N__29032));
    Odrv4 I__4253 (
            .O(N__29032),
            .I(\current_shift_inst.PI_CTRL.integrator_1_28 ));
    InMux I__4252 (
            .O(N__29029),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ));
    CascadeMux I__4251 (
            .O(N__29026),
            .I(N__29023));
    InMux I__4250 (
            .O(N__29023),
            .I(N__29020));
    LocalMux I__4249 (
            .O(N__29020),
            .I(\current_shift_inst.PI_CTRL.integrator_1_29 ));
    InMux I__4248 (
            .O(N__29017),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ));
    CascadeMux I__4247 (
            .O(N__29014),
            .I(N__29011));
    InMux I__4246 (
            .O(N__29011),
            .I(N__29008));
    LocalMux I__4245 (
            .O(N__29008),
            .I(N__29005));
    Span4Mux_v I__4244 (
            .O(N__29005),
            .I(N__29002));
    Sp12to4 I__4243 (
            .O(N__29002),
            .I(N__28999));
    Span12Mux_h I__4242 (
            .O(N__28999),
            .I(N__28996));
    Span12Mux_v I__4241 (
            .O(N__28996),
            .I(N__28993));
    Odrv12 I__4240 (
            .O(N__28993),
            .I(\current_shift_inst.PI_CTRL.integrator_1_13 ));
    InMux I__4239 (
            .O(N__28990),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ));
    CascadeMux I__4238 (
            .O(N__28987),
            .I(N__28984));
    InMux I__4237 (
            .O(N__28984),
            .I(N__28981));
    LocalMux I__4236 (
            .O(N__28981),
            .I(N__28978));
    Span4Mux_h I__4235 (
            .O(N__28978),
            .I(N__28975));
    Span4Mux_h I__4234 (
            .O(N__28975),
            .I(N__28972));
    Sp12to4 I__4233 (
            .O(N__28972),
            .I(N__28969));
    Span12Mux_v I__4232 (
            .O(N__28969),
            .I(N__28966));
    Odrv12 I__4231 (
            .O(N__28966),
            .I(\current_shift_inst.PI_CTRL.integrator_1_14 ));
    InMux I__4230 (
            .O(N__28963),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ));
    CascadeMux I__4229 (
            .O(N__28960),
            .I(N__28957));
    InMux I__4228 (
            .O(N__28957),
            .I(N__28954));
    LocalMux I__4227 (
            .O(N__28954),
            .I(N__28951));
    Span4Mux_v I__4226 (
            .O(N__28951),
            .I(N__28948));
    Sp12to4 I__4225 (
            .O(N__28948),
            .I(N__28945));
    Span12Mux_v I__4224 (
            .O(N__28945),
            .I(N__28942));
    Odrv12 I__4223 (
            .O(N__28942),
            .I(\current_shift_inst.PI_CTRL.integrator_1_15 ));
    InMux I__4222 (
            .O(N__28939),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ));
    CascadeMux I__4221 (
            .O(N__28936),
            .I(N__28933));
    InMux I__4220 (
            .O(N__28933),
            .I(N__28930));
    LocalMux I__4219 (
            .O(N__28930),
            .I(N__28927));
    Span4Mux_h I__4218 (
            .O(N__28927),
            .I(N__28924));
    Odrv4 I__4217 (
            .O(N__28924),
            .I(\current_shift_inst.PI_CTRL.integrator_1_16 ));
    InMux I__4216 (
            .O(N__28921),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ));
    InMux I__4215 (
            .O(N__28918),
            .I(N__28915));
    LocalMux I__4214 (
            .O(N__28915),
            .I(N__28912));
    Odrv4 I__4213 (
            .O(N__28912),
            .I(\current_shift_inst.PI_CTRL.integrator_1_17 ));
    InMux I__4212 (
            .O(N__28909),
            .I(bfn_9_20_0_));
    InMux I__4211 (
            .O(N__28906),
            .I(N__28903));
    LocalMux I__4210 (
            .O(N__28903),
            .I(\current_shift_inst.PI_CTRL.integrator_1_18 ));
    InMux I__4209 (
            .O(N__28900),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ));
    CascadeMux I__4208 (
            .O(N__28897),
            .I(N__28894));
    InMux I__4207 (
            .O(N__28894),
            .I(N__28891));
    LocalMux I__4206 (
            .O(N__28891),
            .I(\current_shift_inst.PI_CTRL.integrator_1_19 ));
    InMux I__4205 (
            .O(N__28888),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ));
    InMux I__4204 (
            .O(N__28885),
            .I(N__28882));
    LocalMux I__4203 (
            .O(N__28882),
            .I(\current_shift_inst.PI_CTRL.integrator_1_20 ));
    InMux I__4202 (
            .O(N__28879),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ));
    CascadeMux I__4201 (
            .O(N__28876),
            .I(N__28873));
    InMux I__4200 (
            .O(N__28873),
            .I(N__28870));
    LocalMux I__4199 (
            .O(N__28870),
            .I(N__28867));
    Span4Mux_v I__4198 (
            .O(N__28867),
            .I(N__28864));
    Sp12to4 I__4197 (
            .O(N__28864),
            .I(N__28861));
    Span12Mux_h I__4196 (
            .O(N__28861),
            .I(N__28858));
    Span12Mux_v I__4195 (
            .O(N__28858),
            .I(N__28855));
    Odrv12 I__4194 (
            .O(N__28855),
            .I(\current_shift_inst.PI_CTRL.integrator_1_5 ));
    InMux I__4193 (
            .O(N__28852),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ));
    CascadeMux I__4192 (
            .O(N__28849),
            .I(N__28846));
    InMux I__4191 (
            .O(N__28846),
            .I(N__28843));
    LocalMux I__4190 (
            .O(N__28843),
            .I(N__28840));
    Span4Mux_h I__4189 (
            .O(N__28840),
            .I(N__28837));
    Sp12to4 I__4188 (
            .O(N__28837),
            .I(N__28834));
    Span12Mux_v I__4187 (
            .O(N__28834),
            .I(N__28831));
    Odrv12 I__4186 (
            .O(N__28831),
            .I(\current_shift_inst.PI_CTRL.integrator_1_6 ));
    InMux I__4185 (
            .O(N__28828),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ));
    CascadeMux I__4184 (
            .O(N__28825),
            .I(N__28822));
    InMux I__4183 (
            .O(N__28822),
            .I(N__28819));
    LocalMux I__4182 (
            .O(N__28819),
            .I(N__28816));
    Span4Mux_v I__4181 (
            .O(N__28816),
            .I(N__28813));
    Sp12to4 I__4180 (
            .O(N__28813),
            .I(N__28810));
    Span12Mux_v I__4179 (
            .O(N__28810),
            .I(N__28807));
    Odrv12 I__4178 (
            .O(N__28807),
            .I(\current_shift_inst.PI_CTRL.integrator_1_7 ));
    InMux I__4177 (
            .O(N__28804),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ));
    CascadeMux I__4176 (
            .O(N__28801),
            .I(N__28798));
    InMux I__4175 (
            .O(N__28798),
            .I(N__28795));
    LocalMux I__4174 (
            .O(N__28795),
            .I(N__28792));
    Sp12to4 I__4173 (
            .O(N__28792),
            .I(N__28789));
    Span12Mux_v I__4172 (
            .O(N__28789),
            .I(N__28786));
    Odrv12 I__4171 (
            .O(N__28786),
            .I(\current_shift_inst.PI_CTRL.integrator_1_8 ));
    InMux I__4170 (
            .O(N__28783),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ));
    InMux I__4169 (
            .O(N__28780),
            .I(N__28777));
    LocalMux I__4168 (
            .O(N__28777),
            .I(N__28774));
    Span4Mux_v I__4167 (
            .O(N__28774),
            .I(N__28771));
    Sp12to4 I__4166 (
            .O(N__28771),
            .I(N__28768));
    Span12Mux_h I__4165 (
            .O(N__28768),
            .I(N__28765));
    Span12Mux_v I__4164 (
            .O(N__28765),
            .I(N__28762));
    Odrv12 I__4163 (
            .O(N__28762),
            .I(\current_shift_inst.PI_CTRL.integrator_1_9 ));
    InMux I__4162 (
            .O(N__28759),
            .I(bfn_9_19_0_));
    CascadeMux I__4161 (
            .O(N__28756),
            .I(N__28753));
    InMux I__4160 (
            .O(N__28753),
            .I(N__28750));
    LocalMux I__4159 (
            .O(N__28750),
            .I(N__28747));
    Span12Mux_h I__4158 (
            .O(N__28747),
            .I(N__28744));
    Span12Mux_v I__4157 (
            .O(N__28744),
            .I(N__28741));
    Odrv12 I__4156 (
            .O(N__28741),
            .I(\current_shift_inst.PI_CTRL.integrator_1_10 ));
    InMux I__4155 (
            .O(N__28738),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ));
    CascadeMux I__4154 (
            .O(N__28735),
            .I(N__28732));
    InMux I__4153 (
            .O(N__28732),
            .I(N__28729));
    LocalMux I__4152 (
            .O(N__28729),
            .I(N__28726));
    Span4Mux_v I__4151 (
            .O(N__28726),
            .I(N__28723));
    Sp12to4 I__4150 (
            .O(N__28723),
            .I(N__28720));
    Span12Mux_h I__4149 (
            .O(N__28720),
            .I(N__28717));
    Odrv12 I__4148 (
            .O(N__28717),
            .I(\current_shift_inst.PI_CTRL.integrator_1_11 ));
    InMux I__4147 (
            .O(N__28714),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ));
    CascadeMux I__4146 (
            .O(N__28711),
            .I(N__28708));
    InMux I__4145 (
            .O(N__28708),
            .I(N__28705));
    LocalMux I__4144 (
            .O(N__28705),
            .I(N__28702));
    Span4Mux_v I__4143 (
            .O(N__28702),
            .I(N__28699));
    Span4Mux_h I__4142 (
            .O(N__28699),
            .I(N__28696));
    Sp12to4 I__4141 (
            .O(N__28696),
            .I(N__28693));
    Span12Mux_v I__4140 (
            .O(N__28693),
            .I(N__28690));
    Odrv12 I__4139 (
            .O(N__28690),
            .I(\current_shift_inst.PI_CTRL.integrator_1_12 ));
    InMux I__4138 (
            .O(N__28687),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ));
    InMux I__4137 (
            .O(N__28684),
            .I(N__28681));
    LocalMux I__4136 (
            .O(N__28681),
            .I(N__28677));
    InMux I__4135 (
            .O(N__28680),
            .I(N__28674));
    Odrv12 I__4134 (
            .O(N__28677),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_25));
    LocalMux I__4133 (
            .O(N__28674),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_25));
    InMux I__4132 (
            .O(N__28669),
            .I(N__28663));
    InMux I__4131 (
            .O(N__28668),
            .I(N__28663));
    LocalMux I__4130 (
            .O(N__28663),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ));
    InMux I__4129 (
            .O(N__28660),
            .I(N__28657));
    LocalMux I__4128 (
            .O(N__28657),
            .I(N__28653));
    InMux I__4127 (
            .O(N__28656),
            .I(N__28650));
    Odrv4 I__4126 (
            .O(N__28653),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_26));
    LocalMux I__4125 (
            .O(N__28650),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_26));
    InMux I__4124 (
            .O(N__28645),
            .I(N__28639));
    InMux I__4123 (
            .O(N__28644),
            .I(N__28639));
    LocalMux I__4122 (
            .O(N__28639),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ));
    InMux I__4121 (
            .O(N__28636),
            .I(N__28633));
    LocalMux I__4120 (
            .O(N__28633),
            .I(N__28629));
    InMux I__4119 (
            .O(N__28632),
            .I(N__28626));
    Odrv4 I__4118 (
            .O(N__28629),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_27));
    LocalMux I__4117 (
            .O(N__28626),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_27));
    InMux I__4116 (
            .O(N__28621),
            .I(N__28615));
    InMux I__4115 (
            .O(N__28620),
            .I(N__28615));
    LocalMux I__4114 (
            .O(N__28615),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ));
    CascadeMux I__4113 (
            .O(N__28612),
            .I(N__28609));
    InMux I__4112 (
            .O(N__28609),
            .I(N__28606));
    LocalMux I__4111 (
            .O(N__28606),
            .I(N__28603));
    Span4Mux_v I__4110 (
            .O(N__28603),
            .I(N__28600));
    Sp12to4 I__4109 (
            .O(N__28600),
            .I(N__28597));
    Span12Mux_h I__4108 (
            .O(N__28597),
            .I(N__28594));
    Span12Mux_v I__4107 (
            .O(N__28594),
            .I(N__28591));
    Odrv12 I__4106 (
            .O(N__28591),
            .I(\current_shift_inst.PI_CTRL.un1_integrator ));
    CascadeMux I__4105 (
            .O(N__28588),
            .I(N__28585));
    InMux I__4104 (
            .O(N__28585),
            .I(N__28582));
    LocalMux I__4103 (
            .O(N__28582),
            .I(N__28579));
    Span4Mux_v I__4102 (
            .O(N__28579),
            .I(N__28576));
    Sp12to4 I__4101 (
            .O(N__28576),
            .I(N__28573));
    Span12Mux_h I__4100 (
            .O(N__28573),
            .I(N__28570));
    Odrv12 I__4099 (
            .O(N__28570),
            .I(\current_shift_inst.PI_CTRL.integrator_1_2 ));
    InMux I__4098 (
            .O(N__28567),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ));
    CascadeMux I__4097 (
            .O(N__28564),
            .I(N__28561));
    InMux I__4096 (
            .O(N__28561),
            .I(N__28558));
    LocalMux I__4095 (
            .O(N__28558),
            .I(N__28555));
    Span4Mux_v I__4094 (
            .O(N__28555),
            .I(N__28552));
    Sp12to4 I__4093 (
            .O(N__28552),
            .I(N__28549));
    Span12Mux_h I__4092 (
            .O(N__28549),
            .I(N__28546));
    Odrv12 I__4091 (
            .O(N__28546),
            .I(\current_shift_inst.PI_CTRL.integrator_1_3 ));
    InMux I__4090 (
            .O(N__28543),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ));
    CascadeMux I__4089 (
            .O(N__28540),
            .I(N__28537));
    InMux I__4088 (
            .O(N__28537),
            .I(N__28534));
    LocalMux I__4087 (
            .O(N__28534),
            .I(N__28531));
    Span4Mux_v I__4086 (
            .O(N__28531),
            .I(N__28528));
    Sp12to4 I__4085 (
            .O(N__28528),
            .I(N__28525));
    Span12Mux_h I__4084 (
            .O(N__28525),
            .I(N__28522));
    Odrv12 I__4083 (
            .O(N__28522),
            .I(\current_shift_inst.PI_CTRL.integrator_1_4 ));
    InMux I__4082 (
            .O(N__28519),
            .I(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ));
    InMux I__4081 (
            .O(N__28516),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6 ));
    InMux I__4080 (
            .O(N__28513),
            .I(N__28510));
    LocalMux I__4079 (
            .O(N__28510),
            .I(N__28507));
    Span12Mux_h I__4078 (
            .O(N__28507),
            .I(N__28504));
    Odrv12 I__4077 (
            .O(N__28504),
            .I(\pwm_generator_inst.un2_threshold_2_8 ));
    InMux I__4076 (
            .O(N__28501),
            .I(N__28498));
    LocalMux I__4075 (
            .O(N__28498),
            .I(N__28495));
    Span4Mux_v I__4074 (
            .O(N__28495),
            .I(N__28492));
    Sp12to4 I__4073 (
            .O(N__28492),
            .I(N__28489));
    Span12Mux_s9_h I__4072 (
            .O(N__28489),
            .I(N__28486));
    Odrv12 I__4071 (
            .O(N__28486),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ));
    InMux I__4070 (
            .O(N__28483),
            .I(bfn_9_16_0_));
    CascadeMux I__4069 (
            .O(N__28480),
            .I(N__28477));
    InMux I__4068 (
            .O(N__28477),
            .I(N__28474));
    LocalMux I__4067 (
            .O(N__28474),
            .I(N__28471));
    Span4Mux_h I__4066 (
            .O(N__28471),
            .I(N__28468));
    Span4Mux_h I__4065 (
            .O(N__28468),
            .I(N__28465));
    Odrv4 I__4064 (
            .O(N__28465),
            .I(\pwm_generator_inst.un2_threshold_2_9 ));
    InMux I__4063 (
            .O(N__28462),
            .I(N__28459));
    LocalMux I__4062 (
            .O(N__28459),
            .I(N__28456));
    Span12Mux_s9_h I__4061 (
            .O(N__28456),
            .I(N__28453));
    Odrv12 I__4060 (
            .O(N__28453),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ));
    InMux I__4059 (
            .O(N__28450),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_8 ));
    InMux I__4058 (
            .O(N__28447),
            .I(N__28444));
    LocalMux I__4057 (
            .O(N__28444),
            .I(N__28441));
    Span12Mux_h I__4056 (
            .O(N__28441),
            .I(N__28438));
    Odrv12 I__4055 (
            .O(N__28438),
            .I(\pwm_generator_inst.un2_threshold_2_10 ));
    InMux I__4054 (
            .O(N__28435),
            .I(N__28432));
    LocalMux I__4053 (
            .O(N__28432),
            .I(N__28429));
    Span4Mux_v I__4052 (
            .O(N__28429),
            .I(N__28426));
    Sp12to4 I__4051 (
            .O(N__28426),
            .I(N__28423));
    Span12Mux_s9_h I__4050 (
            .O(N__28423),
            .I(N__28420));
    Odrv12 I__4049 (
            .O(N__28420),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ));
    InMux I__4048 (
            .O(N__28417),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_9 ));
    CascadeMux I__4047 (
            .O(N__28414),
            .I(N__28406));
    CascadeMux I__4046 (
            .O(N__28413),
            .I(N__28402));
    CascadeMux I__4045 (
            .O(N__28412),
            .I(N__28398));
    CascadeMux I__4044 (
            .O(N__28411),
            .I(N__28395));
    CascadeMux I__4043 (
            .O(N__28410),
            .I(N__28392));
    CascadeMux I__4042 (
            .O(N__28409),
            .I(N__28389));
    InMux I__4041 (
            .O(N__28406),
            .I(N__28385));
    InMux I__4040 (
            .O(N__28405),
            .I(N__28376));
    InMux I__4039 (
            .O(N__28402),
            .I(N__28376));
    InMux I__4038 (
            .O(N__28401),
            .I(N__28376));
    InMux I__4037 (
            .O(N__28398),
            .I(N__28376));
    InMux I__4036 (
            .O(N__28395),
            .I(N__28373));
    InMux I__4035 (
            .O(N__28392),
            .I(N__28366));
    InMux I__4034 (
            .O(N__28389),
            .I(N__28366));
    InMux I__4033 (
            .O(N__28388),
            .I(N__28366));
    LocalMux I__4032 (
            .O(N__28385),
            .I(N__28363));
    LocalMux I__4031 (
            .O(N__28376),
            .I(N__28360));
    LocalMux I__4030 (
            .O(N__28373),
            .I(N__28355));
    LocalMux I__4029 (
            .O(N__28366),
            .I(N__28355));
    Span12Mux_s10_v I__4028 (
            .O(N__28363),
            .I(N__28352));
    Span4Mux_v I__4027 (
            .O(N__28360),
            .I(N__28347));
    Span4Mux_v I__4026 (
            .O(N__28355),
            .I(N__28347));
    Span12Mux_h I__4025 (
            .O(N__28352),
            .I(N__28344));
    Sp12to4 I__4024 (
            .O(N__28347),
            .I(N__28341));
    Span12Mux_h I__4023 (
            .O(N__28344),
            .I(N__28338));
    Span12Mux_h I__4022 (
            .O(N__28341),
            .I(N__28335));
    Odrv12 I__4021 (
            .O(N__28338),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    Odrv12 I__4020 (
            .O(N__28335),
            .I(\pwm_generator_inst.un2_threshold_1_19 ));
    CascadeMux I__4019 (
            .O(N__28330),
            .I(N__28327));
    InMux I__4018 (
            .O(N__28327),
            .I(N__28324));
    LocalMux I__4017 (
            .O(N__28324),
            .I(N__28321));
    Span4Mux_h I__4016 (
            .O(N__28321),
            .I(N__28318));
    Span4Mux_h I__4015 (
            .O(N__28318),
            .I(N__28315));
    Odrv4 I__4014 (
            .O(N__28315),
            .I(\pwm_generator_inst.un2_threshold_2_11 ));
    InMux I__4013 (
            .O(N__28312),
            .I(N__28309));
    LocalMux I__4012 (
            .O(N__28309),
            .I(N__28306));
    Sp12to4 I__4011 (
            .O(N__28306),
            .I(N__28303));
    Span12Mux_v I__4010 (
            .O(N__28303),
            .I(N__28300));
    Odrv12 I__4009 (
            .O(N__28300),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ));
    InMux I__4008 (
            .O(N__28297),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10 ));
    InMux I__4007 (
            .O(N__28294),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11 ));
    InMux I__4006 (
            .O(N__28291),
            .I(N__28288));
    LocalMux I__4005 (
            .O(N__28288),
            .I(N__28285));
    Span12Mux_v I__4004 (
            .O(N__28285),
            .I(N__28282));
    Odrv12 I__4003 (
            .O(N__28282),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO ));
    InMux I__4002 (
            .O(N__28279),
            .I(N__28276));
    LocalMux I__4001 (
            .O(N__28276),
            .I(N__28272));
    InMux I__4000 (
            .O(N__28275),
            .I(N__28269));
    Odrv12 I__3999 (
            .O(N__28272),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_24));
    LocalMux I__3998 (
            .O(N__28269),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_24));
    CascadeMux I__3997 (
            .O(N__28264),
            .I(N__28260));
    CascadeMux I__3996 (
            .O(N__28263),
            .I(N__28257));
    InMux I__3995 (
            .O(N__28260),
            .I(N__28252));
    InMux I__3994 (
            .O(N__28257),
            .I(N__28252));
    LocalMux I__3993 (
            .O(N__28252),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ));
    InMux I__3992 (
            .O(N__28249),
            .I(N__28246));
    LocalMux I__3991 (
            .O(N__28246),
            .I(N__28243));
    Span12Mux_h I__3990 (
            .O(N__28243),
            .I(N__28240));
    Odrv12 I__3989 (
            .O(N__28240),
            .I(\pwm_generator_inst.un2_threshold_2_0 ));
    CascadeMux I__3988 (
            .O(N__28237),
            .I(N__28234));
    InMux I__3987 (
            .O(N__28234),
            .I(N__28231));
    LocalMux I__3986 (
            .O(N__28231),
            .I(N__28228));
    Span4Mux_v I__3985 (
            .O(N__28228),
            .I(N__28225));
    Span4Mux_h I__3984 (
            .O(N__28225),
            .I(N__28222));
    Sp12to4 I__3983 (
            .O(N__28222),
            .I(N__28219));
    Odrv12 I__3982 (
            .O(N__28219),
            .I(\pwm_generator_inst.un2_threshold_1_15 ));
    InMux I__3981 (
            .O(N__28216),
            .I(N__28213));
    LocalMux I__3980 (
            .O(N__28213),
            .I(N__28210));
    Span4Mux_v I__3979 (
            .O(N__28210),
            .I(N__28207));
    Span4Mux_h I__3978 (
            .O(N__28207),
            .I(N__28204));
    Span4Mux_h I__3977 (
            .O(N__28204),
            .I(N__28201));
    Span4Mux_v I__3976 (
            .O(N__28201),
            .I(N__28198));
    Odrv4 I__3975 (
            .O(N__28198),
            .I(\pwm_generator_inst.un3_threshold_axbZ0Z_8 ));
    InMux I__3974 (
            .O(N__28195),
            .I(N__28192));
    LocalMux I__3973 (
            .O(N__28192),
            .I(N__28189));
    Span4Mux_h I__3972 (
            .O(N__28189),
            .I(N__28186));
    Span4Mux_h I__3971 (
            .O(N__28186),
            .I(N__28183));
    Odrv4 I__3970 (
            .O(N__28183),
            .I(\pwm_generator_inst.un2_threshold_2_1 ));
    CascadeMux I__3969 (
            .O(N__28180),
            .I(N__28177));
    InMux I__3968 (
            .O(N__28177),
            .I(N__28174));
    LocalMux I__3967 (
            .O(N__28174),
            .I(N__28171));
    Span4Mux_h I__3966 (
            .O(N__28171),
            .I(N__28168));
    Span4Mux_h I__3965 (
            .O(N__28168),
            .I(N__28165));
    Span4Mux_h I__3964 (
            .O(N__28165),
            .I(N__28162));
    Span4Mux_h I__3963 (
            .O(N__28162),
            .I(N__28159));
    Odrv4 I__3962 (
            .O(N__28159),
            .I(\pwm_generator_inst.un2_threshold_1_16 ));
    InMux I__3961 (
            .O(N__28156),
            .I(N__28153));
    LocalMux I__3960 (
            .O(N__28153),
            .I(N__28150));
    Span12Mux_s9_h I__3959 (
            .O(N__28150),
            .I(N__28147));
    Odrv12 I__3958 (
            .O(N__28147),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ));
    InMux I__3957 (
            .O(N__28144),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_0 ));
    InMux I__3956 (
            .O(N__28141),
            .I(N__28138));
    LocalMux I__3955 (
            .O(N__28138),
            .I(N__28135));
    Span4Mux_v I__3954 (
            .O(N__28135),
            .I(N__28132));
    Sp12to4 I__3953 (
            .O(N__28132),
            .I(N__28129));
    Span12Mux_h I__3952 (
            .O(N__28129),
            .I(N__28126));
    Odrv12 I__3951 (
            .O(N__28126),
            .I(\pwm_generator_inst.un2_threshold_1_17 ));
    CascadeMux I__3950 (
            .O(N__28123),
            .I(N__28120));
    InMux I__3949 (
            .O(N__28120),
            .I(N__28117));
    LocalMux I__3948 (
            .O(N__28117),
            .I(N__28114));
    Span12Mux_h I__3947 (
            .O(N__28114),
            .I(N__28111));
    Odrv12 I__3946 (
            .O(N__28111),
            .I(\pwm_generator_inst.un2_threshold_2_2 ));
    InMux I__3945 (
            .O(N__28108),
            .I(N__28105));
    LocalMux I__3944 (
            .O(N__28105),
            .I(N__28102));
    Span4Mux_v I__3943 (
            .O(N__28102),
            .I(N__28099));
    Span4Mux_h I__3942 (
            .O(N__28099),
            .I(N__28096));
    Span4Mux_h I__3941 (
            .O(N__28096),
            .I(N__28093));
    Span4Mux_v I__3940 (
            .O(N__28093),
            .I(N__28090));
    Odrv4 I__3939 (
            .O(N__28090),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ));
    InMux I__3938 (
            .O(N__28087),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_1 ));
    InMux I__3937 (
            .O(N__28084),
            .I(N__28081));
    LocalMux I__3936 (
            .O(N__28081),
            .I(N__28078));
    Span4Mux_v I__3935 (
            .O(N__28078),
            .I(N__28075));
    Sp12to4 I__3934 (
            .O(N__28075),
            .I(N__28072));
    Span12Mux_h I__3933 (
            .O(N__28072),
            .I(N__28069));
    Odrv12 I__3932 (
            .O(N__28069),
            .I(\pwm_generator_inst.un2_threshold_1_18 ));
    CascadeMux I__3931 (
            .O(N__28066),
            .I(N__28063));
    InMux I__3930 (
            .O(N__28063),
            .I(N__28060));
    LocalMux I__3929 (
            .O(N__28060),
            .I(N__28057));
    Span12Mux_h I__3928 (
            .O(N__28057),
            .I(N__28054));
    Odrv12 I__3927 (
            .O(N__28054),
            .I(\pwm_generator_inst.un2_threshold_2_3 ));
    InMux I__3926 (
            .O(N__28051),
            .I(N__28048));
    LocalMux I__3925 (
            .O(N__28048),
            .I(N__28045));
    Sp12to4 I__3924 (
            .O(N__28045),
            .I(N__28042));
    Span12Mux_v I__3923 (
            .O(N__28042),
            .I(N__28039));
    Odrv12 I__3922 (
            .O(N__28039),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ));
    InMux I__3921 (
            .O(N__28036),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_2 ));
    CascadeMux I__3920 (
            .O(N__28033),
            .I(N__28030));
    InMux I__3919 (
            .O(N__28030),
            .I(N__28027));
    LocalMux I__3918 (
            .O(N__28027),
            .I(N__28024));
    Span4Mux_h I__3917 (
            .O(N__28024),
            .I(N__28021));
    Span4Mux_h I__3916 (
            .O(N__28021),
            .I(N__28018));
    Odrv4 I__3915 (
            .O(N__28018),
            .I(\pwm_generator_inst.un2_threshold_2_4 ));
    InMux I__3914 (
            .O(N__28015),
            .I(N__28012));
    LocalMux I__3913 (
            .O(N__28012),
            .I(N__28009));
    Span12Mux_v I__3912 (
            .O(N__28009),
            .I(N__28006));
    Odrv12 I__3911 (
            .O(N__28006),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ));
    InMux I__3910 (
            .O(N__28003),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_3 ));
    InMux I__3909 (
            .O(N__28000),
            .I(N__27997));
    LocalMux I__3908 (
            .O(N__27997),
            .I(N__27994));
    Odrv12 I__3907 (
            .O(N__27994),
            .I(\pwm_generator_inst.un2_threshold_2_5 ));
    InMux I__3906 (
            .O(N__27991),
            .I(N__27988));
    LocalMux I__3905 (
            .O(N__27988),
            .I(N__27985));
    Span4Mux_v I__3904 (
            .O(N__27985),
            .I(N__27982));
    Sp12to4 I__3903 (
            .O(N__27982),
            .I(N__27979));
    Span12Mux_s9_h I__3902 (
            .O(N__27979),
            .I(N__27976));
    Odrv12 I__3901 (
            .O(N__27976),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ));
    InMux I__3900 (
            .O(N__27973),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_4 ));
    InMux I__3899 (
            .O(N__27970),
            .I(N__27967));
    LocalMux I__3898 (
            .O(N__27967),
            .I(N__27964));
    Odrv12 I__3897 (
            .O(N__27964),
            .I(\pwm_generator_inst.un2_threshold_2_6 ));
    InMux I__3896 (
            .O(N__27961),
            .I(N__27958));
    LocalMux I__3895 (
            .O(N__27958),
            .I(N__27955));
    Span4Mux_v I__3894 (
            .O(N__27955),
            .I(N__27952));
    Sp12to4 I__3893 (
            .O(N__27952),
            .I(N__27949));
    Span12Mux_s9_h I__3892 (
            .O(N__27949),
            .I(N__27946));
    Odrv12 I__3891 (
            .O(N__27946),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ));
    InMux I__3890 (
            .O(N__27943),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_5 ));
    InMux I__3889 (
            .O(N__27940),
            .I(N__27937));
    LocalMux I__3888 (
            .O(N__27937),
            .I(N__27934));
    Sp12to4 I__3887 (
            .O(N__27934),
            .I(N__27931));
    Odrv12 I__3886 (
            .O(N__27931),
            .I(\pwm_generator_inst.un2_threshold_2_7 ));
    InMux I__3885 (
            .O(N__27928),
            .I(N__27925));
    LocalMux I__3884 (
            .O(N__27925),
            .I(N__27922));
    Span4Mux_v I__3883 (
            .O(N__27922),
            .I(N__27919));
    Sp12to4 I__3882 (
            .O(N__27919),
            .I(N__27916));
    Span12Mux_s9_h I__3881 (
            .O(N__27916),
            .I(N__27913));
    Odrv12 I__3880 (
            .O(N__27913),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ));
    InMux I__3879 (
            .O(N__27910),
            .I(N__27906));
    InMux I__3878 (
            .O(N__27909),
            .I(N__27903));
    LocalMux I__3877 (
            .O(N__27906),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ));
    LocalMux I__3876 (
            .O(N__27903),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ));
    InMux I__3875 (
            .O(N__27898),
            .I(bfn_9_14_0_));
    InMux I__3874 (
            .O(N__27895),
            .I(N__27892));
    LocalMux I__3873 (
            .O(N__27892),
            .I(N__27889));
    Odrv4 I__3872 (
            .O(N__27889),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ));
    InMux I__3871 (
            .O(N__27886),
            .I(N__27882));
    InMux I__3870 (
            .O(N__27885),
            .I(N__27879));
    LocalMux I__3869 (
            .O(N__27882),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ));
    LocalMux I__3868 (
            .O(N__27879),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ));
    InMux I__3867 (
            .O(N__27874),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ));
    InMux I__3866 (
            .O(N__27871),
            .I(N__27868));
    LocalMux I__3865 (
            .O(N__27868),
            .I(N__27865));
    Span4Mux_v I__3864 (
            .O(N__27865),
            .I(N__27862));
    Odrv4 I__3863 (
            .O(N__27862),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ));
    InMux I__3862 (
            .O(N__27859),
            .I(N__27855));
    InMux I__3861 (
            .O(N__27858),
            .I(N__27852));
    LocalMux I__3860 (
            .O(N__27855),
            .I(N__27847));
    LocalMux I__3859 (
            .O(N__27852),
            .I(N__27847));
    Span4Mux_v I__3858 (
            .O(N__27847),
            .I(N__27844));
    Odrv4 I__3857 (
            .O(N__27844),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ));
    InMux I__3856 (
            .O(N__27841),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ));
    InMux I__3855 (
            .O(N__27838),
            .I(N__27835));
    LocalMux I__3854 (
            .O(N__27835),
            .I(N__27831));
    InMux I__3853 (
            .O(N__27834),
            .I(N__27828));
    Span4Mux_v I__3852 (
            .O(N__27831),
            .I(N__27825));
    LocalMux I__3851 (
            .O(N__27828),
            .I(N__27822));
    Odrv4 I__3850 (
            .O(N__27825),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ));
    Odrv4 I__3849 (
            .O(N__27822),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ));
    InMux I__3848 (
            .O(N__27817),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ));
    InMux I__3847 (
            .O(N__27814),
            .I(N__27811));
    LocalMux I__3846 (
            .O(N__27811),
            .I(N__27808));
    Span4Mux_h I__3845 (
            .O(N__27808),
            .I(N__27805));
    Odrv4 I__3844 (
            .O(N__27805),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ));
    InMux I__3843 (
            .O(N__27802),
            .I(N__27799));
    LocalMux I__3842 (
            .O(N__27799),
            .I(N__27795));
    InMux I__3841 (
            .O(N__27798),
            .I(N__27792));
    Span4Mux_h I__3840 (
            .O(N__27795),
            .I(N__27789));
    LocalMux I__3839 (
            .O(N__27792),
            .I(N__27786));
    Odrv4 I__3838 (
            .O(N__27789),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ));
    Odrv4 I__3837 (
            .O(N__27786),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ));
    InMux I__3836 (
            .O(N__27781),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ));
    InMux I__3835 (
            .O(N__27778),
            .I(N__27774));
    InMux I__3834 (
            .O(N__27777),
            .I(N__27771));
    LocalMux I__3833 (
            .O(N__27774),
            .I(N__27768));
    LocalMux I__3832 (
            .O(N__27771),
            .I(N__27763));
    Span4Mux_h I__3831 (
            .O(N__27768),
            .I(N__27763));
    Odrv4 I__3830 (
            .O(N__27763),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ));
    InMux I__3829 (
            .O(N__27760),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ));
    InMux I__3828 (
            .O(N__27757),
            .I(N__27754));
    LocalMux I__3827 (
            .O(N__27754),
            .I(N__27751));
    Odrv4 I__3826 (
            .O(N__27751),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ));
    InMux I__3825 (
            .O(N__27748),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ));
    InMux I__3824 (
            .O(N__27745),
            .I(N__27741));
    InMux I__3823 (
            .O(N__27744),
            .I(N__27738));
    LocalMux I__3822 (
            .O(N__27741),
            .I(N__27735));
    LocalMux I__3821 (
            .O(N__27738),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    Odrv12 I__3820 (
            .O(N__27735),
            .I(elapsed_time_ns_1_RNI6HPBB_0_28));
    InMux I__3819 (
            .O(N__27730),
            .I(N__27727));
    LocalMux I__3818 (
            .O(N__27727),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ));
    InMux I__3817 (
            .O(N__27724),
            .I(N__27720));
    InMux I__3816 (
            .O(N__27723),
            .I(N__27717));
    LocalMux I__3815 (
            .O(N__27720),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ));
    LocalMux I__3814 (
            .O(N__27717),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ));
    InMux I__3813 (
            .O(N__27712),
            .I(bfn_9_13_0_));
    InMux I__3812 (
            .O(N__27709),
            .I(N__27706));
    LocalMux I__3811 (
            .O(N__27706),
            .I(N__27703));
    Odrv12 I__3810 (
            .O(N__27703),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ));
    InMux I__3809 (
            .O(N__27700),
            .I(N__27696));
    InMux I__3808 (
            .O(N__27699),
            .I(N__27693));
    LocalMux I__3807 (
            .O(N__27696),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ));
    LocalMux I__3806 (
            .O(N__27693),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ));
    InMux I__3805 (
            .O(N__27688),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ));
    InMux I__3804 (
            .O(N__27685),
            .I(N__27682));
    LocalMux I__3803 (
            .O(N__27682),
            .I(N__27679));
    Odrv4 I__3802 (
            .O(N__27679),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ));
    InMux I__3801 (
            .O(N__27676),
            .I(N__27672));
    InMux I__3800 (
            .O(N__27675),
            .I(N__27669));
    LocalMux I__3799 (
            .O(N__27672),
            .I(N__27664));
    LocalMux I__3798 (
            .O(N__27669),
            .I(N__27664));
    Span4Mux_v I__3797 (
            .O(N__27664),
            .I(N__27661));
    Odrv4 I__3796 (
            .O(N__27661),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ));
    InMux I__3795 (
            .O(N__27658),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ));
    InMux I__3794 (
            .O(N__27655),
            .I(N__27652));
    LocalMux I__3793 (
            .O(N__27652),
            .I(N__27648));
    InMux I__3792 (
            .O(N__27651),
            .I(N__27645));
    Span4Mux_v I__3791 (
            .O(N__27648),
            .I(N__27642));
    LocalMux I__3790 (
            .O(N__27645),
            .I(N__27639));
    Odrv4 I__3789 (
            .O(N__27642),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ));
    Odrv4 I__3788 (
            .O(N__27639),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ));
    InMux I__3787 (
            .O(N__27634),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ));
    InMux I__3786 (
            .O(N__27631),
            .I(N__27628));
    LocalMux I__3785 (
            .O(N__27628),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ));
    InMux I__3784 (
            .O(N__27625),
            .I(N__27622));
    LocalMux I__3783 (
            .O(N__27622),
            .I(N__27618));
    InMux I__3782 (
            .O(N__27621),
            .I(N__27615));
    Span4Mux_v I__3781 (
            .O(N__27618),
            .I(N__27612));
    LocalMux I__3780 (
            .O(N__27615),
            .I(N__27609));
    Odrv4 I__3779 (
            .O(N__27612),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ));
    Odrv4 I__3778 (
            .O(N__27609),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ));
    InMux I__3777 (
            .O(N__27604),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ));
    InMux I__3776 (
            .O(N__27601),
            .I(N__27597));
    InMux I__3775 (
            .O(N__27600),
            .I(N__27594));
    LocalMux I__3774 (
            .O(N__27597),
            .I(N__27591));
    LocalMux I__3773 (
            .O(N__27594),
            .I(N__27588));
    Span4Mux_v I__3772 (
            .O(N__27591),
            .I(N__27585));
    Odrv4 I__3771 (
            .O(N__27588),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ));
    Odrv4 I__3770 (
            .O(N__27585),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ));
    InMux I__3769 (
            .O(N__27580),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ));
    InMux I__3768 (
            .O(N__27577),
            .I(N__27574));
    LocalMux I__3767 (
            .O(N__27574),
            .I(N__27571));
    Span4Mux_v I__3766 (
            .O(N__27571),
            .I(N__27568));
    Odrv4 I__3765 (
            .O(N__27568),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ));
    InMux I__3764 (
            .O(N__27565),
            .I(N__27562));
    LocalMux I__3763 (
            .O(N__27562),
            .I(N__27558));
    InMux I__3762 (
            .O(N__27561),
            .I(N__27555));
    Span4Mux_h I__3761 (
            .O(N__27558),
            .I(N__27550));
    LocalMux I__3760 (
            .O(N__27555),
            .I(N__27550));
    Odrv4 I__3759 (
            .O(N__27550),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ));
    InMux I__3758 (
            .O(N__27547),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ));
    InMux I__3757 (
            .O(N__27544),
            .I(N__27540));
    InMux I__3756 (
            .O(N__27543),
            .I(N__27537));
    LocalMux I__3755 (
            .O(N__27540),
            .I(N__27534));
    LocalMux I__3754 (
            .O(N__27537),
            .I(N__27529));
    Span4Mux_h I__3753 (
            .O(N__27534),
            .I(N__27529));
    Odrv4 I__3752 (
            .O(N__27529),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ));
    InMux I__3751 (
            .O(N__27526),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ));
    InMux I__3750 (
            .O(N__27523),
            .I(N__27520));
    LocalMux I__3749 (
            .O(N__27520),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ));
    InMux I__3748 (
            .O(N__27517),
            .I(N__27514));
    LocalMux I__3747 (
            .O(N__27514),
            .I(N__27510));
    InMux I__3746 (
            .O(N__27513),
            .I(N__27507));
    Span4Mux_h I__3745 (
            .O(N__27510),
            .I(N__27504));
    LocalMux I__3744 (
            .O(N__27507),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ));
    Odrv4 I__3743 (
            .O(N__27504),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ));
    InMux I__3742 (
            .O(N__27499),
            .I(bfn_9_12_0_));
    InMux I__3741 (
            .O(N__27496),
            .I(N__27493));
    LocalMux I__3740 (
            .O(N__27493),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ));
    InMux I__3739 (
            .O(N__27490),
            .I(N__27486));
    InMux I__3738 (
            .O(N__27489),
            .I(N__27483));
    LocalMux I__3737 (
            .O(N__27486),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ));
    LocalMux I__3736 (
            .O(N__27483),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ));
    InMux I__3735 (
            .O(N__27478),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ));
    InMux I__3734 (
            .O(N__27475),
            .I(N__27471));
    InMux I__3733 (
            .O(N__27474),
            .I(N__27468));
    LocalMux I__3732 (
            .O(N__27471),
            .I(N__27463));
    LocalMux I__3731 (
            .O(N__27468),
            .I(N__27463));
    Span4Mux_v I__3730 (
            .O(N__27463),
            .I(N__27460));
    Odrv4 I__3729 (
            .O(N__27460),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ));
    InMux I__3728 (
            .O(N__27457),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ));
    InMux I__3727 (
            .O(N__27454),
            .I(N__27451));
    LocalMux I__3726 (
            .O(N__27451),
            .I(N__27448));
    Odrv4 I__3725 (
            .O(N__27448),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ));
    InMux I__3724 (
            .O(N__27445),
            .I(N__27442));
    LocalMux I__3723 (
            .O(N__27442),
            .I(N__27438));
    InMux I__3722 (
            .O(N__27441),
            .I(N__27435));
    Span4Mux_v I__3721 (
            .O(N__27438),
            .I(N__27432));
    LocalMux I__3720 (
            .O(N__27435),
            .I(N__27429));
    Odrv4 I__3719 (
            .O(N__27432),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ));
    Odrv4 I__3718 (
            .O(N__27429),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ));
    InMux I__3717 (
            .O(N__27424),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ));
    InMux I__3716 (
            .O(N__27421),
            .I(N__27418));
    LocalMux I__3715 (
            .O(N__27418),
            .I(N__27414));
    InMux I__3714 (
            .O(N__27417),
            .I(N__27411));
    Span4Mux_h I__3713 (
            .O(N__27414),
            .I(N__27408));
    LocalMux I__3712 (
            .O(N__27411),
            .I(N__27405));
    Odrv4 I__3711 (
            .O(N__27408),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ));
    Odrv4 I__3710 (
            .O(N__27405),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ));
    InMux I__3709 (
            .O(N__27400),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ));
    InMux I__3708 (
            .O(N__27397),
            .I(N__27394));
    LocalMux I__3707 (
            .O(N__27394),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ));
    InMux I__3706 (
            .O(N__27391),
            .I(N__27387));
    InMux I__3705 (
            .O(N__27390),
            .I(N__27384));
    LocalMux I__3704 (
            .O(N__27387),
            .I(N__27381));
    LocalMux I__3703 (
            .O(N__27384),
            .I(N__27376));
    Span4Mux_h I__3702 (
            .O(N__27381),
            .I(N__27376));
    Odrv4 I__3701 (
            .O(N__27376),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ));
    InMux I__3700 (
            .O(N__27373),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ));
    InMux I__3699 (
            .O(N__27370),
            .I(N__27367));
    LocalMux I__3698 (
            .O(N__27367),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ));
    InMux I__3697 (
            .O(N__27364),
            .I(N__27361));
    LocalMux I__3696 (
            .O(N__27361),
            .I(N__27357));
    InMux I__3695 (
            .O(N__27360),
            .I(N__27354));
    Span4Mux_h I__3694 (
            .O(N__27357),
            .I(N__27351));
    LocalMux I__3693 (
            .O(N__27354),
            .I(N__27348));
    Odrv4 I__3692 (
            .O(N__27351),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ));
    Odrv4 I__3691 (
            .O(N__27348),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ));
    InMux I__3690 (
            .O(N__27343),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ));
    InMux I__3689 (
            .O(N__27340),
            .I(N__27337));
    LocalMux I__3688 (
            .O(N__27337),
            .I(N__27334));
    Odrv4 I__3687 (
            .O(N__27334),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ));
    InMux I__3686 (
            .O(N__27331),
            .I(N__27327));
    InMux I__3685 (
            .O(N__27330),
            .I(N__27324));
    LocalMux I__3684 (
            .O(N__27327),
            .I(N__27321));
    LocalMux I__3683 (
            .O(N__27324),
            .I(N__27316));
    Span4Mux_h I__3682 (
            .O(N__27321),
            .I(N__27316));
    Odrv4 I__3681 (
            .O(N__27316),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ));
    InMux I__3680 (
            .O(N__27313),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ));
    InMux I__3679 (
            .O(N__27310),
            .I(N__27307));
    LocalMux I__3678 (
            .O(N__27307),
            .I(N__27304));
    Span4Mux_v I__3677 (
            .O(N__27304),
            .I(N__27300));
    InMux I__3676 (
            .O(N__27303),
            .I(N__27297));
    Odrv4 I__3675 (
            .O(N__27300),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    LocalMux I__3674 (
            .O(N__27297),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ));
    InMux I__3673 (
            .O(N__27292),
            .I(N__27289));
    LocalMux I__3672 (
            .O(N__27289),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ));
    CascadeMux I__3671 (
            .O(N__27286),
            .I(N__27283));
    InMux I__3670 (
            .O(N__27283),
            .I(N__27280));
    LocalMux I__3669 (
            .O(N__27280),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ));
    InMux I__3668 (
            .O(N__27277),
            .I(N__27274));
    LocalMux I__3667 (
            .O(N__27274),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ));
    InMux I__3666 (
            .O(N__27271),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ));
    InMux I__3665 (
            .O(N__27268),
            .I(N__27265));
    LocalMux I__3664 (
            .O(N__27265),
            .I(N__27261));
    InMux I__3663 (
            .O(N__27264),
            .I(N__27258));
    Span4Mux_v I__3662 (
            .O(N__27261),
            .I(N__27255));
    LocalMux I__3661 (
            .O(N__27258),
            .I(N__27252));
    Odrv4 I__3660 (
            .O(N__27255),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ));
    Odrv4 I__3659 (
            .O(N__27252),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ));
    InMux I__3658 (
            .O(N__27247),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ));
    InMux I__3657 (
            .O(N__27244),
            .I(N__27241));
    LocalMux I__3656 (
            .O(N__27241),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ));
    InMux I__3655 (
            .O(N__27238),
            .I(N__27235));
    LocalMux I__3654 (
            .O(N__27235),
            .I(N__27232));
    Span4Mux_v I__3653 (
            .O(N__27232),
            .I(N__27228));
    InMux I__3652 (
            .O(N__27231),
            .I(N__27225));
    Span4Mux_v I__3651 (
            .O(N__27228),
            .I(N__27220));
    LocalMux I__3650 (
            .O(N__27225),
            .I(N__27220));
    Odrv4 I__3649 (
            .O(N__27220),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ));
    InMux I__3648 (
            .O(N__27217),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ));
    InMux I__3647 (
            .O(N__27214),
            .I(N__27210));
    InMux I__3646 (
            .O(N__27213),
            .I(N__27207));
    LocalMux I__3645 (
            .O(N__27210),
            .I(N__27204));
    LocalMux I__3644 (
            .O(N__27207),
            .I(N__27201));
    Span4Mux_h I__3643 (
            .O(N__27204),
            .I(N__27198));
    Odrv4 I__3642 (
            .O(N__27201),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ));
    Odrv4 I__3641 (
            .O(N__27198),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ));
    InMux I__3640 (
            .O(N__27193),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ));
    InMux I__3639 (
            .O(N__27190),
            .I(N__27187));
    LocalMux I__3638 (
            .O(N__27187),
            .I(N__27184));
    Odrv4 I__3637 (
            .O(N__27184),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ));
    InMux I__3636 (
            .O(N__27181),
            .I(N__27178));
    LocalMux I__3635 (
            .O(N__27178),
            .I(N__27174));
    InMux I__3634 (
            .O(N__27177),
            .I(N__27171));
    Span4Mux_h I__3633 (
            .O(N__27174),
            .I(N__27168));
    LocalMux I__3632 (
            .O(N__27171),
            .I(N__27165));
    Odrv4 I__3631 (
            .O(N__27168),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ));
    Odrv4 I__3630 (
            .O(N__27165),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ));
    InMux I__3629 (
            .O(N__27160),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ));
    InMux I__3628 (
            .O(N__27157),
            .I(N__27153));
    InMux I__3627 (
            .O(N__27156),
            .I(N__27150));
    LocalMux I__3626 (
            .O(N__27153),
            .I(N__27145));
    LocalMux I__3625 (
            .O(N__27150),
            .I(N__27145));
    Span4Mux_h I__3624 (
            .O(N__27145),
            .I(N__27142));
    Odrv4 I__3623 (
            .O(N__27142),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ));
    InMux I__3622 (
            .O(N__27139),
            .I(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ));
    InMux I__3621 (
            .O(N__27136),
            .I(N__27130));
    InMux I__3620 (
            .O(N__27135),
            .I(N__27130));
    LocalMux I__3619 (
            .O(N__27130),
            .I(elapsed_time_ns_1_RNIV8OBB_0_12));
    InMux I__3618 (
            .O(N__27127),
            .I(N__27123));
    InMux I__3617 (
            .O(N__27126),
            .I(N__27120));
    LocalMux I__3616 (
            .O(N__27123),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    LocalMux I__3615 (
            .O(N__27120),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ));
    InMux I__3614 (
            .O(N__27115),
            .I(N__27112));
    LocalMux I__3613 (
            .O(N__27112),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16));
    CascadeMux I__3612 (
            .O(N__27109),
            .I(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_));
    InMux I__3611 (
            .O(N__27106),
            .I(N__27102));
    InMux I__3610 (
            .O(N__27105),
            .I(N__27099));
    LocalMux I__3609 (
            .O(N__27102),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    LocalMux I__3608 (
            .O(N__27099),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ));
    InMux I__3607 (
            .O(N__27094),
            .I(N__27091));
    LocalMux I__3606 (
            .O(N__27091),
            .I(N__27087));
    InMux I__3605 (
            .O(N__27090),
            .I(N__27084));
    Odrv4 I__3604 (
            .O(N__27087),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    LocalMux I__3603 (
            .O(N__27084),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ));
    InMux I__3602 (
            .O(N__27079),
            .I(N__27076));
    LocalMux I__3601 (
            .O(N__27076),
            .I(N__27072));
    InMux I__3600 (
            .O(N__27075),
            .I(N__27069));
    Odrv4 I__3599 (
            .O(N__27072),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    LocalMux I__3598 (
            .O(N__27069),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ));
    InMux I__3597 (
            .O(N__27064),
            .I(N__27061));
    LocalMux I__3596 (
            .O(N__27061),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ));
    InMux I__3595 (
            .O(N__27058),
            .I(N__27055));
    LocalMux I__3594 (
            .O(N__27055),
            .I(N__27051));
    InMux I__3593 (
            .O(N__27054),
            .I(N__27048));
    Odrv4 I__3592 (
            .O(N__27051),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    LocalMux I__3591 (
            .O(N__27048),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ));
    InMux I__3590 (
            .O(N__27043),
            .I(N__27040));
    LocalMux I__3589 (
            .O(N__27040),
            .I(N__27037));
    Odrv4 I__3588 (
            .O(N__27037),
            .I(elapsed_time_ns_1_RNIHG91B_0_5));
    CascadeMux I__3587 (
            .O(N__27034),
            .I(elapsed_time_ns_1_RNIHG91B_0_5_cascade_));
    InMux I__3586 (
            .O(N__27031),
            .I(N__27027));
    InMux I__3585 (
            .O(N__27030),
            .I(N__27024));
    LocalMux I__3584 (
            .O(N__27027),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    LocalMux I__3583 (
            .O(N__27024),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ));
    CascadeMux I__3582 (
            .O(N__27019),
            .I(N__27015));
    InMux I__3581 (
            .O(N__27018),
            .I(N__27012));
    InMux I__3580 (
            .O(N__27015),
            .I(N__27009));
    LocalMux I__3579 (
            .O(N__27012),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    LocalMux I__3578 (
            .O(N__27009),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ));
    InMux I__3577 (
            .O(N__27004),
            .I(N__27001));
    LocalMux I__3576 (
            .O(N__27001),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ));
    InMux I__3575 (
            .O(N__26998),
            .I(N__26994));
    CascadeMux I__3574 (
            .O(N__26997),
            .I(N__26991));
    LocalMux I__3573 (
            .O(N__26994),
            .I(N__26988));
    InMux I__3572 (
            .O(N__26991),
            .I(N__26985));
    Odrv4 I__3571 (
            .O(N__26988),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    LocalMux I__3570 (
            .O(N__26985),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ));
    CascadeMux I__3569 (
            .O(N__26980),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ));
    InMux I__3568 (
            .O(N__26977),
            .I(N__26971));
    InMux I__3567 (
            .O(N__26976),
            .I(N__26971));
    LocalMux I__3566 (
            .O(N__26971),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ));
    InMux I__3565 (
            .O(N__26968),
            .I(N__26964));
    InMux I__3564 (
            .O(N__26967),
            .I(N__26961));
    LocalMux I__3563 (
            .O(N__26964),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    LocalMux I__3562 (
            .O(N__26961),
            .I(elapsed_time_ns_1_RNI5FOBB_0_18));
    InMux I__3561 (
            .O(N__26956),
            .I(N__26953));
    LocalMux I__3560 (
            .O(N__26953),
            .I(N__26949));
    InMux I__3559 (
            .O(N__26952),
            .I(N__26946));
    Odrv4 I__3558 (
            .O(N__26949),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    LocalMux I__3557 (
            .O(N__26946),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ));
    InMux I__3556 (
            .O(N__26941),
            .I(N__26937));
    CascadeMux I__3555 (
            .O(N__26940),
            .I(N__26934));
    LocalMux I__3554 (
            .O(N__26937),
            .I(N__26931));
    InMux I__3553 (
            .O(N__26934),
            .I(N__26928));
    Odrv12 I__3552 (
            .O(N__26931),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    LocalMux I__3551 (
            .O(N__26928),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ));
    InMux I__3550 (
            .O(N__26923),
            .I(N__26917));
    InMux I__3549 (
            .O(N__26922),
            .I(N__26917));
    LocalMux I__3548 (
            .O(N__26917),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ));
    InMux I__3547 (
            .O(N__26914),
            .I(N__26911));
    LocalMux I__3546 (
            .O(N__26911),
            .I(N__26907));
    InMux I__3545 (
            .O(N__26910),
            .I(N__26904));
    Odrv4 I__3544 (
            .O(N__26907),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    LocalMux I__3543 (
            .O(N__26904),
            .I(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ));
    CascadeMux I__3542 (
            .O(N__26899),
            .I(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ));
    InMux I__3541 (
            .O(N__26896),
            .I(N__26886));
    InMux I__3540 (
            .O(N__26895),
            .I(N__26886));
    InMux I__3539 (
            .O(N__26894),
            .I(N__26886));
    InMux I__3538 (
            .O(N__26893),
            .I(N__26883));
    LocalMux I__3537 (
            .O(N__26886),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    LocalMux I__3536 (
            .O(N__26883),
            .I(\phase_controller_inst2.stateZ0Z_2 ));
    CascadeMux I__3535 (
            .O(N__26878),
            .I(N__26874));
    CascadeMux I__3534 (
            .O(N__26877),
            .I(N__26871));
    InMux I__3533 (
            .O(N__26874),
            .I(N__26862));
    InMux I__3532 (
            .O(N__26871),
            .I(N__26862));
    InMux I__3531 (
            .O(N__26870),
            .I(N__26862));
    InMux I__3530 (
            .O(N__26869),
            .I(N__26859));
    LocalMux I__3529 (
            .O(N__26862),
            .I(\phase_controller_inst2.hc_time_passed ));
    LocalMux I__3528 (
            .O(N__26859),
            .I(\phase_controller_inst2.hc_time_passed ));
    InMux I__3527 (
            .O(N__26854),
            .I(N__26851));
    LocalMux I__3526 (
            .O(N__26851),
            .I(\phase_controller_inst2.start_timer_tr_0_sqmuxa ));
    InMux I__3525 (
            .O(N__26848),
            .I(N__26845));
    LocalMux I__3524 (
            .O(N__26845),
            .I(N__26842));
    Span4Mux_v I__3523 (
            .O(N__26842),
            .I(N__26839));
    Sp12to4 I__3522 (
            .O(N__26839),
            .I(N__26836));
    Span12Mux_h I__3521 (
            .O(N__26836),
            .I(N__26833));
    Odrv12 I__3520 (
            .O(N__26833),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_8 ));
    InMux I__3519 (
            .O(N__26830),
            .I(bfn_8_22_0_));
    InMux I__3518 (
            .O(N__26827),
            .I(N__26824));
    LocalMux I__3517 (
            .O(N__26824),
            .I(N__26821));
    Span12Mux_v I__3516 (
            .O(N__26821),
            .I(N__26818));
    Span12Mux_h I__3515 (
            .O(N__26818),
            .I(N__26815));
    Odrv12 I__3514 (
            .O(N__26815),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_9 ));
    InMux I__3513 (
            .O(N__26812),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ));
    InMux I__3512 (
            .O(N__26809),
            .I(N__26806));
    LocalMux I__3511 (
            .O(N__26806),
            .I(N__26803));
    Span4Mux_v I__3510 (
            .O(N__26803),
            .I(N__26800));
    Sp12to4 I__3509 (
            .O(N__26800),
            .I(N__26797));
    Span12Mux_h I__3508 (
            .O(N__26797),
            .I(N__26794));
    Odrv12 I__3507 (
            .O(N__26794),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_10 ));
    InMux I__3506 (
            .O(N__26791),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ));
    InMux I__3505 (
            .O(N__26788),
            .I(N__26785));
    LocalMux I__3504 (
            .O(N__26785),
            .I(N__26782));
    Span4Mux_v I__3503 (
            .O(N__26782),
            .I(N__26779));
    Sp12to4 I__3502 (
            .O(N__26779),
            .I(N__26776));
    Span12Mux_h I__3501 (
            .O(N__26776),
            .I(N__26773));
    Odrv12 I__3500 (
            .O(N__26773),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_11 ));
    InMux I__3499 (
            .O(N__26770),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ));
    InMux I__3498 (
            .O(N__26767),
            .I(N__26764));
    LocalMux I__3497 (
            .O(N__26764),
            .I(N__26761));
    Span4Mux_v I__3496 (
            .O(N__26761),
            .I(N__26758));
    Sp12to4 I__3495 (
            .O(N__26758),
            .I(N__26755));
    Span12Mux_h I__3494 (
            .O(N__26755),
            .I(N__26752));
    Odrv12 I__3493 (
            .O(N__26752),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_12 ));
    InMux I__3492 (
            .O(N__26749),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ));
    InMux I__3491 (
            .O(N__26746),
            .I(N__26743));
    LocalMux I__3490 (
            .O(N__26743),
            .I(N__26740));
    Span4Mux_v I__3489 (
            .O(N__26740),
            .I(N__26737));
    Sp12to4 I__3488 (
            .O(N__26737),
            .I(N__26734));
    Span12Mux_h I__3487 (
            .O(N__26734),
            .I(N__26731));
    Odrv12 I__3486 (
            .O(N__26731),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_13 ));
    InMux I__3485 (
            .O(N__26728),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ));
    InMux I__3484 (
            .O(N__26725),
            .I(N__26722));
    LocalMux I__3483 (
            .O(N__26722),
            .I(N__26719));
    Span4Mux_v I__3482 (
            .O(N__26719),
            .I(N__26716));
    Sp12to4 I__3481 (
            .O(N__26716),
            .I(N__26713));
    Span12Mux_h I__3480 (
            .O(N__26713),
            .I(N__26710));
    Odrv12 I__3479 (
            .O(N__26710),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_14 ));
    InMux I__3478 (
            .O(N__26707),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ));
    InMux I__3477 (
            .O(N__26704),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ));
    InMux I__3476 (
            .O(N__26701),
            .I(N__26698));
    LocalMux I__3475 (
            .O(N__26698),
            .I(N__26695));
    Span4Mux_v I__3474 (
            .O(N__26695),
            .I(N__26692));
    Sp12to4 I__3473 (
            .O(N__26692),
            .I(N__26689));
    Span12Mux_h I__3472 (
            .O(N__26689),
            .I(N__26686));
    Odrv12 I__3471 (
            .O(N__26686),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_0 ));
    CascadeMux I__3470 (
            .O(N__26683),
            .I(N__26680));
    InMux I__3469 (
            .O(N__26680),
            .I(N__26677));
    LocalMux I__3468 (
            .O(N__26677),
            .I(N__26674));
    Span4Mux_v I__3467 (
            .O(N__26674),
            .I(N__26671));
    Sp12to4 I__3466 (
            .O(N__26671),
            .I(N__26668));
    Span12Mux_v I__3465 (
            .O(N__26668),
            .I(N__26665));
    Odrv12 I__3464 (
            .O(N__26665),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_15 ));
    InMux I__3463 (
            .O(N__26662),
            .I(N__26659));
    LocalMux I__3462 (
            .O(N__26659),
            .I(N__26656));
    Span12Mux_v I__3461 (
            .O(N__26656),
            .I(N__26653));
    Span12Mux_h I__3460 (
            .O(N__26653),
            .I(N__26650));
    Odrv12 I__3459 (
            .O(N__26650),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_1 ));
    CascadeMux I__3458 (
            .O(N__26647),
            .I(N__26644));
    InMux I__3457 (
            .O(N__26644),
            .I(N__26641));
    LocalMux I__3456 (
            .O(N__26641),
            .I(N__26638));
    Span12Mux_s11_v I__3455 (
            .O(N__26638),
            .I(N__26635));
    Span12Mux_v I__3454 (
            .O(N__26635),
            .I(N__26632));
    Odrv12 I__3453 (
            .O(N__26632),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_16 ));
    InMux I__3452 (
            .O(N__26629),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ));
    InMux I__3451 (
            .O(N__26626),
            .I(N__26623));
    LocalMux I__3450 (
            .O(N__26623),
            .I(N__26620));
    Span12Mux_h I__3449 (
            .O(N__26620),
            .I(N__26617));
    Span12Mux_h I__3448 (
            .O(N__26617),
            .I(N__26614));
    Odrv12 I__3447 (
            .O(N__26614),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_2 ));
    CascadeMux I__3446 (
            .O(N__26611),
            .I(N__26608));
    InMux I__3445 (
            .O(N__26608),
            .I(N__26605));
    LocalMux I__3444 (
            .O(N__26605),
            .I(N__26602));
    Span4Mux_v I__3443 (
            .O(N__26602),
            .I(N__26599));
    Span4Mux_h I__3442 (
            .O(N__26599),
            .I(N__26596));
    Span4Mux_h I__3441 (
            .O(N__26596),
            .I(N__26593));
    Span4Mux_v I__3440 (
            .O(N__26593),
            .I(N__26590));
    Span4Mux_v I__3439 (
            .O(N__26590),
            .I(N__26587));
    Odrv4 I__3438 (
            .O(N__26587),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_17 ));
    InMux I__3437 (
            .O(N__26584),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ));
    InMux I__3436 (
            .O(N__26581),
            .I(N__26578));
    LocalMux I__3435 (
            .O(N__26578),
            .I(N__26575));
    Span4Mux_v I__3434 (
            .O(N__26575),
            .I(N__26572));
    Sp12to4 I__3433 (
            .O(N__26572),
            .I(N__26569));
    Span12Mux_h I__3432 (
            .O(N__26569),
            .I(N__26566));
    Odrv12 I__3431 (
            .O(N__26566),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_3 ));
    CascadeMux I__3430 (
            .O(N__26563),
            .I(N__26560));
    InMux I__3429 (
            .O(N__26560),
            .I(N__26557));
    LocalMux I__3428 (
            .O(N__26557),
            .I(N__26554));
    Span12Mux_h I__3427 (
            .O(N__26554),
            .I(N__26551));
    Span12Mux_v I__3426 (
            .O(N__26551),
            .I(N__26548));
    Odrv12 I__3425 (
            .O(N__26548),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_1_18 ));
    InMux I__3424 (
            .O(N__26545),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ));
    InMux I__3423 (
            .O(N__26542),
            .I(N__26539));
    LocalMux I__3422 (
            .O(N__26539),
            .I(N__26536));
    Span4Mux_v I__3421 (
            .O(N__26536),
            .I(N__26533));
    Sp12to4 I__3420 (
            .O(N__26533),
            .I(N__26530));
    Span12Mux_h I__3419 (
            .O(N__26530),
            .I(N__26527));
    Odrv12 I__3418 (
            .O(N__26527),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_4 ));
    InMux I__3417 (
            .O(N__26524),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ));
    InMux I__3416 (
            .O(N__26521),
            .I(N__26518));
    LocalMux I__3415 (
            .O(N__26518),
            .I(N__26515));
    Span4Mux_v I__3414 (
            .O(N__26515),
            .I(N__26512));
    Sp12to4 I__3413 (
            .O(N__26512),
            .I(N__26509));
    Span12Mux_h I__3412 (
            .O(N__26509),
            .I(N__26506));
    Odrv12 I__3411 (
            .O(N__26506),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_5 ));
    InMux I__3410 (
            .O(N__26503),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ));
    InMux I__3409 (
            .O(N__26500),
            .I(N__26497));
    LocalMux I__3408 (
            .O(N__26497),
            .I(N__26494));
    Span4Mux_v I__3407 (
            .O(N__26494),
            .I(N__26491));
    Sp12to4 I__3406 (
            .O(N__26491),
            .I(N__26488));
    Span12Mux_h I__3405 (
            .O(N__26488),
            .I(N__26485));
    Odrv12 I__3404 (
            .O(N__26485),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_6 ));
    InMux I__3403 (
            .O(N__26482),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ));
    InMux I__3402 (
            .O(N__26479),
            .I(N__26476));
    LocalMux I__3401 (
            .O(N__26476),
            .I(N__26473));
    Span4Mux_v I__3400 (
            .O(N__26473),
            .I(N__26470));
    Sp12to4 I__3399 (
            .O(N__26470),
            .I(N__26467));
    Span12Mux_h I__3398 (
            .O(N__26467),
            .I(N__26464));
    Odrv12 I__3397 (
            .O(N__26464),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_2_7 ));
    InMux I__3396 (
            .O(N__26461),
            .I(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ));
    InMux I__3395 (
            .O(N__26458),
            .I(N__26452));
    InMux I__3394 (
            .O(N__26457),
            .I(N__26452));
    LocalMux I__3393 (
            .O(N__26452),
            .I(N__26448));
    InMux I__3392 (
            .O(N__26451),
            .I(N__26445));
    Span4Mux_v I__3391 (
            .O(N__26448),
            .I(N__26442));
    LocalMux I__3390 (
            .O(N__26445),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ));
    Odrv4 I__3389 (
            .O(N__26442),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ));
    InMux I__3388 (
            .O(N__26437),
            .I(bfn_8_20_0_));
    CascadeMux I__3387 (
            .O(N__26434),
            .I(N__26430));
    CascadeMux I__3386 (
            .O(N__26433),
            .I(N__26427));
    InMux I__3385 (
            .O(N__26430),
            .I(N__26422));
    InMux I__3384 (
            .O(N__26427),
            .I(N__26422));
    LocalMux I__3383 (
            .O(N__26422),
            .I(N__26418));
    InMux I__3382 (
            .O(N__26421),
            .I(N__26415));
    Span4Mux_v I__3381 (
            .O(N__26418),
            .I(N__26412));
    LocalMux I__3380 (
            .O(N__26415),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ));
    Odrv4 I__3379 (
            .O(N__26412),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ));
    InMux I__3378 (
            .O(N__26407),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_24 ));
    CascadeMux I__3377 (
            .O(N__26404),
            .I(N__26400));
    CascadeMux I__3376 (
            .O(N__26403),
            .I(N__26397));
    InMux I__3375 (
            .O(N__26400),
            .I(N__26392));
    InMux I__3374 (
            .O(N__26397),
            .I(N__26392));
    LocalMux I__3373 (
            .O(N__26392),
            .I(N__26388));
    InMux I__3372 (
            .O(N__26391),
            .I(N__26385));
    Span4Mux_h I__3371 (
            .O(N__26388),
            .I(N__26382));
    LocalMux I__3370 (
            .O(N__26385),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ));
    Odrv4 I__3369 (
            .O(N__26382),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ));
    InMux I__3368 (
            .O(N__26377),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_25 ));
    InMux I__3367 (
            .O(N__26374),
            .I(N__26368));
    InMux I__3366 (
            .O(N__26373),
            .I(N__26368));
    LocalMux I__3365 (
            .O(N__26368),
            .I(N__26364));
    InMux I__3364 (
            .O(N__26367),
            .I(N__26361));
    Span4Mux_h I__3363 (
            .O(N__26364),
            .I(N__26358));
    LocalMux I__3362 (
            .O(N__26361),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    Odrv4 I__3361 (
            .O(N__26358),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ));
    InMux I__3360 (
            .O(N__26353),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_26 ));
    InMux I__3359 (
            .O(N__26350),
            .I(N__26345));
    InMux I__3358 (
            .O(N__26349),
            .I(N__26342));
    InMux I__3357 (
            .O(N__26348),
            .I(N__26339));
    LocalMux I__3356 (
            .O(N__26345),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    LocalMux I__3355 (
            .O(N__26342),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    LocalMux I__3354 (
            .O(N__26339),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ));
    InMux I__3353 (
            .O(N__26332),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_27 ));
    InMux I__3352 (
            .O(N__26329),
            .I(N__26324));
    InMux I__3351 (
            .O(N__26328),
            .I(N__26319));
    InMux I__3350 (
            .O(N__26327),
            .I(N__26319));
    LocalMux I__3349 (
            .O(N__26324),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    LocalMux I__3348 (
            .O(N__26319),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ));
    InMux I__3347 (
            .O(N__26314),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_28 ));
    InMux I__3346 (
            .O(N__26311),
            .I(N__26306));
    InMux I__3345 (
            .O(N__26310),
            .I(N__26301));
    InMux I__3344 (
            .O(N__26309),
            .I(N__26301));
    LocalMux I__3343 (
            .O(N__26306),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    LocalMux I__3342 (
            .O(N__26301),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ));
    InMux I__3341 (
            .O(N__26296),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_29 ));
    InMux I__3340 (
            .O(N__26293),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_30 ));
    InMux I__3339 (
            .O(N__26290),
            .I(N__26285));
    InMux I__3338 (
            .O(N__26289),
            .I(N__26282));
    InMux I__3337 (
            .O(N__26288),
            .I(N__26279));
    LocalMux I__3336 (
            .O(N__26285),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    LocalMux I__3335 (
            .O(N__26282),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    LocalMux I__3334 (
            .O(N__26279),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ));
    CEMux I__3333 (
            .O(N__26272),
            .I(N__26260));
    CEMux I__3332 (
            .O(N__26271),
            .I(N__26260));
    CEMux I__3331 (
            .O(N__26270),
            .I(N__26260));
    CEMux I__3330 (
            .O(N__26269),
            .I(N__26260));
    GlobalMux I__3329 (
            .O(N__26260),
            .I(N__26257));
    gio2CtrlBuf I__3328 (
            .O(N__26257),
            .I(\phase_controller_inst2.stoper_tr.un2_start_0_g ));
    InMux I__3327 (
            .O(N__26254),
            .I(N__26250));
    InMux I__3326 (
            .O(N__26253),
            .I(N__26247));
    LocalMux I__3325 (
            .O(N__26250),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ));
    LocalMux I__3324 (
            .O(N__26247),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ));
    InMux I__3323 (
            .O(N__26242),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_14 ));
    InMux I__3322 (
            .O(N__26239),
            .I(N__26233));
    InMux I__3321 (
            .O(N__26238),
            .I(N__26233));
    LocalMux I__3320 (
            .O(N__26233),
            .I(N__26229));
    InMux I__3319 (
            .O(N__26232),
            .I(N__26226));
    Span4Mux_v I__3318 (
            .O(N__26229),
            .I(N__26223));
    LocalMux I__3317 (
            .O(N__26226),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ));
    Odrv4 I__3316 (
            .O(N__26223),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ));
    InMux I__3315 (
            .O(N__26218),
            .I(bfn_8_19_0_));
    CascadeMux I__3314 (
            .O(N__26215),
            .I(N__26211));
    CascadeMux I__3313 (
            .O(N__26214),
            .I(N__26208));
    InMux I__3312 (
            .O(N__26211),
            .I(N__26203));
    InMux I__3311 (
            .O(N__26208),
            .I(N__26203));
    LocalMux I__3310 (
            .O(N__26203),
            .I(N__26199));
    InMux I__3309 (
            .O(N__26202),
            .I(N__26196));
    Span4Mux_v I__3308 (
            .O(N__26199),
            .I(N__26193));
    LocalMux I__3307 (
            .O(N__26196),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ));
    Odrv4 I__3306 (
            .O(N__26193),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ));
    InMux I__3305 (
            .O(N__26188),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_16 ));
    InMux I__3304 (
            .O(N__26185),
            .I(N__26179));
    InMux I__3303 (
            .O(N__26184),
            .I(N__26179));
    LocalMux I__3302 (
            .O(N__26179),
            .I(N__26175));
    InMux I__3301 (
            .O(N__26178),
            .I(N__26172));
    Span4Mux_h I__3300 (
            .O(N__26175),
            .I(N__26169));
    LocalMux I__3299 (
            .O(N__26172),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ));
    Odrv4 I__3298 (
            .O(N__26169),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ));
    InMux I__3297 (
            .O(N__26164),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_17 ));
    InMux I__3296 (
            .O(N__26161),
            .I(N__26155));
    InMux I__3295 (
            .O(N__26160),
            .I(N__26155));
    LocalMux I__3294 (
            .O(N__26155),
            .I(N__26151));
    InMux I__3293 (
            .O(N__26154),
            .I(N__26148));
    Span4Mux_h I__3292 (
            .O(N__26151),
            .I(N__26145));
    LocalMux I__3291 (
            .O(N__26148),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ));
    Odrv4 I__3290 (
            .O(N__26145),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ));
    InMux I__3289 (
            .O(N__26140),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_18 ));
    CascadeMux I__3288 (
            .O(N__26137),
            .I(N__26133));
    CascadeMux I__3287 (
            .O(N__26136),
            .I(N__26130));
    InMux I__3286 (
            .O(N__26133),
            .I(N__26124));
    InMux I__3285 (
            .O(N__26130),
            .I(N__26124));
    InMux I__3284 (
            .O(N__26129),
            .I(N__26121));
    LocalMux I__3283 (
            .O(N__26124),
            .I(N__26118));
    LocalMux I__3282 (
            .O(N__26121),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ));
    Odrv4 I__3281 (
            .O(N__26118),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ));
    InMux I__3280 (
            .O(N__26113),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_19 ));
    InMux I__3279 (
            .O(N__26110),
            .I(N__26103));
    InMux I__3278 (
            .O(N__26109),
            .I(N__26103));
    InMux I__3277 (
            .O(N__26108),
            .I(N__26100));
    LocalMux I__3276 (
            .O(N__26103),
            .I(N__26097));
    LocalMux I__3275 (
            .O(N__26100),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ));
    Odrv4 I__3274 (
            .O(N__26097),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ));
    InMux I__3273 (
            .O(N__26092),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_20 ));
    CascadeMux I__3272 (
            .O(N__26089),
            .I(N__26085));
    CascadeMux I__3271 (
            .O(N__26088),
            .I(N__26082));
    InMux I__3270 (
            .O(N__26085),
            .I(N__26077));
    InMux I__3269 (
            .O(N__26082),
            .I(N__26077));
    LocalMux I__3268 (
            .O(N__26077),
            .I(N__26073));
    InMux I__3267 (
            .O(N__26076),
            .I(N__26070));
    Span4Mux_h I__3266 (
            .O(N__26073),
            .I(N__26067));
    LocalMux I__3265 (
            .O(N__26070),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ));
    Odrv4 I__3264 (
            .O(N__26067),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ));
    InMux I__3263 (
            .O(N__26062),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_21 ));
    InMux I__3262 (
            .O(N__26059),
            .I(N__26053));
    InMux I__3261 (
            .O(N__26058),
            .I(N__26053));
    LocalMux I__3260 (
            .O(N__26053),
            .I(N__26049));
    InMux I__3259 (
            .O(N__26052),
            .I(N__26046));
    Span4Mux_h I__3258 (
            .O(N__26049),
            .I(N__26043));
    LocalMux I__3257 (
            .O(N__26046),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ));
    Odrv4 I__3256 (
            .O(N__26043),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ));
    InMux I__3255 (
            .O(N__26038),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_22 ));
    InMux I__3254 (
            .O(N__26035),
            .I(N__26031));
    InMux I__3253 (
            .O(N__26034),
            .I(N__26028));
    LocalMux I__3252 (
            .O(N__26031),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ));
    LocalMux I__3251 (
            .O(N__26028),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ));
    InMux I__3250 (
            .O(N__26023),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_6 ));
    InMux I__3249 (
            .O(N__26020),
            .I(N__26016));
    InMux I__3248 (
            .O(N__26019),
            .I(N__26013));
    LocalMux I__3247 (
            .O(N__26016),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ));
    LocalMux I__3246 (
            .O(N__26013),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ));
    InMux I__3245 (
            .O(N__26008),
            .I(bfn_8_18_0_));
    InMux I__3244 (
            .O(N__26005),
            .I(N__26001));
    InMux I__3243 (
            .O(N__26004),
            .I(N__25998));
    LocalMux I__3242 (
            .O(N__26001),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ));
    LocalMux I__3241 (
            .O(N__25998),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ));
    InMux I__3240 (
            .O(N__25993),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_8 ));
    InMux I__3239 (
            .O(N__25990),
            .I(N__25986));
    InMux I__3238 (
            .O(N__25989),
            .I(N__25983));
    LocalMux I__3237 (
            .O(N__25986),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ));
    LocalMux I__3236 (
            .O(N__25983),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ));
    InMux I__3235 (
            .O(N__25978),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_9 ));
    InMux I__3234 (
            .O(N__25975),
            .I(N__25971));
    InMux I__3233 (
            .O(N__25974),
            .I(N__25968));
    LocalMux I__3232 (
            .O(N__25971),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ));
    LocalMux I__3231 (
            .O(N__25968),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ));
    InMux I__3230 (
            .O(N__25963),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_10 ));
    InMux I__3229 (
            .O(N__25960),
            .I(N__25956));
    InMux I__3228 (
            .O(N__25959),
            .I(N__25953));
    LocalMux I__3227 (
            .O(N__25956),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ));
    LocalMux I__3226 (
            .O(N__25953),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ));
    InMux I__3225 (
            .O(N__25948),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_11 ));
    InMux I__3224 (
            .O(N__25945),
            .I(N__25941));
    InMux I__3223 (
            .O(N__25944),
            .I(N__25938));
    LocalMux I__3222 (
            .O(N__25941),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ));
    LocalMux I__3221 (
            .O(N__25938),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ));
    InMux I__3220 (
            .O(N__25933),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_12 ));
    InMux I__3219 (
            .O(N__25930),
            .I(N__25926));
    InMux I__3218 (
            .O(N__25929),
            .I(N__25923));
    LocalMux I__3217 (
            .O(N__25926),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ));
    LocalMux I__3216 (
            .O(N__25923),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ));
    InMux I__3215 (
            .O(N__25918),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_13 ));
    InMux I__3214 (
            .O(N__25915),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ));
    CascadeMux I__3213 (
            .O(N__25912),
            .I(N__25908));
    InMux I__3212 (
            .O(N__25911),
            .I(N__25905));
    InMux I__3211 (
            .O(N__25908),
            .I(N__25902));
    LocalMux I__3210 (
            .O(N__25905),
            .I(N__25897));
    LocalMux I__3209 (
            .O(N__25902),
            .I(N__25897));
    Odrv4 I__3208 (
            .O(N__25897),
            .I(\phase_controller_inst2.stoper_tr.counter ));
    InMux I__3207 (
            .O(N__25894),
            .I(N__25890));
    InMux I__3206 (
            .O(N__25893),
            .I(N__25887));
    LocalMux I__3205 (
            .O(N__25890),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ));
    LocalMux I__3204 (
            .O(N__25887),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ));
    InMux I__3203 (
            .O(N__25882),
            .I(N__25878));
    InMux I__3202 (
            .O(N__25881),
            .I(N__25875));
    LocalMux I__3201 (
            .O(N__25878),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ));
    LocalMux I__3200 (
            .O(N__25875),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ));
    InMux I__3199 (
            .O(N__25870),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_0 ));
    InMux I__3198 (
            .O(N__25867),
            .I(N__25863));
    InMux I__3197 (
            .O(N__25866),
            .I(N__25860));
    LocalMux I__3196 (
            .O(N__25863),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ));
    LocalMux I__3195 (
            .O(N__25860),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ));
    InMux I__3194 (
            .O(N__25855),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_1 ));
    InMux I__3193 (
            .O(N__25852),
            .I(N__25848));
    InMux I__3192 (
            .O(N__25851),
            .I(N__25845));
    LocalMux I__3191 (
            .O(N__25848),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ));
    LocalMux I__3190 (
            .O(N__25845),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ));
    InMux I__3189 (
            .O(N__25840),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_2 ));
    InMux I__3188 (
            .O(N__25837),
            .I(N__25833));
    InMux I__3187 (
            .O(N__25836),
            .I(N__25830));
    LocalMux I__3186 (
            .O(N__25833),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ));
    LocalMux I__3185 (
            .O(N__25830),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ));
    InMux I__3184 (
            .O(N__25825),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_3 ));
    InMux I__3183 (
            .O(N__25822),
            .I(N__25818));
    InMux I__3182 (
            .O(N__25821),
            .I(N__25815));
    LocalMux I__3181 (
            .O(N__25818),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ));
    LocalMux I__3180 (
            .O(N__25815),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ));
    InMux I__3179 (
            .O(N__25810),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_4 ));
    InMux I__3178 (
            .O(N__25807),
            .I(N__25803));
    InMux I__3177 (
            .O(N__25806),
            .I(N__25800));
    LocalMux I__3176 (
            .O(N__25803),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ));
    LocalMux I__3175 (
            .O(N__25800),
            .I(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ));
    InMux I__3174 (
            .O(N__25795),
            .I(\phase_controller_inst2.stoper_tr.counter_cry_5 ));
    InMux I__3173 (
            .O(N__25792),
            .I(N__25789));
    LocalMux I__3172 (
            .O(N__25789),
            .I(N__25785));
    InMux I__3171 (
            .O(N__25788),
            .I(N__25782));
    Span4Mux_v I__3170 (
            .O(N__25785),
            .I(N__25777));
    LocalMux I__3169 (
            .O(N__25782),
            .I(N__25777));
    Odrv4 I__3168 (
            .O(N__25777),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_19));
    InMux I__3167 (
            .O(N__25774),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ));
    InMux I__3166 (
            .O(N__25771),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ));
    InMux I__3165 (
            .O(N__25768),
            .I(N__25765));
    LocalMux I__3164 (
            .O(N__25765),
            .I(N__25762));
    Span4Mux_h I__3163 (
            .O(N__25762),
            .I(N__25758));
    InMux I__3162 (
            .O(N__25761),
            .I(N__25755));
    Odrv4 I__3161 (
            .O(N__25758),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_21));
    LocalMux I__3160 (
            .O(N__25755),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_21));
    InMux I__3159 (
            .O(N__25750),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ));
    InMux I__3158 (
            .O(N__25747),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ));
    InMux I__3157 (
            .O(N__25744),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ));
    InMux I__3156 (
            .O(N__25741),
            .I(bfn_8_16_0_));
    InMux I__3155 (
            .O(N__25738),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ));
    InMux I__3154 (
            .O(N__25735),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ));
    InMux I__3153 (
            .O(N__25732),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ));
    InMux I__3152 (
            .O(N__25729),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ));
    InMux I__3151 (
            .O(N__25726),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ));
    InMux I__3150 (
            .O(N__25723),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ));
    InMux I__3149 (
            .O(N__25720),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ));
    InMux I__3148 (
            .O(N__25717),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ));
    InMux I__3147 (
            .O(N__25714),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ));
    InMux I__3146 (
            .O(N__25711),
            .I(N__25708));
    LocalMux I__3145 (
            .O(N__25708),
            .I(N__25705));
    Span4Mux_v I__3144 (
            .O(N__25705),
            .I(N__25701));
    InMux I__3143 (
            .O(N__25704),
            .I(N__25698));
    Span4Mux_h I__3142 (
            .O(N__25701),
            .I(N__25695));
    LocalMux I__3141 (
            .O(N__25698),
            .I(N__25692));
    Odrv4 I__3140 (
            .O(N__25695),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_16));
    Odrv12 I__3139 (
            .O(N__25692),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_16));
    InMux I__3138 (
            .O(N__25687),
            .I(bfn_8_15_0_));
    InMux I__3137 (
            .O(N__25684),
            .I(N__25681));
    LocalMux I__3136 (
            .O(N__25681),
            .I(N__25677));
    InMux I__3135 (
            .O(N__25680),
            .I(N__25674));
    Span4Mux_v I__3134 (
            .O(N__25677),
            .I(N__25671));
    LocalMux I__3133 (
            .O(N__25674),
            .I(N__25668));
    Odrv4 I__3132 (
            .O(N__25671),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_17));
    Odrv12 I__3131 (
            .O(N__25668),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_17));
    InMux I__3130 (
            .O(N__25663),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ));
    InMux I__3129 (
            .O(N__25660),
            .I(N__25657));
    LocalMux I__3128 (
            .O(N__25657),
            .I(N__25653));
    InMux I__3127 (
            .O(N__25656),
            .I(N__25650));
    Span4Mux_v I__3126 (
            .O(N__25653),
            .I(N__25645));
    LocalMux I__3125 (
            .O(N__25650),
            .I(N__25645));
    Odrv4 I__3124 (
            .O(N__25645),
            .I(phase_controller_inst1_stoper_tr_target_ticks_1_i_18));
    InMux I__3123 (
            .O(N__25642),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ));
    InMux I__3122 (
            .O(N__25639),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ));
    InMux I__3121 (
            .O(N__25636),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ));
    InMux I__3120 (
            .O(N__25633),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ));
    InMux I__3119 (
            .O(N__25630),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ));
    InMux I__3118 (
            .O(N__25627),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ));
    InMux I__3117 (
            .O(N__25624),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ));
    InMux I__3116 (
            .O(N__25621),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ));
    InMux I__3115 (
            .O(N__25618),
            .I(bfn_8_14_0_));
    InMux I__3114 (
            .O(N__25615),
            .I(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ));
    InMux I__3113 (
            .O(N__25612),
            .I(N__25608));
    InMux I__3112 (
            .O(N__25611),
            .I(N__25605));
    LocalMux I__3111 (
            .O(N__25608),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    LocalMux I__3110 (
            .O(N__25605),
            .I(elapsed_time_ns_1_RNIT6OBB_0_10));
    InMux I__3109 (
            .O(N__25600),
            .I(N__25597));
    LocalMux I__3108 (
            .O(N__25597),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26));
    CascadeMux I__3107 (
            .O(N__25594),
            .I(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_));
    InMux I__3106 (
            .O(N__25591),
            .I(N__25587));
    InMux I__3105 (
            .O(N__25590),
            .I(N__25584));
    LocalMux I__3104 (
            .O(N__25587),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    LocalMux I__3103 (
            .O(N__25584),
            .I(elapsed_time_ns_1_RNI2COBB_0_15));
    InMux I__3102 (
            .O(N__25579),
            .I(N__25576));
    LocalMux I__3101 (
            .O(N__25576),
            .I(elapsed_time_ns_1_RNILK91B_0_9));
    CascadeMux I__3100 (
            .O(N__25573),
            .I(elapsed_time_ns_1_RNILK91B_0_9_cascade_));
    InMux I__3099 (
            .O(N__25570),
            .I(N__25566));
    InMux I__3098 (
            .O(N__25569),
            .I(N__25563));
    LocalMux I__3097 (
            .O(N__25566),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    LocalMux I__3096 (
            .O(N__25563),
            .I(elapsed_time_ns_1_RNI1BOBB_0_14));
    InMux I__3095 (
            .O(N__25558),
            .I(N__25555));
    LocalMux I__3094 (
            .O(N__25555),
            .I(\phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ));
    CascadeMux I__3093 (
            .O(N__25552),
            .I(N__25549));
    InMux I__3092 (
            .O(N__25549),
            .I(N__25544));
    InMux I__3091 (
            .O(N__25548),
            .I(N__25541));
    InMux I__3090 (
            .O(N__25547),
            .I(N__25538));
    LocalMux I__3089 (
            .O(N__25544),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3088 (
            .O(N__25541),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    LocalMux I__3087 (
            .O(N__25538),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ));
    InMux I__3086 (
            .O(N__25531),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ));
    CascadeMux I__3085 (
            .O(N__25528),
            .I(N__25525));
    InMux I__3084 (
            .O(N__25525),
            .I(N__25520));
    InMux I__3083 (
            .O(N__25524),
            .I(N__25517));
    InMux I__3082 (
            .O(N__25523),
            .I(N__25514));
    LocalMux I__3081 (
            .O(N__25520),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3080 (
            .O(N__25517),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    LocalMux I__3079 (
            .O(N__25514),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ));
    InMux I__3078 (
            .O(N__25507),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ));
    CascadeMux I__3077 (
            .O(N__25504),
            .I(N__25501));
    InMux I__3076 (
            .O(N__25501),
            .I(N__25496));
    InMux I__3075 (
            .O(N__25500),
            .I(N__25493));
    InMux I__3074 (
            .O(N__25499),
            .I(N__25490));
    LocalMux I__3073 (
            .O(N__25496),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3072 (
            .O(N__25493),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    LocalMux I__3071 (
            .O(N__25490),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ));
    InMux I__3070 (
            .O(N__25483),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ));
    CascadeMux I__3069 (
            .O(N__25480),
            .I(N__25477));
    InMux I__3068 (
            .O(N__25477),
            .I(N__25472));
    InMux I__3067 (
            .O(N__25476),
            .I(N__25469));
    InMux I__3066 (
            .O(N__25475),
            .I(N__25466));
    LocalMux I__3065 (
            .O(N__25472),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3064 (
            .O(N__25469),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    LocalMux I__3063 (
            .O(N__25466),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ));
    InMux I__3062 (
            .O(N__25459),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ));
    CascadeMux I__3061 (
            .O(N__25456),
            .I(N__25453));
    InMux I__3060 (
            .O(N__25453),
            .I(N__25448));
    InMux I__3059 (
            .O(N__25452),
            .I(N__25445));
    InMux I__3058 (
            .O(N__25451),
            .I(N__25442));
    LocalMux I__3057 (
            .O(N__25448),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3056 (
            .O(N__25445),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    LocalMux I__3055 (
            .O(N__25442),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ));
    InMux I__3054 (
            .O(N__25435),
            .I(bfn_8_11_0_));
    CascadeMux I__3053 (
            .O(N__25432),
            .I(N__25429));
    InMux I__3052 (
            .O(N__25429),
            .I(N__25424));
    InMux I__3051 (
            .O(N__25428),
            .I(N__25421));
    InMux I__3050 (
            .O(N__25427),
            .I(N__25418));
    LocalMux I__3049 (
            .O(N__25424),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3048 (
            .O(N__25421),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    LocalMux I__3047 (
            .O(N__25418),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ));
    InMux I__3046 (
            .O(N__25411),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ));
    InMux I__3045 (
            .O(N__25408),
            .I(N__25404));
    InMux I__3044 (
            .O(N__25407),
            .I(N__25401));
    LocalMux I__3043 (
            .O(N__25404),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    LocalMux I__3042 (
            .O(N__25401),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ));
    CascadeMux I__3041 (
            .O(N__25396),
            .I(N__25393));
    InMux I__3040 (
            .O(N__25393),
            .I(N__25388));
    InMux I__3039 (
            .O(N__25392),
            .I(N__25385));
    InMux I__3038 (
            .O(N__25391),
            .I(N__25382));
    LocalMux I__3037 (
            .O(N__25388),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3036 (
            .O(N__25385),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    LocalMux I__3035 (
            .O(N__25382),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ));
    InMux I__3034 (
            .O(N__25375),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ));
    InMux I__3033 (
            .O(N__25372),
            .I(N__25368));
    InMux I__3032 (
            .O(N__25371),
            .I(N__25365));
    LocalMux I__3031 (
            .O(N__25368),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    LocalMux I__3030 (
            .O(N__25365),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ));
    CascadeMux I__3029 (
            .O(N__25360),
            .I(N__25357));
    InMux I__3028 (
            .O(N__25357),
            .I(N__25352));
    InMux I__3027 (
            .O(N__25356),
            .I(N__25349));
    InMux I__3026 (
            .O(N__25355),
            .I(N__25346));
    LocalMux I__3025 (
            .O(N__25352),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__3024 (
            .O(N__25349),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    LocalMux I__3023 (
            .O(N__25346),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ));
    InMux I__3022 (
            .O(N__25339),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ));
    InMux I__3021 (
            .O(N__25336),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ));
    CascadeMux I__3020 (
            .O(N__25333),
            .I(N__25330));
    InMux I__3019 (
            .O(N__25330),
            .I(N__25325));
    InMux I__3018 (
            .O(N__25329),
            .I(N__25322));
    InMux I__3017 (
            .O(N__25328),
            .I(N__25319));
    LocalMux I__3016 (
            .O(N__25325),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3015 (
            .O(N__25322),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    LocalMux I__3014 (
            .O(N__25319),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ));
    InMux I__3013 (
            .O(N__25312),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ));
    CascadeMux I__3012 (
            .O(N__25309),
            .I(N__25306));
    InMux I__3011 (
            .O(N__25306),
            .I(N__25301));
    InMux I__3010 (
            .O(N__25305),
            .I(N__25298));
    InMux I__3009 (
            .O(N__25304),
            .I(N__25295));
    LocalMux I__3008 (
            .O(N__25301),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3007 (
            .O(N__25298),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    LocalMux I__3006 (
            .O(N__25295),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ));
    InMux I__3005 (
            .O(N__25288),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ));
    CascadeMux I__3004 (
            .O(N__25285),
            .I(N__25282));
    InMux I__3003 (
            .O(N__25282),
            .I(N__25277));
    InMux I__3002 (
            .O(N__25281),
            .I(N__25274));
    InMux I__3001 (
            .O(N__25280),
            .I(N__25271));
    LocalMux I__3000 (
            .O(N__25277),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__2999 (
            .O(N__25274),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    LocalMux I__2998 (
            .O(N__25271),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ));
    InMux I__2997 (
            .O(N__25264),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ));
    CascadeMux I__2996 (
            .O(N__25261),
            .I(N__25258));
    InMux I__2995 (
            .O(N__25258),
            .I(N__25253));
    InMux I__2994 (
            .O(N__25257),
            .I(N__25250));
    InMux I__2993 (
            .O(N__25256),
            .I(N__25247));
    LocalMux I__2992 (
            .O(N__25253),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__2991 (
            .O(N__25250),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    LocalMux I__2990 (
            .O(N__25247),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ));
    InMux I__2989 (
            .O(N__25240),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ));
    CascadeMux I__2988 (
            .O(N__25237),
            .I(N__25234));
    InMux I__2987 (
            .O(N__25234),
            .I(N__25229));
    InMux I__2986 (
            .O(N__25233),
            .I(N__25226));
    InMux I__2985 (
            .O(N__25232),
            .I(N__25223));
    LocalMux I__2984 (
            .O(N__25229),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__2983 (
            .O(N__25226),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    LocalMux I__2982 (
            .O(N__25223),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ));
    InMux I__2981 (
            .O(N__25216),
            .I(bfn_8_10_0_));
    InMux I__2980 (
            .O(N__25213),
            .I(N__25208));
    InMux I__2979 (
            .O(N__25212),
            .I(N__25205));
    InMux I__2978 (
            .O(N__25211),
            .I(N__25202));
    LocalMux I__2977 (
            .O(N__25208),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__2976 (
            .O(N__25205),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    LocalMux I__2975 (
            .O(N__25202),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ));
    InMux I__2974 (
            .O(N__25195),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ));
    CascadeMux I__2973 (
            .O(N__25192),
            .I(N__25189));
    InMux I__2972 (
            .O(N__25189),
            .I(N__25184));
    InMux I__2971 (
            .O(N__25188),
            .I(N__25181));
    InMux I__2970 (
            .O(N__25187),
            .I(N__25178));
    LocalMux I__2969 (
            .O(N__25184),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__2968 (
            .O(N__25181),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    LocalMux I__2967 (
            .O(N__25178),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ));
    InMux I__2966 (
            .O(N__25171),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ));
    CascadeMux I__2965 (
            .O(N__25168),
            .I(N__25163));
    CascadeMux I__2964 (
            .O(N__25167),
            .I(N__25160));
    InMux I__2963 (
            .O(N__25166),
            .I(N__25157));
    InMux I__2962 (
            .O(N__25163),
            .I(N__25152));
    InMux I__2961 (
            .O(N__25160),
            .I(N__25152));
    LocalMux I__2960 (
            .O(N__25157),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    LocalMux I__2959 (
            .O(N__25152),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ));
    InMux I__2958 (
            .O(N__25147),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ));
    InMux I__2957 (
            .O(N__25144),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ));
    CascadeMux I__2956 (
            .O(N__25141),
            .I(N__25136));
    CascadeMux I__2955 (
            .O(N__25140),
            .I(N__25133));
    InMux I__2954 (
            .O(N__25139),
            .I(N__25130));
    InMux I__2953 (
            .O(N__25136),
            .I(N__25125));
    InMux I__2952 (
            .O(N__25133),
            .I(N__25125));
    LocalMux I__2951 (
            .O(N__25130),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    LocalMux I__2950 (
            .O(N__25125),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ));
    InMux I__2949 (
            .O(N__25120),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ));
    CascadeMux I__2948 (
            .O(N__25117),
            .I(N__25114));
    InMux I__2947 (
            .O(N__25114),
            .I(N__25109));
    InMux I__2946 (
            .O(N__25113),
            .I(N__25106));
    InMux I__2945 (
            .O(N__25112),
            .I(N__25103));
    LocalMux I__2944 (
            .O(N__25109),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__2943 (
            .O(N__25106),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    LocalMux I__2942 (
            .O(N__25103),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ));
    InMux I__2941 (
            .O(N__25096),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ));
    CascadeMux I__2940 (
            .O(N__25093),
            .I(N__25090));
    InMux I__2939 (
            .O(N__25090),
            .I(N__25085));
    InMux I__2938 (
            .O(N__25089),
            .I(N__25082));
    InMux I__2937 (
            .O(N__25088),
            .I(N__25079));
    LocalMux I__2936 (
            .O(N__25085),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__2935 (
            .O(N__25082),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    LocalMux I__2934 (
            .O(N__25079),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ));
    InMux I__2933 (
            .O(N__25072),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ));
    CascadeMux I__2932 (
            .O(N__25069),
            .I(N__25066));
    InMux I__2931 (
            .O(N__25066),
            .I(N__25061));
    InMux I__2930 (
            .O(N__25065),
            .I(N__25058));
    InMux I__2929 (
            .O(N__25064),
            .I(N__25055));
    LocalMux I__2928 (
            .O(N__25061),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__2927 (
            .O(N__25058),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    LocalMux I__2926 (
            .O(N__25055),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ));
    InMux I__2925 (
            .O(N__25048),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ));
    CascadeMux I__2924 (
            .O(N__25045),
            .I(N__25042));
    InMux I__2923 (
            .O(N__25042),
            .I(N__25037));
    InMux I__2922 (
            .O(N__25041),
            .I(N__25034));
    InMux I__2921 (
            .O(N__25040),
            .I(N__25031));
    LocalMux I__2920 (
            .O(N__25037),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__2919 (
            .O(N__25034),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    LocalMux I__2918 (
            .O(N__25031),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ));
    InMux I__2917 (
            .O(N__25024),
            .I(bfn_8_9_0_));
    InMux I__2916 (
            .O(N__25021),
            .I(N__25016));
    InMux I__2915 (
            .O(N__25020),
            .I(N__25013));
    InMux I__2914 (
            .O(N__25019),
            .I(N__25010));
    LocalMux I__2913 (
            .O(N__25016),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__2912 (
            .O(N__25013),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    LocalMux I__2911 (
            .O(N__25010),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ));
    InMux I__2910 (
            .O(N__25003),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ));
    CascadeMux I__2909 (
            .O(N__25000),
            .I(N__24997));
    InMux I__2908 (
            .O(N__24997),
            .I(N__24992));
    InMux I__2907 (
            .O(N__24996),
            .I(N__24989));
    InMux I__2906 (
            .O(N__24995),
            .I(N__24986));
    LocalMux I__2905 (
            .O(N__24992),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__2904 (
            .O(N__24989),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    LocalMux I__2903 (
            .O(N__24986),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ));
    InMux I__2902 (
            .O(N__24979),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ));
    CascadeMux I__2901 (
            .O(N__24976),
            .I(N__24971));
    CascadeMux I__2900 (
            .O(N__24975),
            .I(N__24968));
    InMux I__2899 (
            .O(N__24974),
            .I(N__24965));
    InMux I__2898 (
            .O(N__24971),
            .I(N__24960));
    InMux I__2897 (
            .O(N__24968),
            .I(N__24960));
    LocalMux I__2896 (
            .O(N__24965),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    LocalMux I__2895 (
            .O(N__24960),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ));
    InMux I__2894 (
            .O(N__24955),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ));
    InMux I__2893 (
            .O(N__24952),
            .I(N__24949));
    LocalMux I__2892 (
            .O(N__24949),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt30 ));
    CascadeMux I__2891 (
            .O(N__24946),
            .I(N__24943));
    InMux I__2890 (
            .O(N__24943),
            .I(N__24940));
    LocalMux I__2889 (
            .O(N__24940),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ));
    InMux I__2888 (
            .O(N__24937),
            .I(N__24934));
    LocalMux I__2887 (
            .O(N__24934),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt28 ));
    InMux I__2886 (
            .O(N__24931),
            .I(N__24928));
    LocalMux I__2885 (
            .O(N__24928),
            .I(N__24925));
    Glb2LocalMux I__2884 (
            .O(N__24925),
            .I(N__24922));
    GlobalMux I__2883 (
            .O(N__24922),
            .I(clk_12mhz));
    IoInMux I__2882 (
            .O(N__24919),
            .I(N__24916));
    LocalMux I__2881 (
            .O(N__24916),
            .I(N__24913));
    Span4Mux_s0_v I__2880 (
            .O(N__24913),
            .I(N__24910));
    Odrv4 I__2879 (
            .O(N__24910),
            .I(GB_BUFFER_clk_12mhz_THRU_CO));
    InMux I__2878 (
            .O(N__24907),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ));
    InMux I__2877 (
            .O(N__24904),
            .I(N__24899));
    InMux I__2876 (
            .O(N__24903),
            .I(N__24894));
    InMux I__2875 (
            .O(N__24902),
            .I(N__24894));
    LocalMux I__2874 (
            .O(N__24899),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    LocalMux I__2873 (
            .O(N__24894),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ));
    InMux I__2872 (
            .O(N__24889),
            .I(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ));
    CascadeMux I__2871 (
            .O(N__24886),
            .I(N__24883));
    InMux I__2870 (
            .O(N__24883),
            .I(N__24878));
    InMux I__2869 (
            .O(N__24882),
            .I(N__24875));
    InMux I__2868 (
            .O(N__24881),
            .I(N__24872));
    LocalMux I__2867 (
            .O(N__24878),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__2866 (
            .O(N__24875),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    LocalMux I__2865 (
            .O(N__24872),
            .I(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ));
    InMux I__2864 (
            .O(N__24865),
            .I(N__24862));
    LocalMux I__2863 (
            .O(N__24862),
            .I(N__24859));
    Odrv4 I__2862 (
            .O(N__24859),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ));
    CascadeMux I__2861 (
            .O(N__24856),
            .I(N__24853));
    InMux I__2860 (
            .O(N__24853),
            .I(N__24850));
    LocalMux I__2859 (
            .O(N__24850),
            .I(N__24847));
    Odrv12 I__2858 (
            .O(N__24847),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt20 ));
    InMux I__2857 (
            .O(N__24844),
            .I(N__24841));
    LocalMux I__2856 (
            .O(N__24841),
            .I(N__24838));
    Span4Mux_v I__2855 (
            .O(N__24838),
            .I(N__24835));
    Odrv4 I__2854 (
            .O(N__24835),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ));
    CascadeMux I__2853 (
            .O(N__24832),
            .I(N__24829));
    InMux I__2852 (
            .O(N__24829),
            .I(N__24826));
    LocalMux I__2851 (
            .O(N__24826),
            .I(N__24823));
    Odrv4 I__2850 (
            .O(N__24823),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt22 ));
    InMux I__2849 (
            .O(N__24820),
            .I(N__24817));
    LocalMux I__2848 (
            .O(N__24817),
            .I(N__24814));
    Odrv4 I__2847 (
            .O(N__24814),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ));
    CascadeMux I__2846 (
            .O(N__24811),
            .I(N__24808));
    InMux I__2845 (
            .O(N__24808),
            .I(N__24805));
    LocalMux I__2844 (
            .O(N__24805),
            .I(N__24802));
    Odrv4 I__2843 (
            .O(N__24802),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt24 ));
    InMux I__2842 (
            .O(N__24799),
            .I(N__24796));
    LocalMux I__2841 (
            .O(N__24796),
            .I(N__24793));
    Odrv4 I__2840 (
            .O(N__24793),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ));
    CascadeMux I__2839 (
            .O(N__24790),
            .I(N__24787));
    InMux I__2838 (
            .O(N__24787),
            .I(N__24784));
    LocalMux I__2837 (
            .O(N__24784),
            .I(N__24781));
    Span4Mux_h I__2836 (
            .O(N__24781),
            .I(N__24778));
    Odrv4 I__2835 (
            .O(N__24778),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt26 ));
    InMux I__2834 (
            .O(N__24775),
            .I(bfn_7_20_0_));
    CascadeMux I__2833 (
            .O(N__24772),
            .I(N__24769));
    InMux I__2832 (
            .O(N__24769),
            .I(N__24766));
    LocalMux I__2831 (
            .O(N__24766),
            .I(N__24763));
    Odrv4 I__2830 (
            .O(N__24763),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ));
    InMux I__2829 (
            .O(N__24760),
            .I(N__24757));
    LocalMux I__2828 (
            .O(N__24757),
            .I(N__24754));
    Odrv12 I__2827 (
            .O(N__24754),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ));
    CascadeMux I__2826 (
            .O(N__24751),
            .I(N__24748));
    InMux I__2825 (
            .O(N__24748),
            .I(N__24745));
    LocalMux I__2824 (
            .O(N__24745),
            .I(\phase_controller_inst2.stoper_tr.counter_i_10 ));
    CascadeMux I__2823 (
            .O(N__24742),
            .I(N__24739));
    InMux I__2822 (
            .O(N__24739),
            .I(N__24736));
    LocalMux I__2821 (
            .O(N__24736),
            .I(N__24733));
    Odrv4 I__2820 (
            .O(N__24733),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ));
    InMux I__2819 (
            .O(N__24730),
            .I(N__24727));
    LocalMux I__2818 (
            .O(N__24727),
            .I(\phase_controller_inst2.stoper_tr.counter_i_11 ));
    InMux I__2817 (
            .O(N__24724),
            .I(N__24721));
    LocalMux I__2816 (
            .O(N__24721),
            .I(N__24718));
    Odrv4 I__2815 (
            .O(N__24718),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ));
    CascadeMux I__2814 (
            .O(N__24715),
            .I(N__24712));
    InMux I__2813 (
            .O(N__24712),
            .I(N__24709));
    LocalMux I__2812 (
            .O(N__24709),
            .I(\phase_controller_inst2.stoper_tr.counter_i_12 ));
    InMux I__2811 (
            .O(N__24706),
            .I(N__24703));
    LocalMux I__2810 (
            .O(N__24703),
            .I(N__24700));
    Odrv4 I__2809 (
            .O(N__24700),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ));
    CascadeMux I__2808 (
            .O(N__24697),
            .I(N__24694));
    InMux I__2807 (
            .O(N__24694),
            .I(N__24691));
    LocalMux I__2806 (
            .O(N__24691),
            .I(N__24688));
    Odrv4 I__2805 (
            .O(N__24688),
            .I(\phase_controller_inst2.stoper_tr.counter_i_13 ));
    CascadeMux I__2804 (
            .O(N__24685),
            .I(N__24682));
    InMux I__2803 (
            .O(N__24682),
            .I(N__24679));
    LocalMux I__2802 (
            .O(N__24679),
            .I(N__24676));
    Odrv12 I__2801 (
            .O(N__24676),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ));
    InMux I__2800 (
            .O(N__24673),
            .I(N__24670));
    LocalMux I__2799 (
            .O(N__24670),
            .I(\phase_controller_inst2.stoper_tr.counter_i_14 ));
    InMux I__2798 (
            .O(N__24667),
            .I(N__24664));
    LocalMux I__2797 (
            .O(N__24664),
            .I(N__24661));
    Odrv12 I__2796 (
            .O(N__24661),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ));
    CascadeMux I__2795 (
            .O(N__24658),
            .I(N__24655));
    InMux I__2794 (
            .O(N__24655),
            .I(N__24652));
    LocalMux I__2793 (
            .O(N__24652),
            .I(\phase_controller_inst2.stoper_tr.counter_i_15 ));
    InMux I__2792 (
            .O(N__24649),
            .I(N__24646));
    LocalMux I__2791 (
            .O(N__24646),
            .I(N__24643));
    Span4Mux_h I__2790 (
            .O(N__24643),
            .I(N__24640));
    Odrv4 I__2789 (
            .O(N__24640),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt16 ));
    CascadeMux I__2788 (
            .O(N__24637),
            .I(N__24634));
    InMux I__2787 (
            .O(N__24634),
            .I(N__24631));
    LocalMux I__2786 (
            .O(N__24631),
            .I(N__24628));
    Span4Mux_h I__2785 (
            .O(N__24628),
            .I(N__24625));
    Odrv4 I__2784 (
            .O(N__24625),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ));
    InMux I__2783 (
            .O(N__24622),
            .I(N__24619));
    LocalMux I__2782 (
            .O(N__24619),
            .I(N__24616));
    Span4Mux_h I__2781 (
            .O(N__24616),
            .I(N__24613));
    Odrv4 I__2780 (
            .O(N__24613),
            .I(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ));
    CascadeMux I__2779 (
            .O(N__24610),
            .I(N__24607));
    InMux I__2778 (
            .O(N__24607),
            .I(N__24604));
    LocalMux I__2777 (
            .O(N__24604),
            .I(N__24601));
    Span4Mux_v I__2776 (
            .O(N__24601),
            .I(N__24598));
    Odrv4 I__2775 (
            .O(N__24598),
            .I(\phase_controller_inst2.stoper_tr.un6_running_lt18 ));
    CascadeMux I__2774 (
            .O(N__24595),
            .I(N__24592));
    InMux I__2773 (
            .O(N__24592),
            .I(N__24589));
    LocalMux I__2772 (
            .O(N__24589),
            .I(N__24586));
    Odrv4 I__2771 (
            .O(N__24586),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ));
    InMux I__2770 (
            .O(N__24583),
            .I(N__24580));
    LocalMux I__2769 (
            .O(N__24580),
            .I(\phase_controller_inst2.stoper_tr.counter_i_2 ));
    CascadeMux I__2768 (
            .O(N__24577),
            .I(N__24574));
    InMux I__2767 (
            .O(N__24574),
            .I(N__24571));
    LocalMux I__2766 (
            .O(N__24571),
            .I(N__24568));
    Odrv4 I__2765 (
            .O(N__24568),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ));
    InMux I__2764 (
            .O(N__24565),
            .I(N__24562));
    LocalMux I__2763 (
            .O(N__24562),
            .I(\phase_controller_inst2.stoper_tr.counter_i_3 ));
    InMux I__2762 (
            .O(N__24559),
            .I(N__24556));
    LocalMux I__2761 (
            .O(N__24556),
            .I(N__24553));
    Span4Mux_h I__2760 (
            .O(N__24553),
            .I(N__24550));
    Span4Mux_h I__2759 (
            .O(N__24550),
            .I(N__24547));
    Odrv4 I__2758 (
            .O(N__24547),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ));
    CascadeMux I__2757 (
            .O(N__24544),
            .I(N__24541));
    InMux I__2756 (
            .O(N__24541),
            .I(N__24538));
    LocalMux I__2755 (
            .O(N__24538),
            .I(\phase_controller_inst2.stoper_tr.counter_i_4 ));
    CascadeMux I__2754 (
            .O(N__24535),
            .I(N__24532));
    InMux I__2753 (
            .O(N__24532),
            .I(N__24529));
    LocalMux I__2752 (
            .O(N__24529),
            .I(N__24526));
    Odrv12 I__2751 (
            .O(N__24526),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ));
    InMux I__2750 (
            .O(N__24523),
            .I(N__24520));
    LocalMux I__2749 (
            .O(N__24520),
            .I(\phase_controller_inst2.stoper_tr.counter_i_5 ));
    InMux I__2748 (
            .O(N__24517),
            .I(N__24514));
    LocalMux I__2747 (
            .O(N__24514),
            .I(N__24511));
    Odrv4 I__2746 (
            .O(N__24511),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ));
    CascadeMux I__2745 (
            .O(N__24508),
            .I(N__24505));
    InMux I__2744 (
            .O(N__24505),
            .I(N__24502));
    LocalMux I__2743 (
            .O(N__24502),
            .I(\phase_controller_inst2.stoper_tr.counter_i_6 ));
    CascadeMux I__2742 (
            .O(N__24499),
            .I(N__24496));
    InMux I__2741 (
            .O(N__24496),
            .I(N__24493));
    LocalMux I__2740 (
            .O(N__24493),
            .I(N__24490));
    Odrv4 I__2739 (
            .O(N__24490),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ));
    InMux I__2738 (
            .O(N__24487),
            .I(N__24484));
    LocalMux I__2737 (
            .O(N__24484),
            .I(\phase_controller_inst2.stoper_tr.counter_i_7 ));
    InMux I__2736 (
            .O(N__24481),
            .I(N__24478));
    LocalMux I__2735 (
            .O(N__24478),
            .I(N__24475));
    Odrv4 I__2734 (
            .O(N__24475),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ));
    CascadeMux I__2733 (
            .O(N__24472),
            .I(N__24469));
    InMux I__2732 (
            .O(N__24469),
            .I(N__24466));
    LocalMux I__2731 (
            .O(N__24466),
            .I(\phase_controller_inst2.stoper_tr.counter_i_8 ));
    CascadeMux I__2730 (
            .O(N__24463),
            .I(N__24460));
    InMux I__2729 (
            .O(N__24460),
            .I(N__24457));
    LocalMux I__2728 (
            .O(N__24457),
            .I(N__24454));
    Odrv4 I__2727 (
            .O(N__24454),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ));
    InMux I__2726 (
            .O(N__24451),
            .I(N__24448));
    LocalMux I__2725 (
            .O(N__24448),
            .I(\phase_controller_inst2.stoper_tr.counter_i_9 ));
    InMux I__2724 (
            .O(N__24445),
            .I(N__24439));
    InMux I__2723 (
            .O(N__24444),
            .I(N__24439));
    LocalMux I__2722 (
            .O(N__24439),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ));
    InMux I__2721 (
            .O(N__24436),
            .I(N__24430));
    InMux I__2720 (
            .O(N__24435),
            .I(N__24430));
    LocalMux I__2719 (
            .O(N__24430),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ));
    InMux I__2718 (
            .O(N__24427),
            .I(N__24421));
    InMux I__2717 (
            .O(N__24426),
            .I(N__24421));
    LocalMux I__2716 (
            .O(N__24421),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ));
    InMux I__2715 (
            .O(N__24418),
            .I(N__24412));
    InMux I__2714 (
            .O(N__24417),
            .I(N__24412));
    LocalMux I__2713 (
            .O(N__24412),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ));
    InMux I__2712 (
            .O(N__24409),
            .I(N__24406));
    LocalMux I__2711 (
            .O(N__24406),
            .I(N__24403));
    Odrv12 I__2710 (
            .O(N__24403),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ));
    CascadeMux I__2709 (
            .O(N__24400),
            .I(N__24397));
    InMux I__2708 (
            .O(N__24397),
            .I(N__24394));
    LocalMux I__2707 (
            .O(N__24394),
            .I(\phase_controller_inst2.stoper_tr.counter_i_0 ));
    CascadeMux I__2706 (
            .O(N__24391),
            .I(N__24388));
    InMux I__2705 (
            .O(N__24388),
            .I(N__24385));
    LocalMux I__2704 (
            .O(N__24385),
            .I(N__24382));
    Odrv12 I__2703 (
            .O(N__24382),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ));
    InMux I__2702 (
            .O(N__24379),
            .I(N__24376));
    LocalMux I__2701 (
            .O(N__24376),
            .I(\phase_controller_inst2.stoper_tr.counter_i_1 ));
    InMux I__2700 (
            .O(N__24373),
            .I(N__24343));
    InMux I__2699 (
            .O(N__24372),
            .I(N__24343));
    InMux I__2698 (
            .O(N__24371),
            .I(N__24343));
    InMux I__2697 (
            .O(N__24370),
            .I(N__24343));
    InMux I__2696 (
            .O(N__24369),
            .I(N__24330));
    InMux I__2695 (
            .O(N__24368),
            .I(N__24330));
    InMux I__2694 (
            .O(N__24367),
            .I(N__24321));
    InMux I__2693 (
            .O(N__24366),
            .I(N__24321));
    InMux I__2692 (
            .O(N__24365),
            .I(N__24321));
    InMux I__2691 (
            .O(N__24364),
            .I(N__24321));
    InMux I__2690 (
            .O(N__24363),
            .I(N__24312));
    InMux I__2689 (
            .O(N__24362),
            .I(N__24312));
    InMux I__2688 (
            .O(N__24361),
            .I(N__24312));
    InMux I__2687 (
            .O(N__24360),
            .I(N__24312));
    InMux I__2686 (
            .O(N__24359),
            .I(N__24303));
    InMux I__2685 (
            .O(N__24358),
            .I(N__24303));
    InMux I__2684 (
            .O(N__24357),
            .I(N__24303));
    InMux I__2683 (
            .O(N__24356),
            .I(N__24303));
    InMux I__2682 (
            .O(N__24355),
            .I(N__24294));
    InMux I__2681 (
            .O(N__24354),
            .I(N__24294));
    InMux I__2680 (
            .O(N__24353),
            .I(N__24294));
    InMux I__2679 (
            .O(N__24352),
            .I(N__24294));
    LocalMux I__2678 (
            .O(N__24343),
            .I(N__24291));
    InMux I__2677 (
            .O(N__24342),
            .I(N__24282));
    InMux I__2676 (
            .O(N__24341),
            .I(N__24282));
    InMux I__2675 (
            .O(N__24340),
            .I(N__24282));
    InMux I__2674 (
            .O(N__24339),
            .I(N__24282));
    InMux I__2673 (
            .O(N__24338),
            .I(N__24273));
    InMux I__2672 (
            .O(N__24337),
            .I(N__24273));
    InMux I__2671 (
            .O(N__24336),
            .I(N__24273));
    InMux I__2670 (
            .O(N__24335),
            .I(N__24273));
    LocalMux I__2669 (
            .O(N__24330),
            .I(N__24268));
    LocalMux I__2668 (
            .O(N__24321),
            .I(N__24268));
    LocalMux I__2667 (
            .O(N__24312),
            .I(N__24257));
    LocalMux I__2666 (
            .O(N__24303),
            .I(N__24257));
    LocalMux I__2665 (
            .O(N__24294),
            .I(N__24257));
    Span4Mux_h I__2664 (
            .O(N__24291),
            .I(N__24257));
    LocalMux I__2663 (
            .O(N__24282),
            .I(N__24257));
    LocalMux I__2662 (
            .O(N__24273),
            .I(N__24254));
    Span4Mux_v I__2661 (
            .O(N__24268),
            .I(N__24249));
    Span4Mux_v I__2660 (
            .O(N__24257),
            .I(N__24249));
    Odrv12 I__2659 (
            .O(N__24254),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    Odrv4 I__2658 (
            .O(N__24249),
            .I(\delay_measurement_inst.delay_tr_timer.running_i ));
    InMux I__2657 (
            .O(N__24244),
            .I(N__24241));
    LocalMux I__2656 (
            .O(N__24241),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19));
    CascadeMux I__2655 (
            .O(N__24238),
            .I(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_));
    InMux I__2654 (
            .O(N__24235),
            .I(N__24232));
    LocalMux I__2653 (
            .O(N__24232),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29));
    CascadeMux I__2652 (
            .O(N__24229),
            .I(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_));
    InMux I__2651 (
            .O(N__24226),
            .I(N__24223));
    LocalMux I__2650 (
            .O(N__24223),
            .I(elapsed_time_ns_1_RNIJI91B_0_7));
    CascadeMux I__2649 (
            .O(N__24220),
            .I(elapsed_time_ns_1_RNIJI91B_0_7_cascade_));
    InMux I__2648 (
            .O(N__24217),
            .I(N__24213));
    InMux I__2647 (
            .O(N__24216),
            .I(N__24210));
    LocalMux I__2646 (
            .O(N__24213),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    LocalMux I__2645 (
            .O(N__24210),
            .I(elapsed_time_ns_1_RNI1CPBB_0_23));
    InMux I__2644 (
            .O(N__24205),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ));
    InMux I__2643 (
            .O(N__24202),
            .I(bfn_7_10_0_));
    InMux I__2642 (
            .O(N__24199),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ));
    InMux I__2641 (
            .O(N__24196),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ));
    InMux I__2640 (
            .O(N__24193),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ));
    InMux I__2639 (
            .O(N__24190),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ));
    InMux I__2638 (
            .O(N__24187),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ));
    InMux I__2637 (
            .O(N__24184),
            .I(N__24181));
    LocalMux I__2636 (
            .O(N__24181),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27));
    CascadeMux I__2635 (
            .O(N__24178),
            .I(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_));
    InMux I__2634 (
            .O(N__24175),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ));
    InMux I__2633 (
            .O(N__24172),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ));
    InMux I__2632 (
            .O(N__24169),
            .I(bfn_7_9_0_));
    InMux I__2631 (
            .O(N__24166),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ));
    InMux I__2630 (
            .O(N__24163),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ));
    InMux I__2629 (
            .O(N__24160),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ));
    InMux I__2628 (
            .O(N__24157),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ));
    InMux I__2627 (
            .O(N__24154),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ));
    InMux I__2626 (
            .O(N__24151),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ));
    InMux I__2625 (
            .O(N__24148),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ));
    InMux I__2624 (
            .O(N__24145),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ));
    InMux I__2623 (
            .O(N__24142),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ));
    InMux I__2622 (
            .O(N__24139),
            .I(bfn_7_8_0_));
    InMux I__2621 (
            .O(N__24136),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ));
    InMux I__2620 (
            .O(N__24133),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ));
    InMux I__2619 (
            .O(N__24130),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ));
    InMux I__2618 (
            .O(N__24127),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ));
    InMux I__2617 (
            .O(N__24124),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ));
    InMux I__2616 (
            .O(N__24121),
            .I(N__24115));
    InMux I__2615 (
            .O(N__24120),
            .I(N__24115));
    LocalMux I__2614 (
            .O(N__24115),
            .I(N__24112));
    Odrv12 I__2613 (
            .O(N__24112),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ));
    InMux I__2612 (
            .O(N__24109),
            .I(N__24103));
    InMux I__2611 (
            .O(N__24108),
            .I(N__24103));
    LocalMux I__2610 (
            .O(N__24103),
            .I(N__24100));
    Odrv4 I__2609 (
            .O(N__24100),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ));
    InMux I__2608 (
            .O(N__24097),
            .I(N__24091));
    InMux I__2607 (
            .O(N__24096),
            .I(N__24091));
    LocalMux I__2606 (
            .O(N__24091),
            .I(N__24088));
    Odrv12 I__2605 (
            .O(N__24088),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ));
    InMux I__2604 (
            .O(N__24085),
            .I(N__24079));
    InMux I__2603 (
            .O(N__24084),
            .I(N__24079));
    LocalMux I__2602 (
            .O(N__24079),
            .I(N__24076));
    Odrv4 I__2601 (
            .O(N__24076),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ));
    InMux I__2600 (
            .O(N__24073),
            .I(bfn_7_7_0_));
    InMux I__2599 (
            .O(N__24070),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ));
    InMux I__2598 (
            .O(N__24067),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ));
    InMux I__2597 (
            .O(N__24064),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ));
    InMux I__2596 (
            .O(N__24061),
            .I(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ));
    InMux I__2595 (
            .O(N__24058),
            .I(N__24052));
    InMux I__2594 (
            .O(N__24057),
            .I(N__24052));
    LocalMux I__2593 (
            .O(N__24052),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ));
    InMux I__2592 (
            .O(N__24049),
            .I(N__24043));
    InMux I__2591 (
            .O(N__24048),
            .I(N__24043));
    LocalMux I__2590 (
            .O(N__24043),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ));
    CascadeMux I__2589 (
            .O(N__24040),
            .I(N__24036));
    CascadeMux I__2588 (
            .O(N__24039),
            .I(N__24033));
    InMux I__2587 (
            .O(N__24036),
            .I(N__24028));
    InMux I__2586 (
            .O(N__24033),
            .I(N__24028));
    LocalMux I__2585 (
            .O(N__24028),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ));
    InMux I__2584 (
            .O(N__24025),
            .I(N__24019));
    InMux I__2583 (
            .O(N__24024),
            .I(N__24019));
    LocalMux I__2582 (
            .O(N__24019),
            .I(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ));
    InMux I__2581 (
            .O(N__24016),
            .I(N__24010));
    InMux I__2580 (
            .O(N__24015),
            .I(N__24010));
    LocalMux I__2579 (
            .O(N__24010),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ));
    InMux I__2578 (
            .O(N__24007),
            .I(N__24001));
    InMux I__2577 (
            .O(N__24006),
            .I(N__24001));
    LocalMux I__2576 (
            .O(N__24001),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ));
    CascadeMux I__2575 (
            .O(N__23998),
            .I(N__23994));
    CascadeMux I__2574 (
            .O(N__23997),
            .I(N__23991));
    InMux I__2573 (
            .O(N__23994),
            .I(N__23986));
    InMux I__2572 (
            .O(N__23991),
            .I(N__23986));
    LocalMux I__2571 (
            .O(N__23986),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ));
    InMux I__2570 (
            .O(N__23983),
            .I(N__23977));
    InMux I__2569 (
            .O(N__23982),
            .I(N__23977));
    LocalMux I__2568 (
            .O(N__23977),
            .I(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ));
    InMux I__2567 (
            .O(N__23974),
            .I(N__23969));
    InMux I__2566 (
            .O(N__23973),
            .I(N__23966));
    InMux I__2565 (
            .O(N__23972),
            .I(N__23963));
    LocalMux I__2564 (
            .O(N__23969),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2563 (
            .O(N__23966),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    LocalMux I__2562 (
            .O(N__23963),
            .I(\pwm_generator_inst.counterZ0Z_4 ));
    InMux I__2561 (
            .O(N__23956),
            .I(\pwm_generator_inst.counter_cry_3 ));
    InMux I__2560 (
            .O(N__23953),
            .I(N__23948));
    InMux I__2559 (
            .O(N__23952),
            .I(N__23945));
    InMux I__2558 (
            .O(N__23951),
            .I(N__23942));
    LocalMux I__2557 (
            .O(N__23948),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2556 (
            .O(N__23945),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    LocalMux I__2555 (
            .O(N__23942),
            .I(\pwm_generator_inst.counterZ0Z_5 ));
    InMux I__2554 (
            .O(N__23935),
            .I(\pwm_generator_inst.counter_cry_4 ));
    InMux I__2553 (
            .O(N__23932),
            .I(N__23927));
    InMux I__2552 (
            .O(N__23931),
            .I(N__23924));
    InMux I__2551 (
            .O(N__23930),
            .I(N__23921));
    LocalMux I__2550 (
            .O(N__23927),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2549 (
            .O(N__23924),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    LocalMux I__2548 (
            .O(N__23921),
            .I(\pwm_generator_inst.counterZ0Z_6 ));
    InMux I__2547 (
            .O(N__23914),
            .I(\pwm_generator_inst.counter_cry_5 ));
    InMux I__2546 (
            .O(N__23911),
            .I(N__23906));
    InMux I__2545 (
            .O(N__23910),
            .I(N__23903));
    InMux I__2544 (
            .O(N__23909),
            .I(N__23900));
    LocalMux I__2543 (
            .O(N__23906),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2542 (
            .O(N__23903),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    LocalMux I__2541 (
            .O(N__23900),
            .I(\pwm_generator_inst.counterZ0Z_7 ));
    InMux I__2540 (
            .O(N__23893),
            .I(\pwm_generator_inst.counter_cry_6 ));
    InMux I__2539 (
            .O(N__23890),
            .I(N__23885));
    InMux I__2538 (
            .O(N__23889),
            .I(N__23882));
    InMux I__2537 (
            .O(N__23888),
            .I(N__23879));
    LocalMux I__2536 (
            .O(N__23885),
            .I(N__23876));
    LocalMux I__2535 (
            .O(N__23882),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    LocalMux I__2534 (
            .O(N__23879),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    Odrv4 I__2533 (
            .O(N__23876),
            .I(\pwm_generator_inst.counterZ0Z_8 ));
    InMux I__2532 (
            .O(N__23869),
            .I(bfn_4_19_0_));
    InMux I__2531 (
            .O(N__23866),
            .I(N__23852));
    InMux I__2530 (
            .O(N__23865),
            .I(N__23852));
    InMux I__2529 (
            .O(N__23864),
            .I(N__23843));
    InMux I__2528 (
            .O(N__23863),
            .I(N__23843));
    InMux I__2527 (
            .O(N__23862),
            .I(N__23843));
    InMux I__2526 (
            .O(N__23861),
            .I(N__23843));
    InMux I__2525 (
            .O(N__23860),
            .I(N__23834));
    InMux I__2524 (
            .O(N__23859),
            .I(N__23834));
    InMux I__2523 (
            .O(N__23858),
            .I(N__23834));
    InMux I__2522 (
            .O(N__23857),
            .I(N__23834));
    LocalMux I__2521 (
            .O(N__23852),
            .I(N__23831));
    LocalMux I__2520 (
            .O(N__23843),
            .I(\pwm_generator_inst.un1_counter_0 ));
    LocalMux I__2519 (
            .O(N__23834),
            .I(\pwm_generator_inst.un1_counter_0 ));
    Odrv4 I__2518 (
            .O(N__23831),
            .I(\pwm_generator_inst.un1_counter_0 ));
    InMux I__2517 (
            .O(N__23824),
            .I(\pwm_generator_inst.counter_cry_8 ));
    InMux I__2516 (
            .O(N__23821),
            .I(N__23816));
    InMux I__2515 (
            .O(N__23820),
            .I(N__23813));
    InMux I__2514 (
            .O(N__23819),
            .I(N__23810));
    LocalMux I__2513 (
            .O(N__23816),
            .I(N__23807));
    LocalMux I__2512 (
            .O(N__23813),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    LocalMux I__2511 (
            .O(N__23810),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    Odrv4 I__2510 (
            .O(N__23807),
            .I(\pwm_generator_inst.counterZ0Z_9 ));
    InMux I__2509 (
            .O(N__23800),
            .I(\pwm_generator_inst.un14_counter_cry_9 ));
    IoInMux I__2508 (
            .O(N__23797),
            .I(N__23794));
    LocalMux I__2507 (
            .O(N__23794),
            .I(N__23791));
    Span4Mux_s3_v I__2506 (
            .O(N__23791),
            .I(N__23788));
    Sp12to4 I__2505 (
            .O(N__23788),
            .I(N__23785));
    Span12Mux_s10_h I__2504 (
            .O(N__23785),
            .I(N__23782));
    Span12Mux_h I__2503 (
            .O(N__23782),
            .I(N__23779));
    Span12Mux_v I__2502 (
            .O(N__23779),
            .I(N__23776));
    Odrv12 I__2501 (
            .O(N__23776),
            .I(pwm_output_c));
    CascadeMux I__2500 (
            .O(N__23773),
            .I(\pwm_generator_inst.un1_counterlto2_0_cascade_ ));
    InMux I__2499 (
            .O(N__23770),
            .I(N__23767));
    LocalMux I__2498 (
            .O(N__23767),
            .I(\pwm_generator_inst.un1_counterlto9_2 ));
    CascadeMux I__2497 (
            .O(N__23764),
            .I(\pwm_generator_inst.un1_counterlt9_cascade_ ));
    InMux I__2496 (
            .O(N__23761),
            .I(N__23756));
    InMux I__2495 (
            .O(N__23760),
            .I(N__23753));
    InMux I__2494 (
            .O(N__23759),
            .I(N__23750));
    LocalMux I__2493 (
            .O(N__23756),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2492 (
            .O(N__23753),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    LocalMux I__2491 (
            .O(N__23750),
            .I(\pwm_generator_inst.counterZ0Z_0 ));
    InMux I__2490 (
            .O(N__23743),
            .I(bfn_4_18_0_));
    InMux I__2489 (
            .O(N__23740),
            .I(N__23735));
    InMux I__2488 (
            .O(N__23739),
            .I(N__23732));
    InMux I__2487 (
            .O(N__23738),
            .I(N__23729));
    LocalMux I__2486 (
            .O(N__23735),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2485 (
            .O(N__23732),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    LocalMux I__2484 (
            .O(N__23729),
            .I(\pwm_generator_inst.counterZ0Z_1 ));
    InMux I__2483 (
            .O(N__23722),
            .I(\pwm_generator_inst.counter_cry_0 ));
    InMux I__2482 (
            .O(N__23719),
            .I(N__23714));
    InMux I__2481 (
            .O(N__23718),
            .I(N__23711));
    InMux I__2480 (
            .O(N__23717),
            .I(N__23708));
    LocalMux I__2479 (
            .O(N__23714),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2478 (
            .O(N__23711),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    LocalMux I__2477 (
            .O(N__23708),
            .I(\pwm_generator_inst.counterZ0Z_2 ));
    InMux I__2476 (
            .O(N__23701),
            .I(\pwm_generator_inst.counter_cry_1 ));
    InMux I__2475 (
            .O(N__23698),
            .I(N__23693));
    InMux I__2474 (
            .O(N__23697),
            .I(N__23690));
    InMux I__2473 (
            .O(N__23696),
            .I(N__23687));
    LocalMux I__2472 (
            .O(N__23693),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2471 (
            .O(N__23690),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    LocalMux I__2470 (
            .O(N__23687),
            .I(\pwm_generator_inst.counterZ0Z_3 ));
    InMux I__2469 (
            .O(N__23680),
            .I(\pwm_generator_inst.counter_cry_2 ));
    CascadeMux I__2468 (
            .O(N__23677),
            .I(N__23674));
    InMux I__2467 (
            .O(N__23674),
            .I(N__23671));
    LocalMux I__2466 (
            .O(N__23671),
            .I(N__23668));
    Span4Mux_v I__2465 (
            .O(N__23668),
            .I(N__23665));
    Odrv4 I__2464 (
            .O(N__23665),
            .I(\pwm_generator_inst.N_181_i ));
    InMux I__2463 (
            .O(N__23662),
            .I(N__23659));
    LocalMux I__2462 (
            .O(N__23659),
            .I(\pwm_generator_inst.counter_i_2 ));
    CascadeMux I__2461 (
            .O(N__23656),
            .I(N__23653));
    InMux I__2460 (
            .O(N__23653),
            .I(N__23650));
    LocalMux I__2459 (
            .O(N__23650),
            .I(N__23647));
    Span12Mux_h I__2458 (
            .O(N__23647),
            .I(N__23644));
    Odrv12 I__2457 (
            .O(N__23644),
            .I(\pwm_generator_inst.N_182_i ));
    InMux I__2456 (
            .O(N__23641),
            .I(N__23638));
    LocalMux I__2455 (
            .O(N__23638),
            .I(\pwm_generator_inst.counter_i_3 ));
    CascadeMux I__2454 (
            .O(N__23635),
            .I(N__23632));
    InMux I__2453 (
            .O(N__23632),
            .I(N__23629));
    LocalMux I__2452 (
            .O(N__23629),
            .I(N__23626));
    Span4Mux_v I__2451 (
            .O(N__23626),
            .I(N__23623));
    Odrv4 I__2450 (
            .O(N__23623),
            .I(\pwm_generator_inst.N_183_i ));
    InMux I__2449 (
            .O(N__23620),
            .I(N__23617));
    LocalMux I__2448 (
            .O(N__23617),
            .I(\pwm_generator_inst.counter_i_4 ));
    InMux I__2447 (
            .O(N__23614),
            .I(N__23611));
    LocalMux I__2446 (
            .O(N__23611),
            .I(\pwm_generator_inst.N_184_i ));
    CascadeMux I__2445 (
            .O(N__23608),
            .I(N__23605));
    InMux I__2444 (
            .O(N__23605),
            .I(N__23602));
    LocalMux I__2443 (
            .O(N__23602),
            .I(\pwm_generator_inst.counter_i_5 ));
    CascadeMux I__2442 (
            .O(N__23599),
            .I(N__23596));
    InMux I__2441 (
            .O(N__23596),
            .I(N__23593));
    LocalMux I__2440 (
            .O(N__23593),
            .I(N__23590));
    Span4Mux_v I__2439 (
            .O(N__23590),
            .I(N__23587));
    Odrv4 I__2438 (
            .O(N__23587),
            .I(\pwm_generator_inst.N_185_i ));
    InMux I__2437 (
            .O(N__23584),
            .I(N__23581));
    LocalMux I__2436 (
            .O(N__23581),
            .I(\pwm_generator_inst.counter_i_6 ));
    CascadeMux I__2435 (
            .O(N__23578),
            .I(N__23575));
    InMux I__2434 (
            .O(N__23575),
            .I(N__23572));
    LocalMux I__2433 (
            .O(N__23572),
            .I(N__23569));
    Odrv4 I__2432 (
            .O(N__23569),
            .I(\pwm_generator_inst.N_186_i ));
    InMux I__2431 (
            .O(N__23566),
            .I(N__23563));
    LocalMux I__2430 (
            .O(N__23563),
            .I(\pwm_generator_inst.counter_i_7 ));
    CascadeMux I__2429 (
            .O(N__23560),
            .I(N__23557));
    InMux I__2428 (
            .O(N__23557),
            .I(N__23554));
    LocalMux I__2427 (
            .O(N__23554),
            .I(\pwm_generator_inst.N_187_i ));
    InMux I__2426 (
            .O(N__23551),
            .I(N__23548));
    LocalMux I__2425 (
            .O(N__23548),
            .I(\pwm_generator_inst.counter_i_8 ));
    CascadeMux I__2424 (
            .O(N__23545),
            .I(N__23542));
    InMux I__2423 (
            .O(N__23542),
            .I(N__23539));
    LocalMux I__2422 (
            .O(N__23539),
            .I(N__23536));
    Span4Mux_h I__2421 (
            .O(N__23536),
            .I(N__23533));
    Odrv4 I__2420 (
            .O(N__23533),
            .I(\pwm_generator_inst.N_188_i ));
    InMux I__2419 (
            .O(N__23530),
            .I(N__23527));
    LocalMux I__2418 (
            .O(N__23527),
            .I(\pwm_generator_inst.counter_i_9 ));
    CascadeMux I__2417 (
            .O(N__23524),
            .I(N__23520));
    InMux I__2416 (
            .O(N__23523),
            .I(N__23517));
    InMux I__2415 (
            .O(N__23520),
            .I(N__23514));
    LocalMux I__2414 (
            .O(N__23517),
            .I(\pwm_generator_inst.un18_threshold1_24 ));
    LocalMux I__2413 (
            .O(N__23514),
            .I(\pwm_generator_inst.un18_threshold1_24 ));
    InMux I__2412 (
            .O(N__23509),
            .I(N__23506));
    LocalMux I__2411 (
            .O(N__23506),
            .I(\pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO ));
    InMux I__2410 (
            .O(N__23503),
            .I(\pwm_generator_inst.un22_threshold_1_cry_6 ));
    InMux I__2409 (
            .O(N__23500),
            .I(bfn_2_18_0_));
    InMux I__2408 (
            .O(N__23497),
            .I(\pwm_generator_inst.un22_threshold_1_cry_8 ));
    CascadeMux I__2407 (
            .O(N__23494),
            .I(N__23491));
    InMux I__2406 (
            .O(N__23491),
            .I(N__23488));
    LocalMux I__2405 (
            .O(N__23488),
            .I(\pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO ));
    InMux I__2404 (
            .O(N__23485),
            .I(N__23482));
    LocalMux I__2403 (
            .O(N__23482),
            .I(N__23478));
    InMux I__2402 (
            .O(N__23481),
            .I(N__23475));
    Odrv4 I__2401 (
            .O(N__23478),
            .I(\pwm_generator_inst.un22_threshold_1 ));
    LocalMux I__2400 (
            .O(N__23475),
            .I(\pwm_generator_inst.un22_threshold_1 ));
    InMux I__2399 (
            .O(N__23470),
            .I(N__23466));
    InMux I__2398 (
            .O(N__23469),
            .I(N__23463));
    LocalMux I__2397 (
            .O(N__23466),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ));
    LocalMux I__2396 (
            .O(N__23463),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ));
    InMux I__2395 (
            .O(N__23458),
            .I(N__23454));
    InMux I__2394 (
            .O(N__23457),
            .I(N__23451));
    LocalMux I__2393 (
            .O(N__23454),
            .I(N__23448));
    LocalMux I__2392 (
            .O(N__23451),
            .I(N__23445));
    Odrv4 I__2391 (
            .O(N__23448),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ));
    Odrv4 I__2390 (
            .O(N__23445),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ));
    CascadeMux I__2389 (
            .O(N__23440),
            .I(N__23436));
    CascadeMux I__2388 (
            .O(N__23439),
            .I(N__23433));
    InMux I__2387 (
            .O(N__23436),
            .I(N__23428));
    InMux I__2386 (
            .O(N__23433),
            .I(N__23428));
    LocalMux I__2385 (
            .O(N__23428),
            .I(\pwm_generator_inst.un18_threshold1_25 ));
    InMux I__2384 (
            .O(N__23425),
            .I(N__23422));
    LocalMux I__2383 (
            .O(N__23422),
            .I(\pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO ));
    InMux I__2382 (
            .O(N__23419),
            .I(N__23416));
    LocalMux I__2381 (
            .O(N__23416),
            .I(\pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO ));
    InMux I__2380 (
            .O(N__23413),
            .I(N__23409));
    CascadeMux I__2379 (
            .O(N__23412),
            .I(N__23406));
    LocalMux I__2378 (
            .O(N__23409),
            .I(N__23403));
    InMux I__2377 (
            .O(N__23406),
            .I(N__23400));
    Odrv4 I__2376 (
            .O(N__23403),
            .I(\pwm_generator_inst.un18_threshold1_18 ));
    LocalMux I__2375 (
            .O(N__23400),
            .I(\pwm_generator_inst.un18_threshold1_18 ));
    CascadeMux I__2374 (
            .O(N__23395),
            .I(N__23388));
    InMux I__2373 (
            .O(N__23394),
            .I(N__23380));
    InMux I__2372 (
            .O(N__23393),
            .I(N__23375));
    InMux I__2371 (
            .O(N__23392),
            .I(N__23375));
    InMux I__2370 (
            .O(N__23391),
            .I(N__23368));
    InMux I__2369 (
            .O(N__23388),
            .I(N__23368));
    InMux I__2368 (
            .O(N__23387),
            .I(N__23368));
    InMux I__2367 (
            .O(N__23386),
            .I(N__23359));
    InMux I__2366 (
            .O(N__23385),
            .I(N__23359));
    InMux I__2365 (
            .O(N__23384),
            .I(N__23359));
    InMux I__2364 (
            .O(N__23383),
            .I(N__23359));
    LocalMux I__2363 (
            .O(N__23380),
            .I(N__23350));
    LocalMux I__2362 (
            .O(N__23375),
            .I(N__23350));
    LocalMux I__2361 (
            .O(N__23368),
            .I(N__23350));
    LocalMux I__2360 (
            .O(N__23359),
            .I(N__23350));
    Span4Mux_v I__2359 (
            .O(N__23350),
            .I(N__23347));
    Odrv4 I__2358 (
            .O(N__23347),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ));
    InMux I__2357 (
            .O(N__23344),
            .I(N__23340));
    InMux I__2356 (
            .O(N__23343),
            .I(N__23337));
    LocalMux I__2355 (
            .O(N__23340),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ));
    LocalMux I__2354 (
            .O(N__23337),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ));
    CascadeMux I__2353 (
            .O(N__23332),
            .I(N__23329));
    InMux I__2352 (
            .O(N__23329),
            .I(N__23326));
    LocalMux I__2351 (
            .O(N__23326),
            .I(\pwm_generator_inst.N_179_i ));
    InMux I__2350 (
            .O(N__23323),
            .I(N__23320));
    LocalMux I__2349 (
            .O(N__23320),
            .I(\pwm_generator_inst.counter_i_0 ));
    CascadeMux I__2348 (
            .O(N__23317),
            .I(N__23314));
    InMux I__2347 (
            .O(N__23314),
            .I(N__23311));
    LocalMux I__2346 (
            .O(N__23311),
            .I(\pwm_generator_inst.N_180_i ));
    InMux I__2345 (
            .O(N__23308),
            .I(N__23305));
    LocalMux I__2344 (
            .O(N__23305),
            .I(\pwm_generator_inst.counter_i_1 ));
    CascadeMux I__2343 (
            .O(N__23302),
            .I(N__23299));
    InMux I__2342 (
            .O(N__23299),
            .I(N__23296));
    LocalMux I__2341 (
            .O(N__23296),
            .I(N__23292));
    InMux I__2340 (
            .O(N__23295),
            .I(N__23289));
    Span4Mux_h I__2339 (
            .O(N__23292),
            .I(N__23284));
    LocalMux I__2338 (
            .O(N__23289),
            .I(N__23284));
    Odrv4 I__2337 (
            .O(N__23284),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ));
    InMux I__2336 (
            .O(N__23281),
            .I(\pwm_generator_inst.un22_threshold_1_cry_0 ));
    InMux I__2335 (
            .O(N__23278),
            .I(N__23274));
    InMux I__2334 (
            .O(N__23277),
            .I(N__23271));
    LocalMux I__2333 (
            .O(N__23274),
            .I(\pwm_generator_inst.un18_threshold1_19 ));
    LocalMux I__2332 (
            .O(N__23271),
            .I(\pwm_generator_inst.un18_threshold1_19 ));
    InMux I__2331 (
            .O(N__23266),
            .I(N__23263));
    LocalMux I__2330 (
            .O(N__23263),
            .I(N__23260));
    Odrv4 I__2329 (
            .O(N__23260),
            .I(\pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO ));
    InMux I__2328 (
            .O(N__23257),
            .I(\pwm_generator_inst.un22_threshold_1_cry_1 ));
    CascadeMux I__2327 (
            .O(N__23254),
            .I(N__23250));
    InMux I__2326 (
            .O(N__23253),
            .I(N__23247));
    InMux I__2325 (
            .O(N__23250),
            .I(N__23244));
    LocalMux I__2324 (
            .O(N__23247),
            .I(\pwm_generator_inst.un18_threshold1_20 ));
    LocalMux I__2323 (
            .O(N__23244),
            .I(\pwm_generator_inst.un18_threshold1_20 ));
    InMux I__2322 (
            .O(N__23239),
            .I(N__23236));
    LocalMux I__2321 (
            .O(N__23236),
            .I(N__23233));
    Odrv4 I__2320 (
            .O(N__23233),
            .I(\pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO ));
    InMux I__2319 (
            .O(N__23230),
            .I(\pwm_generator_inst.un22_threshold_1_cry_2 ));
    InMux I__2318 (
            .O(N__23227),
            .I(N__23223));
    InMux I__2317 (
            .O(N__23226),
            .I(N__23220));
    LocalMux I__2316 (
            .O(N__23223),
            .I(\pwm_generator_inst.un18_threshold1_21 ));
    LocalMux I__2315 (
            .O(N__23220),
            .I(\pwm_generator_inst.un18_threshold1_21 ));
    InMux I__2314 (
            .O(N__23215),
            .I(N__23212));
    LocalMux I__2313 (
            .O(N__23212),
            .I(N__23209));
    Odrv4 I__2312 (
            .O(N__23209),
            .I(\pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO ));
    InMux I__2311 (
            .O(N__23206),
            .I(\pwm_generator_inst.un22_threshold_1_cry_3 ));
    CascadeMux I__2310 (
            .O(N__23203),
            .I(N__23199));
    InMux I__2309 (
            .O(N__23202),
            .I(N__23196));
    InMux I__2308 (
            .O(N__23199),
            .I(N__23193));
    LocalMux I__2307 (
            .O(N__23196),
            .I(\pwm_generator_inst.un18_threshold1_22 ));
    LocalMux I__2306 (
            .O(N__23193),
            .I(\pwm_generator_inst.un18_threshold1_22 ));
    InMux I__2305 (
            .O(N__23188),
            .I(N__23185));
    LocalMux I__2304 (
            .O(N__23185),
            .I(\pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO ));
    InMux I__2303 (
            .O(N__23182),
            .I(\pwm_generator_inst.un22_threshold_1_cry_4 ));
    InMux I__2302 (
            .O(N__23179),
            .I(N__23175));
    InMux I__2301 (
            .O(N__23178),
            .I(N__23172));
    LocalMux I__2300 (
            .O(N__23175),
            .I(\pwm_generator_inst.un18_threshold1_23 ));
    LocalMux I__2299 (
            .O(N__23172),
            .I(\pwm_generator_inst.un18_threshold1_23 ));
    CascadeMux I__2298 (
            .O(N__23167),
            .I(N__23164));
    InMux I__2297 (
            .O(N__23164),
            .I(N__23161));
    LocalMux I__2296 (
            .O(N__23161),
            .I(N__23158));
    Odrv4 I__2295 (
            .O(N__23158),
            .I(\pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO ));
    InMux I__2294 (
            .O(N__23155),
            .I(\pwm_generator_inst.un22_threshold_1_cry_5 ));
    InMux I__2293 (
            .O(N__23152),
            .I(N__23149));
    LocalMux I__2292 (
            .O(N__23149),
            .I(N__23146));
    Odrv4 I__2291 (
            .O(N__23146),
            .I(\pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7 ));
    InMux I__2290 (
            .O(N__23143),
            .I(bfn_1_25_0_));
    InMux I__2289 (
            .O(N__23140),
            .I(N__23137));
    LocalMux I__2288 (
            .O(N__23137),
            .I(\pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7 ));
    InMux I__2287 (
            .O(N__23134),
            .I(\pwm_generator_inst.un3_threshold_cry_16 ));
    InMux I__2286 (
            .O(N__23131),
            .I(N__23128));
    LocalMux I__2285 (
            .O(N__23128),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0 ));
    InMux I__2284 (
            .O(N__23125),
            .I(\pwm_generator_inst.un3_threshold_cry_17 ));
    InMux I__2283 (
            .O(N__23122),
            .I(N__23118));
    InMux I__2282 (
            .O(N__23121),
            .I(N__23115));
    LocalMux I__2281 (
            .O(N__23118),
            .I(N__23110));
    LocalMux I__2280 (
            .O(N__23115),
            .I(N__23110));
    Odrv12 I__2279 (
            .O(N__23110),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ));
    InMux I__2278 (
            .O(N__23107),
            .I(\pwm_generator_inst.un3_threshold_cry_18 ));
    InMux I__2277 (
            .O(N__23104),
            .I(N__23101));
    LocalMux I__2276 (
            .O(N__23101),
            .I(N__23098));
    Span4Mux_v I__2275 (
            .O(N__23098),
            .I(N__23095));
    Span4Mux_v I__2274 (
            .O(N__23095),
            .I(N__23092));
    Odrv4 I__2273 (
            .O(N__23092),
            .I(\pwm_generator_inst.un2_threshold_2_12 ));
    InMux I__2272 (
            .O(N__23089),
            .I(\pwm_generator_inst.un3_threshold_cry_19 ));
    InMux I__2271 (
            .O(N__23086),
            .I(N__23083));
    LocalMux I__2270 (
            .O(N__23083),
            .I(N__23080));
    Odrv4 I__2269 (
            .O(N__23080),
            .I(\pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0 ));
    CascadeMux I__2268 (
            .O(N__23077),
            .I(N__23074));
    InMux I__2267 (
            .O(N__23074),
            .I(N__23071));
    LocalMux I__2266 (
            .O(N__23071),
            .I(N__23067));
    InMux I__2265 (
            .O(N__23070),
            .I(N__23064));
    Span4Mux_h I__2264 (
            .O(N__23067),
            .I(N__23059));
    LocalMux I__2263 (
            .O(N__23064),
            .I(N__23059));
    Odrv4 I__2262 (
            .O(N__23059),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0 ));
    CascadeMux I__2261 (
            .O(N__23056),
            .I(N__23053));
    InMux I__2260 (
            .O(N__23053),
            .I(N__23050));
    LocalMux I__2259 (
            .O(N__23050),
            .I(N__23047));
    Span4Mux_h I__2258 (
            .O(N__23047),
            .I(N__23043));
    InMux I__2257 (
            .O(N__23046),
            .I(N__23040));
    Odrv4 I__2256 (
            .O(N__23043),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ));
    LocalMux I__2255 (
            .O(N__23040),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ));
    CascadeMux I__2254 (
            .O(N__23035),
            .I(N__23032));
    InMux I__2253 (
            .O(N__23032),
            .I(N__23029));
    LocalMux I__2252 (
            .O(N__23029),
            .I(N__23025));
    InMux I__2251 (
            .O(N__23028),
            .I(N__23022));
    Span4Mux_v I__2250 (
            .O(N__23025),
            .I(N__23019));
    LocalMux I__2249 (
            .O(N__23022),
            .I(N__23016));
    Odrv4 I__2248 (
            .O(N__23019),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ));
    Odrv4 I__2247 (
            .O(N__23016),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ));
    InMux I__2246 (
            .O(N__23011),
            .I(N__23008));
    LocalMux I__2245 (
            .O(N__23008),
            .I(N__23004));
    InMux I__2244 (
            .O(N__23007),
            .I(N__23001));
    Span4Mux_v I__2243 (
            .O(N__23004),
            .I(N__22998));
    LocalMux I__2242 (
            .O(N__23001),
            .I(N__22995));
    Odrv4 I__2241 (
            .O(N__22998),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ));
    Odrv4 I__2240 (
            .O(N__22995),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ));
    InMux I__2239 (
            .O(N__22990),
            .I(N__22987));
    LocalMux I__2238 (
            .O(N__22987),
            .I(\pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0 ));
    InMux I__2237 (
            .O(N__22984),
            .I(bfn_1_24_0_));
    InMux I__2236 (
            .O(N__22981),
            .I(N__22978));
    LocalMux I__2235 (
            .O(N__22978),
            .I(\pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8 ));
    InMux I__2234 (
            .O(N__22975),
            .I(\pwm_generator_inst.un3_threshold_cry_8 ));
    InMux I__2233 (
            .O(N__22972),
            .I(N__22969));
    LocalMux I__2232 (
            .O(N__22969),
            .I(\pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8 ));
    InMux I__2231 (
            .O(N__22966),
            .I(\pwm_generator_inst.un3_threshold_cry_9 ));
    InMux I__2230 (
            .O(N__22963),
            .I(N__22960));
    LocalMux I__2229 (
            .O(N__22960),
            .I(\pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7 ));
    InMux I__2228 (
            .O(N__22957),
            .I(\pwm_generator_inst.un3_threshold_cry_10 ));
    InMux I__2227 (
            .O(N__22954),
            .I(N__22951));
    LocalMux I__2226 (
            .O(N__22951),
            .I(\pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7 ));
    InMux I__2225 (
            .O(N__22948),
            .I(\pwm_generator_inst.un3_threshold_cry_11 ));
    InMux I__2224 (
            .O(N__22945),
            .I(N__22942));
    LocalMux I__2223 (
            .O(N__22942),
            .I(\pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7 ));
    InMux I__2222 (
            .O(N__22939),
            .I(\pwm_generator_inst.un3_threshold_cry_12 ));
    InMux I__2221 (
            .O(N__22936),
            .I(N__22933));
    LocalMux I__2220 (
            .O(N__22933),
            .I(\pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7 ));
    InMux I__2219 (
            .O(N__22930),
            .I(\pwm_generator_inst.un3_threshold_cry_13 ));
    InMux I__2218 (
            .O(N__22927),
            .I(N__22924));
    LocalMux I__2217 (
            .O(N__22924),
            .I(\pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7 ));
    InMux I__2216 (
            .O(N__22921),
            .I(\pwm_generator_inst.un3_threshold_cry_14 ));
    CascadeMux I__2215 (
            .O(N__22918),
            .I(N__22915));
    InMux I__2214 (
            .O(N__22915),
            .I(N__22912));
    LocalMux I__2213 (
            .O(N__22912),
            .I(N__22909));
    Span12Mux_v I__2212 (
            .O(N__22909),
            .I(N__22906));
    Span12Mux_h I__2211 (
            .O(N__22906),
            .I(N__22903));
    Span12Mux_h I__2210 (
            .O(N__22903),
            .I(N__22900));
    Odrv12 I__2209 (
            .O(N__22900),
            .I(\pwm_generator_inst.O_0_8 ));
    InMux I__2208 (
            .O(N__22897),
            .I(N__22894));
    LocalMux I__2207 (
            .O(N__22894),
            .I(N__22891));
    Span12Mux_s1_h I__2206 (
            .O(N__22891),
            .I(N__22888));
    Odrv12 I__2205 (
            .O(N__22888),
            .I(\pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0 ));
    InMux I__2204 (
            .O(N__22885),
            .I(\pwm_generator_inst.un3_threshold_cry_0 ));
    CascadeMux I__2203 (
            .O(N__22882),
            .I(N__22879));
    InMux I__2202 (
            .O(N__22879),
            .I(N__22876));
    LocalMux I__2201 (
            .O(N__22876),
            .I(N__22873));
    Span12Mux_v I__2200 (
            .O(N__22873),
            .I(N__22870));
    Span12Mux_h I__2199 (
            .O(N__22870),
            .I(N__22867));
    Span12Mux_h I__2198 (
            .O(N__22867),
            .I(N__22864));
    Odrv12 I__2197 (
            .O(N__22864),
            .I(\pwm_generator_inst.O_0_9 ));
    InMux I__2196 (
            .O(N__22861),
            .I(N__22858));
    LocalMux I__2195 (
            .O(N__22858),
            .I(N__22855));
    Sp12to4 I__2194 (
            .O(N__22855),
            .I(N__22852));
    Odrv12 I__2193 (
            .O(N__22852),
            .I(\pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0 ));
    InMux I__2192 (
            .O(N__22849),
            .I(\pwm_generator_inst.un3_threshold_cry_1 ));
    InMux I__2191 (
            .O(N__22846),
            .I(N__22843));
    LocalMux I__2190 (
            .O(N__22843),
            .I(N__22840));
    Span4Mux_v I__2189 (
            .O(N__22840),
            .I(N__22837));
    Span4Mux_h I__2188 (
            .O(N__22837),
            .I(N__22834));
    Span4Mux_v I__2187 (
            .O(N__22834),
            .I(N__22831));
    Sp12to4 I__2186 (
            .O(N__22831),
            .I(N__22828));
    Span12Mux_h I__2185 (
            .O(N__22828),
            .I(N__22825));
    Odrv12 I__2184 (
            .O(N__22825),
            .I(\pwm_generator_inst.O_0_10 ));
    InMux I__2183 (
            .O(N__22822),
            .I(N__22819));
    LocalMux I__2182 (
            .O(N__22819),
            .I(N__22816));
    Span4Mux_v I__2181 (
            .O(N__22816),
            .I(N__22813));
    Span4Mux_v I__2180 (
            .O(N__22813),
            .I(N__22810));
    Odrv4 I__2179 (
            .O(N__22810),
            .I(\pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0 ));
    InMux I__2178 (
            .O(N__22807),
            .I(\pwm_generator_inst.un3_threshold_cry_2 ));
    InMux I__2177 (
            .O(N__22804),
            .I(N__22801));
    LocalMux I__2176 (
            .O(N__22801),
            .I(N__22798));
    Span12Mux_s11_v I__2175 (
            .O(N__22798),
            .I(N__22795));
    Span12Mux_h I__2174 (
            .O(N__22795),
            .I(N__22792));
    Span12Mux_h I__2173 (
            .O(N__22792),
            .I(N__22789));
    Odrv12 I__2172 (
            .O(N__22789),
            .I(\pwm_generator_inst.O_0_11 ));
    InMux I__2171 (
            .O(N__22786),
            .I(N__22783));
    LocalMux I__2170 (
            .O(N__22783),
            .I(N__22780));
    Odrv4 I__2169 (
            .O(N__22780),
            .I(\pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0 ));
    InMux I__2168 (
            .O(N__22777),
            .I(\pwm_generator_inst.un3_threshold_cry_3 ));
    InMux I__2167 (
            .O(N__22774),
            .I(N__22771));
    LocalMux I__2166 (
            .O(N__22771),
            .I(N__22768));
    Span4Mux_v I__2165 (
            .O(N__22768),
            .I(N__22765));
    Span4Mux_h I__2164 (
            .O(N__22765),
            .I(N__22762));
    Span4Mux_v I__2163 (
            .O(N__22762),
            .I(N__22759));
    Sp12to4 I__2162 (
            .O(N__22759),
            .I(N__22756));
    Span12Mux_h I__2161 (
            .O(N__22756),
            .I(N__22753));
    Odrv12 I__2160 (
            .O(N__22753),
            .I(\pwm_generator_inst.O_0_12 ));
    InMux I__2159 (
            .O(N__22750),
            .I(N__22747));
    LocalMux I__2158 (
            .O(N__22747),
            .I(N__22744));
    Span4Mux_s1_h I__2157 (
            .O(N__22744),
            .I(N__22741));
    Odrv4 I__2156 (
            .O(N__22741),
            .I(\pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0 ));
    InMux I__2155 (
            .O(N__22738),
            .I(\pwm_generator_inst.un3_threshold_cry_4 ));
    InMux I__2154 (
            .O(N__22735),
            .I(N__22732));
    LocalMux I__2153 (
            .O(N__22732),
            .I(N__22729));
    Span12Mux_s9_v I__2152 (
            .O(N__22729),
            .I(N__22726));
    Span12Mux_h I__2151 (
            .O(N__22726),
            .I(N__22723));
    Span12Mux_h I__2150 (
            .O(N__22723),
            .I(N__22720));
    Odrv12 I__2149 (
            .O(N__22720),
            .I(\pwm_generator_inst.O_0_13 ));
    InMux I__2148 (
            .O(N__22717),
            .I(N__22714));
    LocalMux I__2147 (
            .O(N__22714),
            .I(N__22711));
    Odrv4 I__2146 (
            .O(N__22711),
            .I(\pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0 ));
    InMux I__2145 (
            .O(N__22708),
            .I(\pwm_generator_inst.un3_threshold_cry_5 ));
    InMux I__2144 (
            .O(N__22705),
            .I(N__22702));
    LocalMux I__2143 (
            .O(N__22702),
            .I(N__22699));
    Span12Mux_s8_v I__2142 (
            .O(N__22699),
            .I(N__22696));
    Span12Mux_h I__2141 (
            .O(N__22696),
            .I(N__22693));
    Span12Mux_h I__2140 (
            .O(N__22693),
            .I(N__22690));
    Odrv12 I__2139 (
            .O(N__22690),
            .I(\pwm_generator_inst.O_0_14 ));
    InMux I__2138 (
            .O(N__22687),
            .I(N__22684));
    LocalMux I__2137 (
            .O(N__22684),
            .I(N__22681));
    Span4Mux_s1_h I__2136 (
            .O(N__22681),
            .I(N__22678));
    Odrv4 I__2135 (
            .O(N__22678),
            .I(\pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0 ));
    InMux I__2134 (
            .O(N__22675),
            .I(\pwm_generator_inst.un3_threshold_cry_6 ));
    CascadeMux I__2133 (
            .O(N__22672),
            .I(N__22669));
    InMux I__2132 (
            .O(N__22669),
            .I(N__22666));
    LocalMux I__2131 (
            .O(N__22666),
            .I(N__22663));
    Span4Mux_h I__2130 (
            .O(N__22663),
            .I(N__22660));
    Odrv4 I__2129 (
            .O(N__22660),
            .I(\pwm_generator_inst.un5_threshold_2_11 ));
    InMux I__2128 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__2127 (
            .O(N__22654),
            .I(N__22651));
    Odrv4 I__2126 (
            .O(N__22651),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0 ));
    InMux I__2125 (
            .O(N__22648),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_10 ));
    InMux I__2124 (
            .O(N__22645),
            .I(N__22642));
    LocalMux I__2123 (
            .O(N__22642),
            .I(N__22639));
    Span4Mux_h I__2122 (
            .O(N__22639),
            .I(N__22636));
    Odrv4 I__2121 (
            .O(N__22636),
            .I(\pwm_generator_inst.un5_threshold_2_12 ));
    CascadeMux I__2120 (
            .O(N__22633),
            .I(N__22630));
    InMux I__2119 (
            .O(N__22630),
            .I(N__22627));
    LocalMux I__2118 (
            .O(N__22627),
            .I(N__22624));
    Span4Mux_h I__2117 (
            .O(N__22624),
            .I(N__22621));
    Odrv4 I__2116 (
            .O(N__22621),
            .I(\pwm_generator_inst.un5_threshold_2_13 ));
    InMux I__2115 (
            .O(N__22618),
            .I(N__22615));
    LocalMux I__2114 (
            .O(N__22615),
            .I(N__22612));
    Span4Mux_v I__2113 (
            .O(N__22612),
            .I(N__22609));
    Odrv4 I__2112 (
            .O(N__22609),
            .I(\pwm_generator_inst.un5_threshold_2_14 ));
    InMux I__2111 (
            .O(N__22606),
            .I(bfn_1_21_0_));
    CascadeMux I__2110 (
            .O(N__22603),
            .I(N__22600));
    InMux I__2109 (
            .O(N__22600),
            .I(N__22597));
    LocalMux I__2108 (
            .O(N__22597),
            .I(N__22594));
    Odrv4 I__2107 (
            .O(N__22594),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0 ));
    CascadeMux I__2106 (
            .O(N__22591),
            .I(N__22584));
    CascadeMux I__2105 (
            .O(N__22590),
            .I(N__22580));
    InMux I__2104 (
            .O(N__22589),
            .I(N__22576));
    InMux I__2103 (
            .O(N__22588),
            .I(N__22573));
    InMux I__2102 (
            .O(N__22587),
            .I(N__22562));
    InMux I__2101 (
            .O(N__22584),
            .I(N__22562));
    InMux I__2100 (
            .O(N__22583),
            .I(N__22562));
    InMux I__2099 (
            .O(N__22580),
            .I(N__22562));
    InMux I__2098 (
            .O(N__22579),
            .I(N__22562));
    LocalMux I__2097 (
            .O(N__22576),
            .I(N__22557));
    LocalMux I__2096 (
            .O(N__22573),
            .I(N__22557));
    LocalMux I__2095 (
            .O(N__22562),
            .I(N__22552));
    Span4Mux_v I__2094 (
            .O(N__22557),
            .I(N__22552));
    Span4Mux_v I__2093 (
            .O(N__22552),
            .I(N__22549));
    Odrv4 I__2092 (
            .O(N__22549),
            .I(\pwm_generator_inst.un5_threshold_1_26 ));
    InMux I__2091 (
            .O(N__22546),
            .I(N__22543));
    LocalMux I__2090 (
            .O(N__22543),
            .I(N__22540));
    Odrv4 I__2089 (
            .O(N__22540),
            .I(\pwm_generator_inst.un5_threshold_2_1_16 ));
    CascadeMux I__2088 (
            .O(N__22537),
            .I(\pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_ ));
    InMux I__2087 (
            .O(N__22534),
            .I(N__22530));
    InMux I__2086 (
            .O(N__22533),
            .I(N__22527));
    LocalMux I__2085 (
            .O(N__22530),
            .I(N__22524));
    LocalMux I__2084 (
            .O(N__22527),
            .I(N__22521));
    Span4Mux_h I__2083 (
            .O(N__22524),
            .I(N__22518));
    Span4Mux_h I__2082 (
            .O(N__22521),
            .I(N__22515));
    Odrv4 I__2081 (
            .O(N__22518),
            .I(\pwm_generator_inst.un5_threshold_2_1_15 ));
    Odrv4 I__2080 (
            .O(N__22515),
            .I(\pwm_generator_inst.un5_threshold_2_1_15 ));
    InMux I__2079 (
            .O(N__22510),
            .I(N__22507));
    LocalMux I__2078 (
            .O(N__22507),
            .I(\pwm_generator_inst.un5_threshold_add_1_axb_16 ));
    InMux I__2077 (
            .O(N__22504),
            .I(N__22501));
    LocalMux I__2076 (
            .O(N__22501),
            .I(N__22498));
    Span4Mux_v I__2075 (
            .O(N__22498),
            .I(N__22495));
    Odrv4 I__2074 (
            .O(N__22495),
            .I(\pwm_generator_inst.un5_threshold_1_19 ));
    CascadeMux I__2073 (
            .O(N__22492),
            .I(N__22489));
    InMux I__2072 (
            .O(N__22489),
            .I(N__22486));
    LocalMux I__2071 (
            .O(N__22486),
            .I(N__22483));
    Span4Mux_h I__2070 (
            .O(N__22483),
            .I(N__22480));
    Odrv4 I__2069 (
            .O(N__22480),
            .I(\pwm_generator_inst.un5_threshold_2_4 ));
    InMux I__2068 (
            .O(N__22477),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_3 ));
    InMux I__2067 (
            .O(N__22474),
            .I(N__22471));
    LocalMux I__2066 (
            .O(N__22471),
            .I(N__22468));
    Span4Mux_v I__2065 (
            .O(N__22468),
            .I(N__22465));
    Odrv4 I__2064 (
            .O(N__22465),
            .I(\pwm_generator_inst.un5_threshold_1_20 ));
    CascadeMux I__2063 (
            .O(N__22462),
            .I(N__22459));
    InMux I__2062 (
            .O(N__22459),
            .I(N__22456));
    LocalMux I__2061 (
            .O(N__22456),
            .I(N__22453));
    Span4Mux_h I__2060 (
            .O(N__22453),
            .I(N__22450));
    Odrv4 I__2059 (
            .O(N__22450),
            .I(\pwm_generator_inst.un5_threshold_2_5 ));
    InMux I__2058 (
            .O(N__22447),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_4 ));
    InMux I__2057 (
            .O(N__22444),
            .I(N__22441));
    LocalMux I__2056 (
            .O(N__22441),
            .I(N__22438));
    Span4Mux_v I__2055 (
            .O(N__22438),
            .I(N__22435));
    Odrv4 I__2054 (
            .O(N__22435),
            .I(\pwm_generator_inst.un5_threshold_1_21 ));
    CascadeMux I__2053 (
            .O(N__22432),
            .I(N__22429));
    InMux I__2052 (
            .O(N__22429),
            .I(N__22426));
    LocalMux I__2051 (
            .O(N__22426),
            .I(N__22423));
    Span4Mux_v I__2050 (
            .O(N__22423),
            .I(N__22420));
    Odrv4 I__2049 (
            .O(N__22420),
            .I(\pwm_generator_inst.un5_threshold_2_6 ));
    InMux I__2048 (
            .O(N__22417),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_5 ));
    InMux I__2047 (
            .O(N__22414),
            .I(N__22411));
    LocalMux I__2046 (
            .O(N__22411),
            .I(N__22408));
    Span4Mux_v I__2045 (
            .O(N__22408),
            .I(N__22405));
    Odrv4 I__2044 (
            .O(N__22405),
            .I(\pwm_generator_inst.un5_threshold_1_22 ));
    CascadeMux I__2043 (
            .O(N__22402),
            .I(N__22399));
    InMux I__2042 (
            .O(N__22399),
            .I(N__22396));
    LocalMux I__2041 (
            .O(N__22396),
            .I(N__22393));
    Span4Mux_v I__2040 (
            .O(N__22393),
            .I(N__22390));
    Odrv4 I__2039 (
            .O(N__22390),
            .I(\pwm_generator_inst.un5_threshold_2_7 ));
    InMux I__2038 (
            .O(N__22387),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_6 ));
    InMux I__2037 (
            .O(N__22384),
            .I(N__22381));
    LocalMux I__2036 (
            .O(N__22381),
            .I(N__22378));
    Span4Mux_v I__2035 (
            .O(N__22378),
            .I(N__22375));
    Span4Mux_v I__2034 (
            .O(N__22375),
            .I(N__22372));
    Odrv4 I__2033 (
            .O(N__22372),
            .I(\pwm_generator_inst.un5_threshold_1_23 ));
    CascadeMux I__2032 (
            .O(N__22369),
            .I(N__22366));
    InMux I__2031 (
            .O(N__22366),
            .I(N__22363));
    LocalMux I__2030 (
            .O(N__22363),
            .I(N__22360));
    Span4Mux_h I__2029 (
            .O(N__22360),
            .I(N__22357));
    Odrv4 I__2028 (
            .O(N__22357),
            .I(\pwm_generator_inst.un5_threshold_2_8 ));
    InMux I__2027 (
            .O(N__22354),
            .I(bfn_1_20_0_));
    InMux I__2026 (
            .O(N__22351),
            .I(N__22348));
    LocalMux I__2025 (
            .O(N__22348),
            .I(N__22345));
    Span4Mux_v I__2024 (
            .O(N__22345),
            .I(N__22342));
    Span4Mux_v I__2023 (
            .O(N__22342),
            .I(N__22339));
    Odrv4 I__2022 (
            .O(N__22339),
            .I(\pwm_generator_inst.un5_threshold_1_24 ));
    CascadeMux I__2021 (
            .O(N__22336),
            .I(N__22333));
    InMux I__2020 (
            .O(N__22333),
            .I(N__22330));
    LocalMux I__2019 (
            .O(N__22330),
            .I(N__22327));
    Span4Mux_h I__2018 (
            .O(N__22327),
            .I(N__22324));
    Odrv4 I__2017 (
            .O(N__22324),
            .I(\pwm_generator_inst.un5_threshold_2_9 ));
    CascadeMux I__2016 (
            .O(N__22321),
            .I(N__22318));
    InMux I__2015 (
            .O(N__22318),
            .I(N__22314));
    InMux I__2014 (
            .O(N__22317),
            .I(N__22311));
    LocalMux I__2013 (
            .O(N__22314),
            .I(N__22308));
    LocalMux I__2012 (
            .O(N__22311),
            .I(N__22305));
    Odrv4 I__2011 (
            .O(N__22308),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ));
    Odrv4 I__2010 (
            .O(N__22305),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ));
    InMux I__2009 (
            .O(N__22300),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_8 ));
    InMux I__2008 (
            .O(N__22297),
            .I(N__22294));
    LocalMux I__2007 (
            .O(N__22294),
            .I(N__22291));
    Span4Mux_v I__2006 (
            .O(N__22291),
            .I(N__22288));
    Span4Mux_v I__2005 (
            .O(N__22288),
            .I(N__22285));
    Odrv4 I__2004 (
            .O(N__22285),
            .I(\pwm_generator_inst.un5_threshold_1_25 ));
    CascadeMux I__2003 (
            .O(N__22282),
            .I(N__22279));
    InMux I__2002 (
            .O(N__22279),
            .I(N__22276));
    LocalMux I__2001 (
            .O(N__22276),
            .I(N__22273));
    Span4Mux_h I__2000 (
            .O(N__22273),
            .I(N__22270));
    Odrv4 I__1999 (
            .O(N__22270),
            .I(\pwm_generator_inst.un5_threshold_2_10 ));
    InMux I__1998 (
            .O(N__22267),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_9 ));
    InMux I__1997 (
            .O(N__22264),
            .I(N__22261));
    LocalMux I__1996 (
            .O(N__22261),
            .I(N__22258));
    Odrv4 I__1995 (
            .O(N__22258),
            .I(\pwm_generator_inst.un18_threshold_1_axb_17 ));
    InMux I__1994 (
            .O(N__22255),
            .I(N__22252));
    LocalMux I__1993 (
            .O(N__22252),
            .I(\pwm_generator_inst.un18_threshold_1_axb_25 ));
    InMux I__1992 (
            .O(N__22249),
            .I(N__22246));
    LocalMux I__1991 (
            .O(N__22246),
            .I(N__22243));
    Odrv4 I__1990 (
            .O(N__22243),
            .I(\pwm_generator_inst.un18_threshold_1_axb_20 ));
    InMux I__1989 (
            .O(N__22240),
            .I(N__22237));
    LocalMux I__1988 (
            .O(N__22237),
            .I(\pwm_generator_inst.un18_threshold_1_axb_24 ));
    InMux I__1987 (
            .O(N__22234),
            .I(N__22231));
    LocalMux I__1986 (
            .O(N__22231),
            .I(N__22228));
    Odrv4 I__1985 (
            .O(N__22228),
            .I(\pwm_generator_inst.un18_threshold_1_axb_18 ));
    InMux I__1984 (
            .O(N__22225),
            .I(N__22222));
    LocalMux I__1983 (
            .O(N__22222),
            .I(N__22219));
    Span4Mux_h I__1982 (
            .O(N__22219),
            .I(N__22216));
    Odrv4 I__1981 (
            .O(N__22216),
            .I(\pwm_generator_inst.un5_threshold_2_0 ));
    CascadeMux I__1980 (
            .O(N__22213),
            .I(N__22210));
    InMux I__1979 (
            .O(N__22210),
            .I(N__22207));
    LocalMux I__1978 (
            .O(N__22207),
            .I(N__22204));
    Span12Mux_v I__1977 (
            .O(N__22204),
            .I(N__22201));
    Odrv12 I__1976 (
            .O(N__22201),
            .I(\pwm_generator_inst.un5_threshold_1_15 ));
    InMux I__1975 (
            .O(N__22198),
            .I(N__22195));
    LocalMux I__1974 (
            .O(N__22195),
            .I(N__22192));
    Odrv12 I__1973 (
            .O(N__22192),
            .I(\pwm_generator_inst.un18_threshold_1_axb_15 ));
    InMux I__1972 (
            .O(N__22189),
            .I(N__22186));
    LocalMux I__1971 (
            .O(N__22186),
            .I(N__22183));
    Span4Mux_h I__1970 (
            .O(N__22183),
            .I(N__22180));
    Odrv4 I__1969 (
            .O(N__22180),
            .I(\pwm_generator_inst.un5_threshold_2_1 ));
    CascadeMux I__1968 (
            .O(N__22177),
            .I(N__22174));
    InMux I__1967 (
            .O(N__22174),
            .I(N__22171));
    LocalMux I__1966 (
            .O(N__22171),
            .I(N__22168));
    Span4Mux_v I__1965 (
            .O(N__22168),
            .I(N__22165));
    Span4Mux_v I__1964 (
            .O(N__22165),
            .I(N__22162));
    Odrv4 I__1963 (
            .O(N__22162),
            .I(\pwm_generator_inst.un5_threshold_1_16 ));
    InMux I__1962 (
            .O(N__22159),
            .I(N__22156));
    LocalMux I__1961 (
            .O(N__22156),
            .I(N__22153));
    Odrv12 I__1960 (
            .O(N__22153),
            .I(\pwm_generator_inst.un18_threshold_1_axb_16 ));
    InMux I__1959 (
            .O(N__22150),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_0 ));
    InMux I__1958 (
            .O(N__22147),
            .I(N__22144));
    LocalMux I__1957 (
            .O(N__22144),
            .I(N__22141));
    Span4Mux_h I__1956 (
            .O(N__22141),
            .I(N__22138));
    Odrv4 I__1955 (
            .O(N__22138),
            .I(\pwm_generator_inst.un5_threshold_2_2 ));
    CascadeMux I__1954 (
            .O(N__22135),
            .I(N__22132));
    InMux I__1953 (
            .O(N__22132),
            .I(N__22129));
    LocalMux I__1952 (
            .O(N__22129),
            .I(N__22126));
    Span4Mux_v I__1951 (
            .O(N__22126),
            .I(N__22123));
    Span4Mux_v I__1950 (
            .O(N__22123),
            .I(N__22120));
    Odrv4 I__1949 (
            .O(N__22120),
            .I(\pwm_generator_inst.un5_threshold_1_17 ));
    InMux I__1948 (
            .O(N__22117),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_1 ));
    InMux I__1947 (
            .O(N__22114),
            .I(N__22111));
    LocalMux I__1946 (
            .O(N__22111),
            .I(N__22108));
    Span4Mux_h I__1945 (
            .O(N__22108),
            .I(N__22105));
    Odrv4 I__1944 (
            .O(N__22105),
            .I(\pwm_generator_inst.un5_threshold_2_3 ));
    CascadeMux I__1943 (
            .O(N__22102),
            .I(N__22099));
    InMux I__1942 (
            .O(N__22099),
            .I(N__22096));
    LocalMux I__1941 (
            .O(N__22096),
            .I(N__22093));
    Span4Mux_v I__1940 (
            .O(N__22093),
            .I(N__22090));
    Odrv4 I__1939 (
            .O(N__22090),
            .I(\pwm_generator_inst.un5_threshold_1_18 ));
    InMux I__1938 (
            .O(N__22087),
            .I(\pwm_generator_inst.un5_threshold_add_1_cry_2 ));
    InMux I__1937 (
            .O(N__22084),
            .I(\pwm_generator_inst.un18_threshold_1_cry_22 ));
    InMux I__1936 (
            .O(N__22081),
            .I(bfn_1_17_0_));
    InMux I__1935 (
            .O(N__22078),
            .I(\pwm_generator_inst.un18_threshold_1_cry_24 ));
    InMux I__1934 (
            .O(N__22075),
            .I(\pwm_generator_inst.un18_threshold_1_cry_25 ));
    InMux I__1933 (
            .O(N__22072),
            .I(N__22069));
    LocalMux I__1932 (
            .O(N__22069),
            .I(\pwm_generator_inst.un18_threshold_1_axb_19 ));
    InMux I__1931 (
            .O(N__22066),
            .I(N__22063));
    LocalMux I__1930 (
            .O(N__22063),
            .I(\pwm_generator_inst.un18_threshold_1_axb_21 ));
    InMux I__1929 (
            .O(N__22060),
            .I(N__22057));
    LocalMux I__1928 (
            .O(N__22057),
            .I(\pwm_generator_inst.un18_threshold_1_axb_22 ));
    InMux I__1927 (
            .O(N__22054),
            .I(N__22051));
    LocalMux I__1926 (
            .O(N__22051),
            .I(\pwm_generator_inst.un18_threshold_1_axb_23 ));
    InMux I__1925 (
            .O(N__22048),
            .I(N__22045));
    LocalMux I__1924 (
            .O(N__22045),
            .I(N__22042));
    Span4Mux_v I__1923 (
            .O(N__22042),
            .I(N__22039));
    Odrv4 I__1922 (
            .O(N__22039),
            .I(\pwm_generator_inst.O_14 ));
    InMux I__1921 (
            .O(N__22036),
            .I(N__22033));
    LocalMux I__1920 (
            .O(N__22033),
            .I(\pwm_generator_inst.un18_threshold_1_axb_14 ));
    InMux I__1919 (
            .O(N__22030),
            .I(\pwm_generator_inst.un18_threshold_1_cry_16 ));
    InMux I__1918 (
            .O(N__22027),
            .I(\pwm_generator_inst.un18_threshold_1_cry_17 ));
    InMux I__1917 (
            .O(N__22024),
            .I(\pwm_generator_inst.un18_threshold_1_cry_18 ));
    InMux I__1916 (
            .O(N__22021),
            .I(\pwm_generator_inst.un18_threshold_1_cry_19 ));
    InMux I__1915 (
            .O(N__22018),
            .I(\pwm_generator_inst.un18_threshold_1_cry_20 ));
    InMux I__1914 (
            .O(N__22015),
            .I(\pwm_generator_inst.un18_threshold_1_cry_21 ));
    InMux I__1913 (
            .O(N__22012),
            .I(N__22009));
    LocalMux I__1912 (
            .O(N__22009),
            .I(N__22006));
    Span4Mux_v I__1911 (
            .O(N__22006),
            .I(N__22003));
    Odrv4 I__1910 (
            .O(N__22003),
            .I(\pwm_generator_inst.O_6 ));
    InMux I__1909 (
            .O(N__22000),
            .I(N__21997));
    LocalMux I__1908 (
            .O(N__21997),
            .I(\pwm_generator_inst.un18_threshold_1_axb_6 ));
    InMux I__1907 (
            .O(N__21994),
            .I(N__21991));
    LocalMux I__1906 (
            .O(N__21991),
            .I(N__21988));
    Span4Mux_v I__1905 (
            .O(N__21988),
            .I(N__21985));
    Odrv4 I__1904 (
            .O(N__21985),
            .I(\pwm_generator_inst.O_7 ));
    InMux I__1903 (
            .O(N__21982),
            .I(N__21979));
    LocalMux I__1902 (
            .O(N__21979),
            .I(\pwm_generator_inst.un18_threshold_1_axb_7 ));
    InMux I__1901 (
            .O(N__21976),
            .I(N__21973));
    LocalMux I__1900 (
            .O(N__21973),
            .I(N__21970));
    Span4Mux_v I__1899 (
            .O(N__21970),
            .I(N__21967));
    Odrv4 I__1898 (
            .O(N__21967),
            .I(\pwm_generator_inst.O_8 ));
    InMux I__1897 (
            .O(N__21964),
            .I(N__21961));
    LocalMux I__1896 (
            .O(N__21961),
            .I(\pwm_generator_inst.un18_threshold_1_axb_8 ));
    InMux I__1895 (
            .O(N__21958),
            .I(N__21955));
    LocalMux I__1894 (
            .O(N__21955),
            .I(N__21952));
    Span4Mux_v I__1893 (
            .O(N__21952),
            .I(N__21949));
    Odrv4 I__1892 (
            .O(N__21949),
            .I(\pwm_generator_inst.O_9 ));
    InMux I__1891 (
            .O(N__21946),
            .I(N__21943));
    LocalMux I__1890 (
            .O(N__21943),
            .I(\pwm_generator_inst.un18_threshold_1_axb_9 ));
    InMux I__1889 (
            .O(N__21940),
            .I(N__21937));
    LocalMux I__1888 (
            .O(N__21937),
            .I(N__21934));
    Span4Mux_v I__1887 (
            .O(N__21934),
            .I(N__21931));
    Odrv4 I__1886 (
            .O(N__21931),
            .I(\pwm_generator_inst.O_10 ));
    InMux I__1885 (
            .O(N__21928),
            .I(N__21925));
    LocalMux I__1884 (
            .O(N__21925),
            .I(\pwm_generator_inst.un18_threshold_1_axb_10 ));
    InMux I__1883 (
            .O(N__21922),
            .I(N__21919));
    LocalMux I__1882 (
            .O(N__21919),
            .I(N__21916));
    Span4Mux_v I__1881 (
            .O(N__21916),
            .I(N__21913));
    Odrv4 I__1880 (
            .O(N__21913),
            .I(\pwm_generator_inst.O_11 ));
    InMux I__1879 (
            .O(N__21910),
            .I(N__21907));
    LocalMux I__1878 (
            .O(N__21907),
            .I(\pwm_generator_inst.un18_threshold_1_axb_11 ));
    InMux I__1877 (
            .O(N__21904),
            .I(N__21901));
    LocalMux I__1876 (
            .O(N__21901),
            .I(N__21898));
    Span4Mux_v I__1875 (
            .O(N__21898),
            .I(N__21895));
    Odrv4 I__1874 (
            .O(N__21895),
            .I(\pwm_generator_inst.O_12 ));
    InMux I__1873 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__1872 (
            .O(N__21889),
            .I(\pwm_generator_inst.un18_threshold_1_axb_12 ));
    InMux I__1871 (
            .O(N__21886),
            .I(N__21883));
    LocalMux I__1870 (
            .O(N__21883),
            .I(N__21880));
    Span4Mux_v I__1869 (
            .O(N__21880),
            .I(N__21877));
    Odrv4 I__1868 (
            .O(N__21877),
            .I(\pwm_generator_inst.O_13 ));
    InMux I__1867 (
            .O(N__21874),
            .I(N__21871));
    LocalMux I__1866 (
            .O(N__21871),
            .I(\pwm_generator_inst.un18_threshold_1_axb_13 ));
    InMux I__1865 (
            .O(N__21868),
            .I(N__21865));
    LocalMux I__1864 (
            .O(N__21865),
            .I(N__21862));
    Span4Mux_v I__1863 (
            .O(N__21862),
            .I(N__21859));
    Odrv4 I__1862 (
            .O(N__21859),
            .I(\pwm_generator_inst.O_0 ));
    InMux I__1861 (
            .O(N__21856),
            .I(N__21853));
    LocalMux I__1860 (
            .O(N__21853),
            .I(\pwm_generator_inst.un18_threshold_1_axb_0 ));
    InMux I__1859 (
            .O(N__21850),
            .I(N__21847));
    LocalMux I__1858 (
            .O(N__21847),
            .I(N__21844));
    Span4Mux_v I__1857 (
            .O(N__21844),
            .I(N__21841));
    Odrv4 I__1856 (
            .O(N__21841),
            .I(\pwm_generator_inst.O_1 ));
    InMux I__1855 (
            .O(N__21838),
            .I(N__21835));
    LocalMux I__1854 (
            .O(N__21835),
            .I(\pwm_generator_inst.un18_threshold_1_axb_1 ));
    InMux I__1853 (
            .O(N__21832),
            .I(N__21829));
    LocalMux I__1852 (
            .O(N__21829),
            .I(N__21826));
    Span4Mux_v I__1851 (
            .O(N__21826),
            .I(N__21823));
    Odrv4 I__1850 (
            .O(N__21823),
            .I(\pwm_generator_inst.O_2 ));
    InMux I__1849 (
            .O(N__21820),
            .I(N__21817));
    LocalMux I__1848 (
            .O(N__21817),
            .I(\pwm_generator_inst.un18_threshold_1_axb_2 ));
    InMux I__1847 (
            .O(N__21814),
            .I(N__21811));
    LocalMux I__1846 (
            .O(N__21811),
            .I(N__21808));
    Span4Mux_v I__1845 (
            .O(N__21808),
            .I(N__21805));
    Odrv4 I__1844 (
            .O(N__21805),
            .I(\pwm_generator_inst.O_3 ));
    InMux I__1843 (
            .O(N__21802),
            .I(N__21799));
    LocalMux I__1842 (
            .O(N__21799),
            .I(\pwm_generator_inst.un18_threshold_1_axb_3 ));
    InMux I__1841 (
            .O(N__21796),
            .I(N__21793));
    LocalMux I__1840 (
            .O(N__21793),
            .I(N__21790));
    Span4Mux_v I__1839 (
            .O(N__21790),
            .I(N__21787));
    Odrv4 I__1838 (
            .O(N__21787),
            .I(\pwm_generator_inst.O_4 ));
    InMux I__1837 (
            .O(N__21784),
            .I(N__21781));
    LocalMux I__1836 (
            .O(N__21781),
            .I(\pwm_generator_inst.un18_threshold_1_axb_4 ));
    InMux I__1835 (
            .O(N__21778),
            .I(N__21775));
    LocalMux I__1834 (
            .O(N__21775),
            .I(N__21772));
    Span4Mux_v I__1833 (
            .O(N__21772),
            .I(N__21769));
    Odrv4 I__1832 (
            .O(N__21769),
            .I(\pwm_generator_inst.O_5 ));
    InMux I__1831 (
            .O(N__21766),
            .I(N__21763));
    LocalMux I__1830 (
            .O(N__21763),
            .I(\pwm_generator_inst.un18_threshold_1_axb_5 ));
    InMux I__1829 (
            .O(N__21760),
            .I(N__21757));
    LocalMux I__1828 (
            .O(N__21757),
            .I(N__21754));
    Span4Mux_v I__1827 (
            .O(N__21754),
            .I(N__21751));
    Sp12to4 I__1826 (
            .O(N__21751),
            .I(N__21748));
    Span12Mux_s8_h I__1825 (
            .O(N__21748),
            .I(N__21745));
    Span12Mux_h I__1824 (
            .O(N__21745),
            .I(N__21742));
    Odrv12 I__1823 (
            .O(N__21742),
            .I(\pwm_generator_inst.O_0_1 ));
    InMux I__1822 (
            .O(N__21739),
            .I(N__21736));
    LocalMux I__1821 (
            .O(N__21736),
            .I(N__21733));
    Span4Mux_v I__1820 (
            .O(N__21733),
            .I(N__21730));
    Sp12to4 I__1819 (
            .O(N__21730),
            .I(N__21727));
    Span12Mux_s9_h I__1818 (
            .O(N__21727),
            .I(N__21724));
    Span12Mux_h I__1817 (
            .O(N__21724),
            .I(N__21721));
    Odrv12 I__1816 (
            .O(N__21721),
            .I(\pwm_generator_inst.O_0_0 ));
    InMux I__1815 (
            .O(N__21718),
            .I(N__21715));
    LocalMux I__1814 (
            .O(N__21715),
            .I(N__21712));
    Span4Mux_h I__1813 (
            .O(N__21712),
            .I(N__21709));
    Sp12to4 I__1812 (
            .O(N__21709),
            .I(N__21706));
    Span12Mux_v I__1811 (
            .O(N__21706),
            .I(N__21703));
    Span12Mux_h I__1810 (
            .O(N__21703),
            .I(N__21700));
    Span12Mux_v I__1809 (
            .O(N__21700),
            .I(N__21697));
    Odrv12 I__1808 (
            .O(N__21697),
            .I(\pwm_generator_inst.O_0_5 ));
    InMux I__1807 (
            .O(N__21694),
            .I(N__21691));
    LocalMux I__1806 (
            .O(N__21691),
            .I(N__21688));
    Span4Mux_v I__1805 (
            .O(N__21688),
            .I(N__21685));
    Sp12to4 I__1804 (
            .O(N__21685),
            .I(N__21682));
    Span12Mux_s6_h I__1803 (
            .O(N__21682),
            .I(N__21679));
    Span12Mux_h I__1802 (
            .O(N__21679),
            .I(N__21676));
    Odrv12 I__1801 (
            .O(N__21676),
            .I(\pwm_generator_inst.O_0_3 ));
    InMux I__1800 (
            .O(N__21673),
            .I(N__21670));
    LocalMux I__1799 (
            .O(N__21670),
            .I(N__21667));
    Span4Mux_v I__1798 (
            .O(N__21667),
            .I(N__21664));
    Span4Mux_h I__1797 (
            .O(N__21664),
            .I(N__21661));
    Span4Mux_h I__1796 (
            .O(N__21661),
            .I(N__21658));
    Span4Mux_h I__1795 (
            .O(N__21658),
            .I(N__21655));
    Span4Mux_h I__1794 (
            .O(N__21655),
            .I(N__21652));
    Sp12to4 I__1793 (
            .O(N__21652),
            .I(N__21649));
    Odrv12 I__1792 (
            .O(N__21649),
            .I(\pwm_generator_inst.O_0_4 ));
    InMux I__1791 (
            .O(N__21646),
            .I(N__21643));
    LocalMux I__1790 (
            .O(N__21643),
            .I(N__21640));
    Span4Mux_v I__1789 (
            .O(N__21640),
            .I(N__21637));
    Sp12to4 I__1788 (
            .O(N__21637),
            .I(N__21634));
    Span12Mux_s7_h I__1787 (
            .O(N__21634),
            .I(N__21631));
    Span12Mux_h I__1786 (
            .O(N__21631),
            .I(N__21628));
    Odrv12 I__1785 (
            .O(N__21628),
            .I(\pwm_generator_inst.O_0_2 ));
    InMux I__1784 (
            .O(N__21625),
            .I(N__21622));
    LocalMux I__1783 (
            .O(N__21622),
            .I(N__21619));
    Span4Mux_v I__1782 (
            .O(N__21619),
            .I(N__21616));
    Sp12to4 I__1781 (
            .O(N__21616),
            .I(N__21613));
    Span12Mux_h I__1780 (
            .O(N__21613),
            .I(N__21610));
    Span12Mux_h I__1779 (
            .O(N__21610),
            .I(N__21607));
    Odrv12 I__1778 (
            .O(N__21607),
            .I(\pwm_generator_inst.O_0_6 ));
    IoInMux I__1777 (
            .O(N__21604),
            .I(N__21601));
    LocalMux I__1776 (
            .O(N__21601),
            .I(N__21598));
    Span4Mux_s3_v I__1775 (
            .O(N__21598),
            .I(N__21595));
    Span4Mux_h I__1774 (
            .O(N__21595),
            .I(N__21592));
    Sp12to4 I__1773 (
            .O(N__21592),
            .I(N__21589));
    Span12Mux_v I__1772 (
            .O(N__21589),
            .I(N__21586));
    Span12Mux_v I__1771 (
            .O(N__21586),
            .I(N__21583));
    Odrv12 I__1770 (
            .O(N__21583),
            .I(delay_tr_input_ibuf_gb_io_gb_input));
    IoInMux I__1769 (
            .O(N__21580),
            .I(N__21577));
    LocalMux I__1768 (
            .O(N__21577),
            .I(N__21574));
    IoSpan4Mux I__1767 (
            .O(N__21574),
            .I(N__21571));
    IoSpan4Mux I__1766 (
            .O(N__21571),
            .I(N__21568));
    Odrv4 I__1765 (
            .O(N__21568),
            .I(delay_hc_input_ibuf_gb_io_gb_input));
    defparam IN_MUX_bfv_1_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_23_0_));
    defparam IN_MUX_bfv_1_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_24_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_7 ),
            .carryinitout(bfn_1_24_0_));
    defparam IN_MUX_bfv_1_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_25_0_ (
            .carryinitin(\pwm_generator_inst.un3_threshold_cry_15 ),
            .carryinitout(bfn_1_25_0_));
    defparam IN_MUX_bfv_2_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_17_0_));
    defparam IN_MUX_bfv_2_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_18_0_ (
            .carryinitin(\pwm_generator_inst.un22_threshold_1_cry_7 ),
            .carryinitout(bfn_2_18_0_));
    defparam IN_MUX_bfv_18_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_17_0_));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_17_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_18_0_));
    defparam IN_MUX_bfv_17_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_19_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .carryinitout(bfn_17_19_0_));
    defparam IN_MUX_bfv_17_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_20_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .carryinitout(bfn_17_20_0_));
    defparam IN_MUX_bfv_17_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_21_0_ (
            .carryinitin(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .carryinitout(bfn_17_21_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_7 ),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_15 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_15_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_19_0_ (
            .carryinitin(\current_shift_inst.un10_control_input_cry_23 ),
            .carryinitout(bfn_15_19_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_12_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .carryinitout(bfn_12_21_0_));
    defparam IN_MUX_bfv_12_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .carryinitout(bfn_12_22_0_));
    defparam IN_MUX_bfv_12_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_23_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .carryinitout(bfn_12_23_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_1_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_19_0_));
    defparam IN_MUX_bfv_1_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_20_0_ (
            .carryinitin(\pwm_generator_inst.un5_threshold_add_1_cry_7 ),
            .carryinitout(bfn_1_20_0_));
    defparam IN_MUX_bfv_1_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_21_0_ (
            .carryinitin(\pwm_generator_inst.un5_threshold_add_1_cry_15 ),
            .carryinitout(bfn_1_21_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\pwm_generator_inst.un18_threshold_1_cry_7 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_1_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_16_0_ (
            .carryinitin(\pwm_generator_inst.un18_threshold_1_cry_15 ),
            .carryinitout(bfn_1_16_0_));
    defparam IN_MUX_bfv_1_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_17_0_ (
            .carryinitin(\pwm_generator_inst.un18_threshold_1_cry_23 ),
            .carryinitout(bfn_1_17_0_));
    defparam IN_MUX_bfv_3_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_17_0_));
    defparam IN_MUX_bfv_3_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_18_0_ (
            .carryinitin(\pwm_generator_inst.un14_counter_cry_7 ),
            .carryinitout(bfn_3_18_0_));
    defparam IN_MUX_bfv_4_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_18_0_));
    defparam IN_MUX_bfv_4_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_19_0_ (
            .carryinitin(\pwm_generator_inst.counter_cry_7 ),
            .carryinitout(bfn_4_19_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .carryinitout(bfn_7_18_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .carryinitout(bfn_7_19_0_));
    defparam IN_MUX_bfv_7_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.un6_running_cry_30 ),
            .carryinitout(bfn_7_20_0_));
    defparam IN_MUX_bfv_8_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_17_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_7 ),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_19_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_15 ),
            .carryinitout(bfn_8_19_0_));
    defparam IN_MUX_bfv_8_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_20_0_ (
            .carryinitin(\phase_controller_inst2.stoper_tr.counter_cry_23 ),
            .carryinitout(bfn_8_20_0_));
    defparam IN_MUX_bfv_11_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_5_0_));
    defparam IN_MUX_bfv_11_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_6_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .carryinitout(bfn_11_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.un6_running_cry_30 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_7 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_15 ),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\phase_controller_inst2.stoper_hc.counter_cry_23 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_10_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un6_running_cry_30 ),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_8_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_13_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_7 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_15 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\phase_controller_inst1.stoper_tr.counter_cry_23 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_14_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_5_0_));
    defparam IN_MUX_bfv_14_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_6_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .carryinitout(bfn_14_6_0_));
    defparam IN_MUX_bfv_14_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_7_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .carryinitout(bfn_14_7_0_));
    defparam IN_MUX_bfv_14_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un6_running_cry_30 ),
            .carryinitout(bfn_14_8_0_));
    defparam IN_MUX_bfv_16_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_8_0_));
    defparam IN_MUX_bfv_16_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ),
            .carryinitout(bfn_16_9_0_));
    defparam IN_MUX_bfv_16_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ),
            .carryinitout(bfn_16_10_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ),
            .carryinitout(bfn_15_9_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_7 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_15 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\phase_controller_inst1.stoper_hc.counter_cry_23 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .carryinitout(bfn_7_10_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_13_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_17_13_0_));
    defparam IN_MUX_bfv_18_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_7_0_));
    defparam IN_MUX_bfv_18_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_8_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .carryinitout(bfn_18_8_0_));
    defparam IN_MUX_bfv_18_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_9_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .carryinitout(bfn_18_9_0_));
    defparam IN_MUX_bfv_18_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_10_0_ (
            .carryinitin(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .carryinitout(bfn_18_10_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_14_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_20_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_7 ),
            .carryinitout(bfn_14_20_0_));
    defparam IN_MUX_bfv_14_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_21_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_15 ),
            .carryinitout(bfn_14_21_0_));
    defparam IN_MUX_bfv_14_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_22_0_ (
            .carryinitin(\current_shift_inst.control_input_cry_23 ),
            .carryinitout(bfn_14_22_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_16_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_13_0_));
    defparam IN_MUX_bfv_16_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_14_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_8 ),
            .carryinitout(bfn_16_14_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_16 ),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\current_shift_inst.un4_control_input_1_cry_24 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_7 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_15 ),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(\current_shift_inst.timer_s1.counter_cry_23 ),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_9_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_9_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_21_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .carryinitout(bfn_9_21_0_));
    defparam IN_MUX_bfv_8_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_21_0_));
    defparam IN_MUX_bfv_8_22_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_22_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .carryinitout(bfn_8_22_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .carryinitout(bfn_13_20_0_));
    ICE_GB delay_tr_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21604),
            .GLOBALBUFFEROUTPUT(delay_tr_input_c_g));
    ICE_GB delay_hc_input_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__21580),
            .GLOBALBUFFEROUTPUT(delay_hc_input_c_g));
    ICE_GB \phase_controller_inst1.stoper_tr.running_RNI6D081_0  (
            .USERSIGNALTOGLOBALBUFFER(N__30499),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst1.stoper_tr.un2_start_0_g ));
    ICE_GB \phase_controller_inst2.stoper_tr.running_RNI96ON_0  (
            .USERSIGNALTOGLOBALBUFFER(N__29281),
            .GLOBALBUFFEROUTPUT(\phase_controller_inst2.stoper_tr.un2_start_0_g ));
    ICE_GB \current_shift_inst.timer_s1.running_RNII51H_0  (
            .USERSIGNALTOGLOBALBUFFER(N__47017),
            .GLOBALBUFFEROUTPUT(\current_shift_inst.timer_s1.N_163_i_g ));
    defparam osc.CLKHF_DIV="0b10";
    SB_HFOSC osc (
            .CLKHFPU(N__51292),
            .CLKHFEN(N__51293),
            .CLKHF(clk_12mhz));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_14_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_0_c_inv_LC_1_14_0  (
            .in0(N__21868),
            .in1(N__21856),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_0 ),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_14_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_1_c_inv_LC_1_14_1  (
            .in0(_gnd_net_),
            .in1(N__21838),
            .in2(_gnd_net_),
            .in3(N__21850),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_14_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_14_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_2_c_inv_LC_1_14_2  (
            .in0(N__21832),
            .in1(N__21820),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_14_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_3_c_inv_LC_1_14_3  (
            .in0(N__21814),
            .in1(N__21802),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_14_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_4_c_inv_LC_1_14_4  (
            .in0(_gnd_net_),
            .in1(N__21784),
            .in2(_gnd_net_),
            .in3(N__21796),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_14_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_5_c_inv_LC_1_14_5  (
            .in0(_gnd_net_),
            .in1(N__21766),
            .in2(_gnd_net_),
            .in3(N__21778),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_14_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_6_c_inv_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__22000),
            .in2(_gnd_net_),
            .in3(N__22012),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_14_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_7_c_inv_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__21982),
            .in2(_gnd_net_),
            .in3(N__21994),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_8_c_inv_LC_1_15_0  (
            .in0(_gnd_net_),
            .in1(N__21964),
            .in2(_gnd_net_),
            .in3(N__21976),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_8 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_9_c_inv_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__21946),
            .in2(_gnd_net_),
            .in3(N__21958),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_8 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_10_c_inv_LC_1_15_2  (
            .in0(_gnd_net_),
            .in1(N__21928),
            .in2(_gnd_net_),
            .in3(N__21940),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_10 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_9 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_11_c_inv_LC_1_15_3  (
            .in0(_gnd_net_),
            .in1(N__21910),
            .in2(_gnd_net_),
            .in3(N__21922),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_11 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_10 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_12_c_inv_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__21892),
            .in2(_gnd_net_),
            .in3(N__21904),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_12 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_11 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_13_c_inv_LC_1_15_5  (
            .in0(_gnd_net_),
            .in1(N__21874),
            .in2(_gnd_net_),
            .in3(N__21886),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_13 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_12 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_14_c_inv_LC_1_15_6  (
            .in0(_gnd_net_),
            .in1(N__22036),
            .in2(_gnd_net_),
            .in3(N__22048),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_14 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_13 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_15_c_LC_1_15_7  (
            .in0(_gnd_net_),
            .in1(N__22198),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_14 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(N__22159),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_16_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_RNIL8HR_LC_1_16_1  (
            .in0(_gnd_net_),
            .in1(N__22264),
            .in2(_gnd_net_),
            .in3(N__22030),
            .lcout(\pwm_generator_inst.un22_threshold_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_16 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_17_c_RNINCJR_LC_1_16_2  (
            .in0(_gnd_net_),
            .in1(N__22234),
            .in2(_gnd_net_),
            .in3(N__22027),
            .lcout(\pwm_generator_inst.un18_threshold1_18 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_17 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_18_c_RNIPGLR_LC_1_16_3  (
            .in0(_gnd_net_),
            .in1(N__22072),
            .in2(_gnd_net_),
            .in3(N__22024),
            .lcout(\pwm_generator_inst.un18_threshold1_19 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_18 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_16_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_19_c_RNIRKNR_LC_1_16_4  (
            .in0(_gnd_net_),
            .in1(N__22249),
            .in2(_gnd_net_),
            .in3(N__22021),
            .lcout(\pwm_generator_inst.un18_threshold1_20 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_19 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_16_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_20_c_RNIK7IS_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__22066),
            .in2(_gnd_net_),
            .in3(N__22018),
            .lcout(\pwm_generator_inst.un18_threshold1_21 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_20 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_16_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_21_c_RNIMBKS_LC_1_16_6  (
            .in0(_gnd_net_),
            .in1(N__22060),
            .in2(_gnd_net_),
            .in3(N__22015),
            .lcout(\pwm_generator_inst.un18_threshold1_22 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_21 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_16_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_22_c_RNIOFMS_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(N__22054),
            .in2(_gnd_net_),
            .in3(N__22084),
            .lcout(\pwm_generator_inst.un18_threshold1_23 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_22 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_23_c_RNIQJOS_LC_1_17_0  (
            .in0(_gnd_net_),
            .in1(N__22240),
            .in2(_gnd_net_),
            .in3(N__22081),
            .lcout(\pwm_generator_inst.un18_threshold1_24 ),
            .ltout(),
            .carryin(bfn_1_17_0_),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_24_c_RNISNQS_LC_1_17_1  (
            .in0(_gnd_net_),
            .in1(N__22255),
            .in2(_gnd_net_),
            .in3(N__22078),
            .lcout(\pwm_generator_inst.un18_threshold1_25 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un18_threshold_1_cry_24 ),
            .carryout(\pwm_generator_inst.un18_threshold_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_17_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_17_2 .LUT_INIT=16'b0110101010100110;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_25_c_RNIK5UE2_LC_1_17_2  (
            .in0(N__22657),
            .in1(N__23393),
            .in2(N__23494),
            .in3(N__22075),
            .lcout(\pwm_generator_inst.N_188_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_1_17_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_1_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_1_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_0_LC_1_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23070),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_1_17_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_1_17_4 .LUT_INIT=16'b0111010010111000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_6_c_RNI1I2H3_LC_1_17_4  (
            .in0(N__23509),
            .in1(N__23392),
            .in2(N__22321),
            .in3(N__23523),
            .lcout(\pwm_generator_inst.N_186_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_17_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_0_LC_1_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23028),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_0_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23295),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_1_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_1_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_0_LC_1_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23007),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_18_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_0_LC_1_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23469),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_1_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_1_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_1_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_0_LC_1_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23457),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_18_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_0_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23046),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_1_18_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_1_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_0_LC_1_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22317),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_18_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_0_LC_1_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23343),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_19_0 .LUT_INIT=16'b1100001111000011;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_15_c_RNO_LC_1_19_0  (
            .in0(_gnd_net_),
            .in1(N__22225),
            .in2(N__22213),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_15 ),
            .ltout(),
            .carryin(bfn_1_19_0_),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_19_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_19_1 .LUT_INIT=16'b0011110011000011;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_RNO_LC_1_19_1  (
            .in0(_gnd_net_),
            .in1(N__22189),
            .in2(N__22177),
            .in3(N__22150),
            .lcout(\pwm_generator_inst.un18_threshold_1_axb_16 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_19_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPO_LC_1_19_2  (
            .in0(_gnd_net_),
            .in1(N__22147),
            .in2(N__22135),
            .in3(N__22117),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_1_c_RNIJNPOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_19_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQO_LC_1_19_3  (
            .in0(_gnd_net_),
            .in1(N__22114),
            .in2(N__22102),
            .in3(N__22087),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_2_c_RNIKPQOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_19_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRRO_LC_1_19_4  (
            .in0(_gnd_net_),
            .in1(N__22504),
            .in2(N__22492),
            .in3(N__22477),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_3_c_RNILRROZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_19_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSO_LC_1_19_5  (
            .in0(_gnd_net_),
            .in1(N__22474),
            .in2(N__22462),
            .in3(N__22447),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_4_c_RNIMTSOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_19_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_19_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTO_LC_1_19_6  (
            .in0(_gnd_net_),
            .in1(N__22444),
            .in2(N__22432),
            .in3(N__22417),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_5_c_RNINVTOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_19_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VO_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__22414),
            .in2(N__22402),
            .in3(N__22387),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_6_c_RNIO1VOZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_20_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30P_LC_1_20_0  (
            .in0(_gnd_net_),
            .in1(N__22384),
            .in2(N__22369),
            .in3(N__22354),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_7_c_RNIP30PZ0 ),
            .ltout(),
            .carryin(bfn_1_20_0_),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_20_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51P_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__22351),
            .in2(N__22336),
            .in3(N__22300),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_8_c_RNIQ51PZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_20_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72P_LC_1_20_2  (
            .in0(_gnd_net_),
            .in1(N__22297),
            .in2(N__22282),
            .in3(N__22267),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_9_c_RNIR72PZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_20_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPF_LC_1_20_3  (
            .in0(_gnd_net_),
            .in1(N__22579),
            .in2(N__22672),
            .in3(N__22648),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_10_c_RNI3NPFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_20_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_20_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_20_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_12_c_LC_1_20_4  (
            .in0(_gnd_net_),
            .in1(N__22645),
            .in2(N__22590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_11 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_20_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_20_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_13_c_LC_1_20_5  (
            .in0(_gnd_net_),
            .in1(N__22583),
            .in2(N__22633),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_12 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_20_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_20_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_20_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_14_c_LC_1_20_6  (
            .in0(_gnd_net_),
            .in1(N__22618),
            .in2(N__22591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_13 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_20_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_20_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_15_c_LC_1_20_7  (
            .in0(_gnd_net_),
            .in1(N__22587),
            .in2(N__22603),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\pwm_generator_inst.un5_threshold_add_1_cry_14 ),
            .carryout(\pwm_generator_inst.un5_threshold_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_21_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJ1_LC_1_21_0  (
            .in0(_gnd_net_),
            .in1(N__22510),
            .in2(_gnd_net_),
            .in3(N__22606),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNI1OUJZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_21_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_21_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_21_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNO_LC_1_21_4  (
            .in0(N__22589),
            .in1(N__23121),
            .in2(_gnd_net_),
            .in3(N__22533),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_1_22_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_1_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \pwm_generator_inst.un5_threshold_add_1_axb_16_1_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(N__22588),
            .in2(_gnd_net_),
            .in3(N__22546),
            .lcout(),
            .ltout(\pwm_generator_inst.un5_threshold_add_1_axb_16Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_1_22_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_1_22_4 .LUT_INIT=16'b0101101010010110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNICSGJ1_LC_1_22_4  (
            .in0(N__23086),
            .in1(N__23122),
            .in2(N__22537),
            .in3(N__22534),
            .lcout(\pwm_generator_inst.un5_threshold_add_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_23_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_23_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_LC_1_23_0  (
            .in0(_gnd_net_),
            .in1(N__51949),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_23_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_23_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_23_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_23_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_0_c_RNI53CC_LC_1_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22918),
            .in3(N__22885),
            .lcout(\pwm_generator_inst.un3_threshold_cry_0_c_RNI53CCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_0 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_23_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_1_c_RNI65DC_LC_1_23_2  (
            .in0(_gnd_net_),
            .in1(N__50900),
            .in2(N__22882),
            .in3(N__22849),
            .lcout(\pwm_generator_inst.un3_threshold_cry_1_c_RNI65DCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_1 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_23_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_23_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_2_c_RNI77EC_LC_1_23_3  (
            .in0(_gnd_net_),
            .in1(N__22846),
            .in2(N__51060),
            .in3(N__22807),
            .lcout(\pwm_generator_inst.un3_threshold_cry_2_c_RNI77ECZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_2 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_23_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_3_c_RNI89FC_LC_1_23_4  (
            .in0(_gnd_net_),
            .in1(N__22804),
            .in2(_gnd_net_),
            .in3(N__22777),
            .lcout(\pwm_generator_inst.un3_threshold_cry_3_c_RNI89FCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_3 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_23_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGC_LC_1_23_5  (
            .in0(_gnd_net_),
            .in1(N__22774),
            .in2(N__51061),
            .in3(N__22738),
            .lcout(\pwm_generator_inst.un3_threshold_cry_4_c_RNI9BGCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_4 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_23_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_5_c_RNIADHC_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(N__22735),
            .in2(_gnd_net_),
            .in3(N__22708),
            .lcout(\pwm_generator_inst.un3_threshold_cry_5_c_RNIADHCZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_5 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_23_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_23_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_6_c_RNIBFIC_LC_1_23_7  (
            .in0(_gnd_net_),
            .in1(N__22705),
            .in2(_gnd_net_),
            .in3(N__22675),
            .lcout(\pwm_generator_inst.un3_threshold_cry_6_c_RNIBFICZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_6 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_24_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_24_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FO_LC_1_24_0  (
            .in0(_gnd_net_),
            .in1(N__28216),
            .in2(_gnd_net_),
            .in3(N__22984),
            .lcout(\pwm_generator_inst.un3_threshold_cry_7_c_RNIA8FOZ0 ),
            .ltout(),
            .carryin(bfn_1_24_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_24_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_8_c_RNIQDI8_LC_1_24_1  (
            .in0(_gnd_net_),
            .in1(N__28156),
            .in2(_gnd_net_),
            .in3(N__22975),
            .lcout(\pwm_generator_inst.un3_threshold_cry_8_c_RNIQDIZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_8 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_24_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_24_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_24_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_9_c_RNISHK8_LC_1_24_2  (
            .in0(_gnd_net_),
            .in1(N__28108),
            .in2(_gnd_net_),
            .in3(N__22966),
            .lcout(\pwm_generator_inst.un3_threshold_cry_9_c_RNISHKZ0Z8 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_9 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_24_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_24_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_24_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_10_c_RNI59G7_LC_1_24_3  (
            .in0(_gnd_net_),
            .in1(N__28051),
            .in2(_gnd_net_),
            .in3(N__22957),
            .lcout(\pwm_generator_inst.un3_threshold_cry_10_c_RNI59GZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_10 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_24_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_24_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_11_c_RNI7DI7_LC_1_24_4  (
            .in0(_gnd_net_),
            .in1(N__28015),
            .in2(_gnd_net_),
            .in3(N__22948),
            .lcout(\pwm_generator_inst.un3_threshold_cry_11_c_RNI7DIZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_11 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_24_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_24_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_12_c_RNI9HK7_LC_1_24_5  (
            .in0(_gnd_net_),
            .in1(N__27991),
            .in2(_gnd_net_),
            .in3(N__22939),
            .lcout(\pwm_generator_inst.un3_threshold_cry_12_c_RNI9HKZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_12 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_24_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_24_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_13_c_RNIBLM7_LC_1_24_6  (
            .in0(_gnd_net_),
            .in1(N__27961),
            .in2(_gnd_net_),
            .in3(N__22930),
            .lcout(\pwm_generator_inst.un3_threshold_cry_13_c_RNIBLMZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_13 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_24_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_24_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_14_c_RNIDPO7_LC_1_24_7  (
            .in0(_gnd_net_),
            .in1(N__27928),
            .in2(_gnd_net_),
            .in3(N__22921),
            .lcout(\pwm_generator_inst.un3_threshold_cry_14_c_RNIDPOZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_14 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_25_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQ7_LC_1_25_0  (
            .in0(_gnd_net_),
            .in1(N__28501),
            .in2(_gnd_net_),
            .in3(N__23143),
            .lcout(\pwm_generator_inst.un3_threshold_cry_15_c_RNIFTQZ0Z7 ),
            .ltout(),
            .carryin(bfn_1_25_0_),
            .carryout(\pwm_generator_inst.un3_threshold_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_25_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un3_threshold_cry_16_c_RNIH1T7_LC_1_25_1  (
            .in0(_gnd_net_),
            .in1(N__28462),
            .in2(_gnd_net_),
            .in3(N__23134),
            .lcout(\pwm_generator_inst.un3_threshold_cry_16_c_RNIH1TZ0Z7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_16 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_25_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFD_LC_1_25_2  (
            .in0(_gnd_net_),
            .in1(N__28435),
            .in2(_gnd_net_),
            .in3(N__23125),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_10_s_RNIQFDZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_17 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_25_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJF_LC_1_25_3  (
            .in0(_gnd_net_),
            .in1(N__28312),
            .in2(_gnd_net_),
            .in3(N__23107),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_s_RNISJFZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un3_threshold_cry_18 ),
            .carryout(\pwm_generator_inst.un3_threshold_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_25_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSON_LC_1_25_4  (
            .in0(N__23104),
            .in1(N__28291),
            .in2(N__28414),
            .in3(N__23089),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_c_RNIBSONZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_2_15_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_2_15_0 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_1_c_RNIMQKF3_LC_2_15_0  (
            .in0(N__23266),
            .in1(N__23278),
            .in2(N__23077),
            .in3(N__23383),
            .lcout(\pwm_generator_inst.N_181_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_2_15_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_2_15_2 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_2_c_RNIQ2PF3_LC_2_15_2  (
            .in0(N__23253),
            .in1(N__23239),
            .in2(N__23056),
            .in3(N__23384),
            .lcout(\pwm_generator_inst.N_182_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_2_15_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_2_15_4 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_3_c_RNILPLG3_LC_2_15_4  (
            .in0(N__23215),
            .in1(N__23227),
            .in2(N__23035),
            .in3(N__23385),
            .lcout(\pwm_generator_inst.N_183_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_15_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_15_5 .LUT_INIT=16'b0111110100101000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_5_c_RNIT9UG3_LC_2_15_5  (
            .in0(N__23386),
            .in1(N__23179),
            .in2(N__23167),
            .in3(N__23011),
            .lcout(\pwm_generator_inst.N_185_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_2_16_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_2_16_1 .LUT_INIT=16'b0110011011110000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_4_c_RNIP1QG3_LC_2_16_1  (
            .in0(N__23188),
            .in1(N__23202),
            .in2(N__23302),
            .in3(N__23394),
            .lcout(\pwm_generator_inst.N_184_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_0_c_LC_2_17_0  (
            .in0(_gnd_net_),
            .in1(N__23481),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_17_0_),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_0_THRU_LUT4_0_LC_2_17_1  (
            .in0(_gnd_net_),
            .in1(N__51062),
            .in2(N__23412),
            .in3(N__23281),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_0 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_1_THRU_LUT4_0_LC_2_17_2  (
            .in0(_gnd_net_),
            .in1(N__23277),
            .in2(N__51289),
            .in3(N__23257),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_1 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_2_THRU_LUT4_0_LC_2_17_3  (
            .in0(_gnd_net_),
            .in1(N__51066),
            .in2(N__23254),
            .in3(N__23230),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_2 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_3_THRU_LUT4_0_LC_2_17_4  (
            .in0(_gnd_net_),
            .in1(N__23226),
            .in2(N__51290),
            .in3(N__23206),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_3 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_4_THRU_LUT4_0_LC_2_17_5  (
            .in0(_gnd_net_),
            .in1(N__51070),
            .in2(N__23203),
            .in3(N__23182),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_4 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_5_THRU_LUT4_0_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__23178),
            .in2(N__51291),
            .in3(N__23155),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_5 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_6_THRU_LUT4_0_LC_2_17_7  (
            .in0(_gnd_net_),
            .in1(N__51074),
            .in2(N__23524),
            .in3(N__23503),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\pwm_generator_inst.un22_threshold_1_cry_6 ),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_7_THRU_LUT4_0_LC_2_18_0  (
            .in0(_gnd_net_),
            .in1(N__50989),
            .in2(N__23439),
            .in3(N__23500),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_18_0_),
            .carryout(\pwm_generator_inst.un22_threshold_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_18_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_8_THRU_LUT4_0_LC_2_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23497),
            .lcout(\pwm_generator_inst.un22_threshold_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_18_3 .C_ON=1'b0;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \pwm_generator_inst.un18_threshold_1_cry_16_c_RNI9O983_LC_2_18_3  (
            .in0(N__23387),
            .in1(N__23485),
            .in2(_gnd_net_),
            .in3(N__23470),
            .lcout(\pwm_generator_inst.N_179_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_18_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_18_4 .LUT_INIT=16'b0010111011100010;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_7_c_RNI5Q6H3_LC_2_18_4  (
            .in0(N__23458),
            .in1(N__23391),
            .in2(N__23440),
            .in3(N__23425),
            .lcout(\pwm_generator_inst.N_187_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_18_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_18_5 .LUT_INIT=16'b0110111101100000;
    LogicCell40 \pwm_generator_inst.un22_threshold_1_cry_0_c_RNIIIGF3_LC_2_18_5  (
            .in0(N__23419),
            .in1(N__23413),
            .in2(N__23395),
            .in3(N__23344),
            .lcout(\pwm_generator_inst.N_180_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_17_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_17_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_0_c_inv_LC_3_17_0  (
            .in0(N__23759),
            .in1(N__23323),
            .in2(N__23332),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_0 ),
            .ltout(),
            .carryin(bfn_3_17_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_17_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_17_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_1_c_inv_LC_3_17_1  (
            .in0(N__23739),
            .in1(N__23308),
            .in2(N__23317),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_0 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_17_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_2_c_inv_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__23662),
            .in2(N__23677),
            .in3(N__23717),
            .lcout(\pwm_generator_inst.counter_i_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_1 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_17_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_3_c_inv_LC_3_17_3  (
            .in0(N__23696),
            .in1(N__23641),
            .in2(N__23656),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.counter_i_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_2 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_17_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_4_c_inv_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__23620),
            .in2(N__23635),
            .in3(N__23972),
            .lcout(\pwm_generator_inst.counter_i_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_3 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_17_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_5_c_inv_LC_3_17_5  (
            .in0(_gnd_net_),
            .in1(N__23614),
            .in2(N__23608),
            .in3(N__23952),
            .lcout(\pwm_generator_inst.counter_i_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_4 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_17_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_6_c_inv_LC_3_17_6  (
            .in0(_gnd_net_),
            .in1(N__23584),
            .in2(N__23599),
            .in3(N__23930),
            .lcout(\pwm_generator_inst.counter_i_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_5 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_17_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_7_c_inv_LC_3_17_7  (
            .in0(_gnd_net_),
            .in1(N__23566),
            .in2(N__23578),
            .in3(N__23909),
            .lcout(\pwm_generator_inst.counter_i_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_6 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_8_c_inv_LC_3_18_0  (
            .in0(_gnd_net_),
            .in1(N__23551),
            .in2(N__23560),
            .in3(N__23888),
            .lcout(\pwm_generator_inst.counter_i_8 ),
            .ltout(),
            .carryin(bfn_3_18_0_),
            .carryout(\pwm_generator_inst.un14_counter_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pwm_generator_inst.un14_counter_cry_9_c_inv_LC_3_18_1  (
            .in0(_gnd_net_),
            .in1(N__23530),
            .in2(N__23545),
            .in3(N__23819),
            .lcout(\pwm_generator_inst.counter_i_9 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un14_counter_cry_8 ),
            .carryout(\pwm_generator_inst.un14_counter_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.pwm_out_LC_3_18_2 .C_ON=1'b0;
    defparam \pwm_generator_inst.pwm_out_LC_3_18_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.pwm_out_LC_3_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.pwm_out_LC_3_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23800),
            .lcout(pwm_output_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52609),
            .ce(),
            .sr(N__52268));
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_4_17_0 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNITBL3_9_LC_4_17_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNITBL3_9_LC_4_17_0  (
            .in0(N__23890),
            .in1(N__23821),
            .in2(_gnd_net_),
            .in3(N__23951),
            .lcout(\pwm_generator_inst.un1_counterlto9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_4_17_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_4_17_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIRPD2_0_LC_4_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIRPD2_0_LC_4_17_5  (
            .in0(_gnd_net_),
            .in1(N__23760),
            .in2(_gnd_net_),
            .in3(N__23738),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlto2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_4_17_6 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_4_17_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIBO26_2_LC_4_17_6 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \pwm_generator_inst.counter_RNIBO26_2_LC_4_17_6  (
            .in0(N__23973),
            .in1(N__23697),
            .in2(N__23773),
            .in3(N__23718),
            .lcout(),
            .ltout(\pwm_generator_inst.un1_counterlt9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_4_17_7 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.counter_RNIFA6C_6_LC_4_17_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \pwm_generator_inst.counter_RNIFA6C_6_LC_4_17_7  (
            .in0(N__23770),
            .in1(N__23910),
            .in2(N__23764),
            .in3(N__23932),
            .lcout(\pwm_generator_inst.un1_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.counter_0_LC_4_18_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_0_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_0_LC_4_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_0_LC_4_18_0  (
            .in0(N__23861),
            .in1(N__23761),
            .in2(_gnd_net_),
            .in3(N__23743),
            .lcout(\pwm_generator_inst.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_4_18_0_),
            .carryout(\pwm_generator_inst.counter_cry_0 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_1_LC_4_18_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_1_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_1_LC_4_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_1_LC_4_18_1  (
            .in0(N__23857),
            .in1(N__23740),
            .in2(_gnd_net_),
            .in3(N__23722),
            .lcout(\pwm_generator_inst.counterZ0Z_1 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_0 ),
            .carryout(\pwm_generator_inst.counter_cry_1 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_2_LC_4_18_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_2_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_2_LC_4_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_2_LC_4_18_2  (
            .in0(N__23862),
            .in1(N__23719),
            .in2(_gnd_net_),
            .in3(N__23701),
            .lcout(\pwm_generator_inst.counterZ0Z_2 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_1 ),
            .carryout(\pwm_generator_inst.counter_cry_2 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_3_LC_4_18_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_3_LC_4_18_3 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_3_LC_4_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_3_LC_4_18_3  (
            .in0(N__23858),
            .in1(N__23698),
            .in2(_gnd_net_),
            .in3(N__23680),
            .lcout(\pwm_generator_inst.counterZ0Z_3 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_2 ),
            .carryout(\pwm_generator_inst.counter_cry_3 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_4_LC_4_18_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_4_LC_4_18_4 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_4_LC_4_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_4_LC_4_18_4  (
            .in0(N__23863),
            .in1(N__23974),
            .in2(_gnd_net_),
            .in3(N__23956),
            .lcout(\pwm_generator_inst.counterZ0Z_4 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_3 ),
            .carryout(\pwm_generator_inst.counter_cry_4 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_5_LC_4_18_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_5_LC_4_18_5 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_5_LC_4_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_5_LC_4_18_5  (
            .in0(N__23859),
            .in1(N__23953),
            .in2(_gnd_net_),
            .in3(N__23935),
            .lcout(\pwm_generator_inst.counterZ0Z_5 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_4 ),
            .carryout(\pwm_generator_inst.counter_cry_5 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_6_LC_4_18_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_6_LC_4_18_6 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_6_LC_4_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_6_LC_4_18_6  (
            .in0(N__23864),
            .in1(N__23931),
            .in2(_gnd_net_),
            .in3(N__23914),
            .lcout(\pwm_generator_inst.counterZ0Z_6 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_5 ),
            .carryout(\pwm_generator_inst.counter_cry_6 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_7_LC_4_18_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_7_LC_4_18_7 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_7_LC_4_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_7_LC_4_18_7  (
            .in0(N__23860),
            .in1(N__23911),
            .in2(_gnd_net_),
            .in3(N__23893),
            .lcout(\pwm_generator_inst.counterZ0Z_7 ),
            .ltout(),
            .carryin(\pwm_generator_inst.counter_cry_6 ),
            .carryout(\pwm_generator_inst.counter_cry_7 ),
            .clk(N__52601),
            .ce(),
            .sr(N__52266));
    defparam \pwm_generator_inst.counter_8_LC_4_19_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.counter_8_LC_4_19_0 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_8_LC_4_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \pwm_generator_inst.counter_8_LC_4_19_0  (
            .in0(N__23866),
            .in1(N__23889),
            .in2(_gnd_net_),
            .in3(N__23869),
            .lcout(\pwm_generator_inst.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_4_19_0_),
            .carryout(\pwm_generator_inst.counter_cry_8 ),
            .clk(N__52594),
            .ce(),
            .sr(N__52269));
    defparam \pwm_generator_inst.counter_9_LC_4_19_1 .C_ON=1'b0;
    defparam \pwm_generator_inst.counter_9_LC_4_19_1 .SEQ_MODE=4'b1010;
    defparam \pwm_generator_inst.counter_9_LC_4_19_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \pwm_generator_inst.counter_9_LC_4_19_1  (
            .in0(N__23820),
            .in1(N__23865),
            .in2(_gnd_net_),
            .in3(N__23824),
            .lcout(\pwm_generator_inst.counterZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52594),
            .ce(),
            .sr(N__52269));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_15_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_15_0  (
            .in0(N__24016),
            .in1(N__31810),
            .in2(N__31840),
            .in3(N__24007),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_5_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_5_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_16_LC_5_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_16_LC_5_15_1  (
            .in0(N__25704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52621),
            .ce(N__36636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_5_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_5_15_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_16_LC_5_15_2  (
            .in0(N__24015),
            .in1(N__31809),
            .in2(N__31839),
            .in3(N__24006),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_5_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_5_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_17_LC_5_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_17_LC_5_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25680),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52621),
            .ce(N__36636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_15_4 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_15_4  (
            .in0(N__32047),
            .in1(N__32067),
            .in2(N__23997),
            .in3(N__23983),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_5_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_5_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_18_LC_5_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_18_LC_5_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25656),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52621),
            .ce(N__36636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_5_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_5_15_6 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_18_LC_5_15_6  (
            .in0(N__32046),
            .in1(N__32068),
            .in2(N__23998),
            .in3(N__23982),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_5_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_19_LC_5_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_19_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25788),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52621),
            .ce(N__36636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_16_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_25_LC_5_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28684),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52610),
            .ce(N__32635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_5_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_5_16_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_27_LC_5_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_27_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28636),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52610),
            .ce(N__32635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_5_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_26_LC_5_16_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_26_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(N__28660),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52610),
            .ce(N__32635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_5_16_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_24_LC_5_16_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_24_LC_5_16_5  (
            .in0(N__28279),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52610),
            .ce(N__32635),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_5_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_21_LC_5_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_21_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25768),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52602),
            .ce(N__36637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_18_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_18_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_16_LC_5_18_0  (
            .in0(N__26239),
            .in1(N__24049),
            .in2(N__26215),
            .in3(N__24058),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_5_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_16_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_16_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25711),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52595),
            .ce(N__32636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_5_18_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_5_18_2 .LUT_INIT=16'b1100111101001101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_16_LC_5_18_2  (
            .in0(N__26238),
            .in1(N__24048),
            .in2(N__26214),
            .in3(N__24057),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_5_18_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_5_18_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_17_LC_5_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_17_LC_5_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25684),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52595),
            .ce(N__32636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_18_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_18_4 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_18_LC_5_18_4  (
            .in0(N__26161),
            .in1(N__26184),
            .in2(N__24039),
            .in3(N__24025),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_5_18_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_5_18_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_18_LC_5_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_18_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25660),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52595),
            .ce(N__32636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_5_18_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_5_18_6 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_18_LC_5_18_6  (
            .in0(N__26160),
            .in1(N__26185),
            .in2(N__24040),
            .in3(N__24024),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_5_18_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_19_LC_5_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_19_LC_5_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25792),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52595),
            .ce(N__32636),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_5_19_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_5_19_0 .LUT_INIT=16'b0100110100001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_24_LC_5_19_0  (
            .in0(N__26458),
            .in1(N__24121),
            .in2(N__26434),
            .in3(N__24109),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_5_19_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_5_19_2 .LUT_INIT=16'b1100111101001101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_24_LC_5_19_2  (
            .in0(N__26457),
            .in1(N__24120),
            .in2(N__26433),
            .in3(N__24108),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_5_19_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_5_19_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_26_LC_5_19_4  (
            .in0(N__24097),
            .in1(N__26374),
            .in2(N__26403),
            .in3(N__24085),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_5_19_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_5_19_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_26_LC_5_19_6  (
            .in0(N__24096),
            .in1(N__26373),
            .in2(N__26404),
            .in3(N__24084),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_5_22_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_5_22_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_5_22_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_5_22_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_0_LC_7_7_0  (
            .in0(N__24335),
            .in1(N__29828),
            .in2(_gnd_net_),
            .in3(N__24073),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_1_LC_7_7_1  (
            .in0(N__24370),
            .in1(N__29783),
            .in2(_gnd_net_),
            .in3(N__24070),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_2_LC_7_7_2  (
            .in0(N__24336),
            .in1(N__24904),
            .in2(_gnd_net_),
            .in3(N__24067),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_3_LC_7_7_3  (
            .in0(N__24371),
            .in1(N__24882),
            .in2(_gnd_net_),
            .in3(N__24064),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_4_LC_7_7_4  (
            .in0(N__24337),
            .in1(N__25139),
            .in2(_gnd_net_),
            .in3(N__24061),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_5_LC_7_7_5  (
            .in0(N__24372),
            .in1(N__25113),
            .in2(_gnd_net_),
            .in3(N__24148),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_6_LC_7_7_6  (
            .in0(N__24338),
            .in1(N__25089),
            .in2(_gnd_net_),
            .in3(N__24145),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_7_LC_7_7_7  (
            .in0(N__24373),
            .in1(N__25065),
            .in2(_gnd_net_),
            .in3(N__24142),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_7 ),
            .clk(N__52656),
            .ce(N__36565),
            .sr(N__52211));
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_8_LC_7_8_0  (
            .in0(N__24342),
            .in1(N__25041),
            .in2(_gnd_net_),
            .in3(N__24139),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_9_LC_7_8_1  (
            .in0(N__24355),
            .in1(N__25020),
            .in2(_gnd_net_),
            .in3(N__24136),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_10_LC_7_8_2  (
            .in0(N__24339),
            .in1(N__24996),
            .in2(_gnd_net_),
            .in3(N__24133),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_11_LC_7_8_3  (
            .in0(N__24352),
            .in1(N__24974),
            .in2(_gnd_net_),
            .in3(N__24130),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_12_LC_7_8_4  (
            .in0(N__24340),
            .in1(N__25329),
            .in2(_gnd_net_),
            .in3(N__24127),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_13_LC_7_8_5  (
            .in0(N__24353),
            .in1(N__25305),
            .in2(_gnd_net_),
            .in3(N__24124),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_14_LC_7_8_6  (
            .in0(N__24341),
            .in1(N__25281),
            .in2(_gnd_net_),
            .in3(N__24175),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_15_LC_7_8_7  (
            .in0(N__24354),
            .in1(N__25257),
            .in2(_gnd_net_),
            .in3(N__24172),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_15 ),
            .clk(N__52651),
            .ce(N__36564),
            .sr(N__52218));
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_16_LC_7_9_0  (
            .in0(N__24364),
            .in1(N__25233),
            .in2(_gnd_net_),
            .in3(N__24169),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_17_LC_7_9_1  (
            .in0(N__24360),
            .in1(N__25212),
            .in2(_gnd_net_),
            .in3(N__24166),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_18_LC_7_9_2  (
            .in0(N__24365),
            .in1(N__25188),
            .in2(_gnd_net_),
            .in3(N__24163),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_19_LC_7_9_3  (
            .in0(N__24361),
            .in1(N__25166),
            .in2(_gnd_net_),
            .in3(N__24160),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_20_LC_7_9_4  (
            .in0(N__24366),
            .in1(N__25548),
            .in2(_gnd_net_),
            .in3(N__24157),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_21_LC_7_9_5  (
            .in0(N__24362),
            .in1(N__25524),
            .in2(_gnd_net_),
            .in3(N__24154),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_22_LC_7_9_6  (
            .in0(N__24367),
            .in1(N__25500),
            .in2(_gnd_net_),
            .in3(N__24151),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_23_LC_7_9_7  (
            .in0(N__24363),
            .in1(N__25476),
            .in2(_gnd_net_),
            .in3(N__24205),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_23 ),
            .clk(N__52644),
            .ce(N__36557),
            .sr(N__52224));
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_24_LC_7_10_0  (
            .in0(N__24356),
            .in1(N__25452),
            .in2(_gnd_net_),
            .in3(N__24202),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_7_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .clk(N__52639),
            .ce(N__36556),
            .sr(N__52233));
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_25_LC_7_10_1  (
            .in0(N__24368),
            .in1(N__25428),
            .in2(_gnd_net_),
            .in3(N__24199),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .clk(N__52639),
            .ce(N__36556),
            .sr(N__52233));
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_26_LC_7_10_2  (
            .in0(N__24357),
            .in1(N__25392),
            .in2(_gnd_net_),
            .in3(N__24196),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .clk(N__52639),
            .ce(N__36556),
            .sr(N__52233));
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_27_LC_7_10_3  (
            .in0(N__24369),
            .in1(N__25356),
            .in2(_gnd_net_),
            .in3(N__24193),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .clk(N__52639),
            .ce(N__36556),
            .sr(N__52233));
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_28_LC_7_10_4  (
            .in0(N__24358),
            .in1(N__25408),
            .in2(_gnd_net_),
            .in3(N__24190),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.counter_cry_28 ),
            .clk(N__52639),
            .ce(N__36556),
            .sr(N__52233));
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.counter_29_LC_7_10_5  (
            .in0(N__25372),
            .in1(N__24359),
            .in2(_gnd_net_),
            .in3(N__24187),
            .lcout(\delay_measurement_inst.delay_tr_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52639),
            .ce(N__36556),
            .sr(N__52233));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_7_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_7_11_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5GPBB_27_LC_7_11_0  (
            .in0(N__33752),
            .in1(N__24184),
            .in2(_gnd_net_),
            .in3(N__27106),
            .lcout(elapsed_time_ns_1_RNI5GPBB_0_27),
            .ltout(elapsed_time_ns_1_RNI5GPBB_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_7_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_7_11_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_27_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24178),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_11_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7IPBB_29_LC_7_11_2  (
            .in0(N__33753),
            .in1(N__24235),
            .in2(_gnd_net_),
            .in3(N__27031),
            .lcout(elapsed_time_ns_1_RNI7IPBB_0_29),
            .ltout(elapsed_time_ns_1_RNI7IPBB_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_7_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_7_11_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_29_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24229),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_7_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_7_11_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIT6OBB_10_LC_7_11_4  (
            .in0(N__33750),
            .in1(N__25612),
            .in2(_gnd_net_),
            .in3(N__26956),
            .lcout(elapsed_time_ns_1_RNIT6OBB_0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJI91B_7_LC_7_11_5  (
            .in0(N__33749),
            .in1(N__24226),
            .in2(_gnd_net_),
            .in3(N__29628),
            .lcout(elapsed_time_ns_1_RNIJI91B_0_7),
            .ltout(elapsed_time_ns_1_RNIJI91B_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_7_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_7_11_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_7_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24220),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_11_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1CPBB_23_LC_7_11_7  (
            .in0(N__24217),
            .in1(N__27018),
            .in2(_gnd_net_),
            .in3(N__33751),
            .lcout(elapsed_time_ns_1_RNI1CPBB_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_12_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_0_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__36699),
            .in2(_gnd_net_),
            .in3(N__36740),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52626),
            .ce(N__32596),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_12_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI1BOBB_14_LC_7_12_2  (
            .in0(N__26914),
            .in1(N__25570),
            .in2(_gnd_net_),
            .in3(N__33776),
            .lcout(elapsed_time_ns_1_RNI1BOBB_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_7_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_7_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_23_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24216),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2COBB_15_LC_7_12_6  (
            .in0(N__26998),
            .in1(N__25591),
            .in2(_gnd_net_),
            .in3(N__33777),
            .lcout(elapsed_time_ns_1_RNI2COBB_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNI2DO8_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36502),
            .lcout(\delay_measurement_inst.delay_tr_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_7_13_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_7_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6GOBB_19_LC_7_13_6  (
            .in0(N__24244),
            .in1(N__27310),
            .in2(_gnd_net_),
            .in3(N__33778),
            .lcout(elapsed_time_ns_1_RNI6GOBB_0_19),
            .ltout(elapsed_time_ns_1_RNI6GOBB_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_7_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_7_13_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_19_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24238),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_5_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30090),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_1_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30120),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_3_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30264),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_6_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30105),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_7_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30057),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_7_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_15_LC_7_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_15_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34227),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_7_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_14_LC_7_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_14_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34281),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_4_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30042),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52611),
            .ce(N__32615),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_7_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_2_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_2_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30028),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_10_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34107),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_7_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_13_LC_7_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_13_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30069),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_15_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_8_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__34167),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_11_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34194),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_9_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34137),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_7_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_7_15_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_12_LC_7_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_12_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34254),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_15_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_15_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_22_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32754),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52603),
            .ce(N__32637),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_16_0 .LUT_INIT=16'b0100110101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_20_LC_7_16_0  (
            .in0(N__26109),
            .in1(N__24436),
            .in2(N__26136),
            .in3(N__24445),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_20_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32154),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52596),
            .ce(N__32619),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_16_2 .LUT_INIT=16'b1101110101001101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_20_LC_7_16_2  (
            .in0(N__26110),
            .in1(N__24435),
            .in2(N__26137),
            .in3(N__24444),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_21_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25761),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52596),
            .ce(N__32619),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_16_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_22_LC_7_16_4  (
            .in0(N__26059),
            .in1(N__24427),
            .in2(N__26089),
            .in3(N__24418),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_16_6 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_22_LC_7_16_6  (
            .in0(N__26058),
            .in1(N__24426),
            .in2(N__26088),
            .in3(N__24417),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_23_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32679),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52596),
            .ce(N__32619),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_7_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_7_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__24409),
            .in2(N__24400),
            .in3(N__25893),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_0 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_7_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_7_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__24379),
            .in2(N__24391),
            .in3(N__25881),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_7_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_7_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_2_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__24583),
            .in2(N__24595),
            .in3(N__25866),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_7_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_7_17_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_3_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__24565),
            .in2(N__24577),
            .in3(N__25851),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_7_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_7_17_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__24559),
            .in2(N__24544),
            .in3(N__25836),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_7_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_7_17_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_7_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_5_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__24523),
            .in2(N__24535),
            .in3(N__25821),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_7_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_7_17_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__24517),
            .in2(N__24508),
            .in3(N__25806),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_7_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_7_17_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_7_LC_7_17_7  (
            .in0(N__26034),
            .in1(N__24487),
            .in2(N__24499),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_7_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_7_18_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_8_LC_7_18_0  (
            .in0(N__26019),
            .in1(N__24481),
            .in2(N__24472),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_8 ),
            .ltout(),
            .carryin(bfn_7_18_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_7_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_7_18_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_9_LC_7_18_1  (
            .in0(N__26004),
            .in1(N__24451),
            .in2(N__24463),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_7_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_7_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_10_LC_7_18_2  (
            .in0(_gnd_net_),
            .in1(N__24760),
            .in2(N__24751),
            .in3(N__25989),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_7_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_7_18_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_11_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__24730),
            .in2(N__24742),
            .in3(N__25974),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_7_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_7_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_12_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__24724),
            .in2(N__24715),
            .in3(N__25959),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_7_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_7_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_13_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__24706),
            .in2(N__24697),
            .in3(N__25944),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_7_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_7_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_14_LC_7_18_6  (
            .in0(_gnd_net_),
            .in1(N__24673),
            .in2(N__24685),
            .in3(N__25929),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_7_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_7_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_inv_15_LC_7_18_7  (
            .in0(_gnd_net_),
            .in1(N__24667),
            .in2(N__24658),
            .in3(N__26253),
            .lcout(\phase_controller_inst2.stoper_tr.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_7_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_7_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_16_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__24649),
            .in2(N__24637),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_7_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_7_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_18_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__24622),
            .in2(N__24610),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_7_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_7_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_20_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__24865),
            .in2(N__24856),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_7_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_7_19_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_7_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_22_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__24844),
            .in2(N__24832),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_7_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_7_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_24_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__24820),
            .in2(N__24811),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_7_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_7_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_26_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__24799),
            .in2(N__24790),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_7_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_7_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_28_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__24937),
            .in2(N__24946),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_7_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_7_19_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_30_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__24952),
            .in2(N__24772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.un6_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_7_20_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_7_20_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_7_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24775),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_7_20_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_7_20_1 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_30_LC_7_20_1  (
            .in0(N__32658),
            .in1(N__26289),
            .in2(_gnd_net_),
            .in3(N__26309),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_7_20_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_7_20_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_30_LC_7_20_2  (
            .in0(N__26310),
            .in1(N__26288),
            .in2(_gnd_net_),
            .in3(N__32659),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_7_20_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_7_20_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_28_LC_7_20_3  (
            .in0(N__32656),
            .in1(N__26327),
            .in2(_gnd_net_),
            .in3(N__26348),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_2_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_7_20_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_7_20_4 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNO_0_28_LC_7_20_4  (
            .in0(N__26328),
            .in1(N__26349),
            .in2(_gnd_net_),
            .in3(N__32657),
            .lcout(\phase_controller_inst2.stoper_tr.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_7_20_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_7_20_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_tr.un6_running_cry_c_RNI781H_30_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__32556),
            .in2(_gnd_net_),
            .in3(N__29220),
            .lcout(\phase_controller_inst2.stoper_tr.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_7_30_1.C_ON=1'b0;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_7_30_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_7_30_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_clk_12mhz_THRU_LUT4_0_LC_7_30_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24931),
            .lcout(GB_BUFFER_clk_12mhz_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.start_latched_LC_8_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29269),
            .lcout(\phase_controller_inst2.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52652),
            .ce(),
            .sr(N__52199));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_8_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_3_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__24902),
            .in2(N__29835),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_3 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_4_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__24881),
            .in2(N__29790),
            .in3(N__24907),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_5_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__24903),
            .in2(N__25140),
            .in3(N__24889),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_6_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__25112),
            .in2(N__24886),
            .in3(N__25144),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_7_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__25088),
            .in2(N__25141),
            .in3(N__25120),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_8_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__25064),
            .in2(N__25117),
            .in3(N__25096),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_9_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__25040),
            .in2(N__25093),
            .in3(N__25072),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_10_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__25019),
            .in2(N__25069),
            .in3(N__25048),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__52645),
            .ce(N__36478),
            .sr(N__52212));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_11_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__24995),
            .in2(N__25045),
            .in3(N__25024),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_11 ),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_12_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__25021),
            .in2(N__24975),
            .in3(N__25003),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_13_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__25328),
            .in2(N__25000),
            .in3(N__24979),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_14_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__25304),
            .in2(N__24976),
            .in3(N__24955),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_15_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__25280),
            .in2(N__25333),
            .in3(N__25312),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_16_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__25256),
            .in2(N__25309),
            .in3(N__25288),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_17_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__25232),
            .in2(N__25285),
            .in3(N__25264),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_18_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__25211),
            .in2(N__25261),
            .in3(N__25240),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__52640),
            .ce(N__36477),
            .sr(N__52219));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_19_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__25187),
            .in2(N__25237),
            .in3(N__25216),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_19 ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_20_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__25213),
            .in2(N__25167),
            .in3(N__25195),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_21_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__25547),
            .in2(N__25192),
            .in3(N__25171),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_22_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__25523),
            .in2(N__25168),
            .in3(N__25147),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_23_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__25499),
            .in2(N__25552),
            .in3(N__25531),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_24_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__25475),
            .in2(N__25528),
            .in3(N__25507),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_25_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__25451),
            .in2(N__25504),
            .in3(N__25483),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_26_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(N__25427),
            .in2(N__25480),
            .in3(N__25459),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__52633),
            .ce(N__36476),
            .sr(N__52225));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_27_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__25391),
            .in2(N__25456),
            .in3(N__25435),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_27 ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__52627),
            .ce(N__36475),
            .sr(N__52234));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_28_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__25355),
            .in2(N__25432),
            .in3(N__25411),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__52627),
            .ce(N__36475),
            .sr(N__52234));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_29_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__25407),
            .in2(N__25396),
            .in3(N__25375),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__52627),
            .ce(N__36475),
            .sr(N__52234));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_30_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__25371),
            .in2(N__25360),
            .in3(N__25339),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_tr_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__52627),
            .ce(N__36475),
            .sr(N__52234));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_31_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25336),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52627),
            .ce(N__36475),
            .sr(N__52234));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_8_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_8_12_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_10_LC_8_12_0  (
            .in0(N__25611),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_12_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4FPBB_26_LC_8_12_1  (
            .in0(N__33772),
            .in1(N__25600),
            .in2(_gnd_net_),
            .in3(N__27094),
            .lcout(elapsed_time_ns_1_RNI4FPBB_0_26),
            .ltout(elapsed_time_ns_1_RNI4FPBB_0_26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_8_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_8_12_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_26_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25594),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_15_LC_8_12_3  (
            .in0(N__25590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_12_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNILK91B_9_LC_8_12_4  (
            .in0(N__25579),
            .in1(N__26941),
            .in2(_gnd_net_),
            .in3(N__33771),
            .lcout(elapsed_time_ns_1_RNILK91B_0_9),
            .ltout(elapsed_time_ns_1_RNILK91B_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_8_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_8_12_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_9_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25573),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_8_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_8_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_14_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25569),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_8_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_8_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_21_LC_8_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33796),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_13_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_inv_LC_8_13_0  (
            .in0(N__36691),
            .in1(N__25558),
            .in2(N__36742),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.measured_delay_tr_i_31 ),
            .ltout(),
            .carryin(bfn_8_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_13_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_0_c_RNIC7NP_LC_8_13_1  (
            .in0(N__27268),
            .in1(N__27264),
            .in2(N__51471),
            .in3(N__25639),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_1),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_13_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_1_c_RNIEBPP_LC_8_13_2  (
            .in0(N__27238),
            .in1(N__27231),
            .in2(N__51495),
            .in3(N__25636),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_2),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_13_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_2_c_RNIGFRP_LC_8_13_3  (
            .in0(N__27213),
            .in1(N__27214),
            .in2(N__51472),
            .in3(N__25633),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_3),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_13_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_3_c_RNIIJTP_LC_8_13_4  (
            .in0(N__27181),
            .in1(N__27177),
            .in2(N__51496),
            .in3(N__25630),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_4),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_13_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_4_c_RNIKNVP_LC_8_13_5  (
            .in0(N__27157),
            .in1(N__27156),
            .in2(N__51473),
            .in3(N__25627),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_5),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_13_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_5_c_RNIMR1Q_LC_8_13_6  (
            .in0(N__27513),
            .in1(N__27517),
            .in2(N__51497),
            .in3(N__25624),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_6),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_13_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_6_c_RNIOV3Q_LC_8_13_7  (
            .in0(N__27490),
            .in1(N__27489),
            .in2(N__51474),
            .in3(N__25621),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_7),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_14_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_7_c_RNI19MO_LC_8_14_0  (
            .in0(N__27475),
            .in1(N__27474),
            .in2(N__51469),
            .in3(N__25618),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_8),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_14_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_8_c_RNI3DOO_LC_8_14_1  (
            .in0(N__27445),
            .in1(N__27441),
            .in2(N__51466),
            .in3(N__25615),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_9),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_14_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_9_c_RNI5HQO_LC_8_14_2  (
            .in0(N__27421),
            .in1(N__27417),
            .in2(N__51470),
            .in3(N__25729),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_10),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_14_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_10_c_RNIELQC_LC_8_14_3  (
            .in0(N__27390),
            .in1(N__27391),
            .in2(N__51463),
            .in3(N__25726),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_11),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_14_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_11_c_RNIGPSC_LC_8_14_4  (
            .in0(N__27364),
            .in1(N__27360),
            .in2(N__51467),
            .in3(N__25723),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_12),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_14_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_12_c_RNIITUC_LC_8_14_5  (
            .in0(N__27330),
            .in1(N__27331),
            .in2(N__51464),
            .in3(N__25720),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_13),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_14_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_13_c_RNIK11D_LC_8_14_6  (
            .in0(N__27724),
            .in1(N__27723),
            .in2(N__51468),
            .in3(N__25717),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_14),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_14_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_14_c_RNIM53D_LC_8_14_7  (
            .in0(N__27700),
            .in1(N__27699),
            .in2(N__51465),
            .in3(N__25714),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_15),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_15_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_15_c_RNIO95D_LC_8_15_0  (
            .in0(N__27676),
            .in1(N__27675),
            .in2(N__51298),
            .in3(N__25687),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_16),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_15_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_16_c_RNIQD7D_LC_8_15_1  (
            .in0(N__27655),
            .in1(N__27651),
            .in2(N__51373),
            .in3(N__25663),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_17),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_15_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_17_c_RNIJ02E_LC_8_15_2  (
            .in0(N__27625),
            .in1(N__27621),
            .in2(N__51299),
            .in3(N__25642),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_18),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_15_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_18_c_RNIL44E_LC_8_15_3  (
            .in0(N__27600),
            .in1(N__27601),
            .in2(N__51374),
            .in3(N__25774),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_19),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_15_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_19_c_RNIN86E_LC_8_15_4  (
            .in0(N__27565),
            .in1(N__27561),
            .in2(N__51300),
            .in3(N__25771),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_20),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_15_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_20_c_RNIGR0F_LC_8_15_5  (
            .in0(N__27543),
            .in1(N__27544),
            .in2(N__51375),
            .in3(N__25750),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_21),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_15_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_21_c_RNIIV2F_LC_8_15_6  (
            .in0(N__27910),
            .in1(N__27909),
            .in2(N__51301),
            .in3(N__25747),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_22),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_15_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_22_c_RNIK35F_LC_8_15_7  (
            .in0(N__27886),
            .in1(N__27885),
            .in2(N__51376),
            .in3(N__25744),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_23),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_16_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_23_c_RNIM77F_LC_8_16_0  (
            .in0(N__27859),
            .in1(N__27858),
            .in2(N__51294),
            .in3(N__25741),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_24),
            .ltout(),
            .carryin(bfn_8_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_16_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_24_c_RNIOB9F_LC_8_16_1  (
            .in0(N__27838),
            .in1(N__27834),
            .in2(N__51296),
            .in3(N__25738),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_25),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_16_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_25_c_RNIQFBF_LC_8_16_2  (
            .in0(N__27802),
            .in1(N__27798),
            .in2(N__51295),
            .in3(N__25735),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_26),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_16_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_26_c_RNISJDF_LC_8_16_3  (
            .in0(N__27777),
            .in1(N__27778),
            .in2(N__51297),
            .in3(N__25732),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_27),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_LUT4_0_LC_8_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25915),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_8_17_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_8_17_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_0_LC_8_17_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_0_LC_8_17_0  (
            .in0(N__32503),
            .in1(N__25894),
            .in2(N__25912),
            .in3(N__25911),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_17_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_0 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_8_17_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_8_17_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_1_LC_8_17_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_1_LC_8_17_1  (
            .in0(N__32490),
            .in1(N__25882),
            .in2(_gnd_net_),
            .in3(N__25870),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_1 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_8_17_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_8_17_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_2_LC_8_17_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_2_LC_8_17_2  (
            .in0(N__32504),
            .in1(N__25867),
            .in2(_gnd_net_),
            .in3(N__25855),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_2 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_8_17_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_8_17_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_3_LC_8_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_3_LC_8_17_3  (
            .in0(N__32491),
            .in1(N__25852),
            .in2(_gnd_net_),
            .in3(N__25840),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_3 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_8_17_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_8_17_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_4_LC_8_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_4_LC_8_17_4  (
            .in0(N__32505),
            .in1(N__25837),
            .in2(_gnd_net_),
            .in3(N__25825),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_4 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_8_17_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_8_17_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_5_LC_8_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_5_LC_8_17_5  (
            .in0(N__32492),
            .in1(N__25822),
            .in2(_gnd_net_),
            .in3(N__25810),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_5 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_8_17_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_8_17_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_6_LC_8_17_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_6_LC_8_17_6  (
            .in0(N__32506),
            .in1(N__25807),
            .in2(_gnd_net_),
            .in3(N__25795),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_6 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_8_17_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_8_17_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_7_LC_8_17_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_7_LC_8_17_7  (
            .in0(N__32493),
            .in1(N__26035),
            .in2(_gnd_net_),
            .in3(N__26023),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_7 ),
            .clk(N__52584),
            .ce(N__26269),
            .sr(N__52251));
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_8_18_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_8_18_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_8_LC_8_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_8_LC_8_18_0  (
            .in0(N__32489),
            .in1(N__26020),
            .in2(_gnd_net_),
            .in3(N__26008),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_8 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_8_18_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_8_18_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_9_LC_8_18_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_9_LC_8_18_1  (
            .in0(N__32499),
            .in1(N__26005),
            .in2(_gnd_net_),
            .in3(N__25993),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_9 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_8_18_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_8_18_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_10_LC_8_18_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_10_LC_8_18_2  (
            .in0(N__32486),
            .in1(N__25990),
            .in2(_gnd_net_),
            .in3(N__25978),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_10 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_8_18_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_8_18_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_11_LC_8_18_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_11_LC_8_18_3  (
            .in0(N__32500),
            .in1(N__25975),
            .in2(_gnd_net_),
            .in3(N__25963),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_11 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_8_18_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_8_18_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_12_LC_8_18_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_12_LC_8_18_4  (
            .in0(N__32487),
            .in1(N__25960),
            .in2(_gnd_net_),
            .in3(N__25948),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_12 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_8_18_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_8_18_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_13_LC_8_18_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_13_LC_8_18_5  (
            .in0(N__32501),
            .in1(N__25945),
            .in2(_gnd_net_),
            .in3(N__25933),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_13 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_8_18_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_8_18_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_14_LC_8_18_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_14_LC_8_18_6  (
            .in0(N__32488),
            .in1(N__25930),
            .in2(_gnd_net_),
            .in3(N__25918),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_14 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_8_18_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_8_18_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_15_LC_8_18_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_15_LC_8_18_7  (
            .in0(N__32502),
            .in1(N__26254),
            .in2(_gnd_net_),
            .in3(N__26242),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_15 ),
            .clk(N__52578),
            .ce(N__26270),
            .sr(N__52256));
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_8_19_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_8_19_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_16_LC_8_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_16_LC_8_19_0  (
            .in0(N__32478),
            .in1(N__26232),
            .in2(_gnd_net_),
            .in3(N__26218),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_8_19_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_16 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_8_19_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_8_19_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_17_LC_8_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_17_LC_8_19_1  (
            .in0(N__32482),
            .in1(N__26202),
            .in2(_gnd_net_),
            .in3(N__26188),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_17 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_8_19_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_8_19_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_18_LC_8_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_18_LC_8_19_2  (
            .in0(N__32479),
            .in1(N__26178),
            .in2(_gnd_net_),
            .in3(N__26164),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_18 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_8_19_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_8_19_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_19_LC_8_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_19_LC_8_19_3  (
            .in0(N__32483),
            .in1(N__26154),
            .in2(_gnd_net_),
            .in3(N__26140),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_19 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_8_19_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_8_19_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_20_LC_8_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_20_LC_8_19_4  (
            .in0(N__32480),
            .in1(N__26129),
            .in2(_gnd_net_),
            .in3(N__26113),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_20 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_8_19_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_8_19_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_21_LC_8_19_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_21_LC_8_19_5  (
            .in0(N__32484),
            .in1(N__26108),
            .in2(_gnd_net_),
            .in3(N__26092),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_21 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_8_19_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_8_19_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_22_LC_8_19_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_22_LC_8_19_6  (
            .in0(N__32481),
            .in1(N__26076),
            .in2(_gnd_net_),
            .in3(N__26062),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_22 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_8_19_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_8_19_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_23_LC_8_19_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_23_LC_8_19_7  (
            .in0(N__32485),
            .in1(N__26052),
            .in2(_gnd_net_),
            .in3(N__26038),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_23 ),
            .clk(N__52573),
            .ce(N__26271),
            .sr(N__52260));
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_8_20_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_8_20_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_24_LC_8_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_24_LC_8_20_0  (
            .in0(N__32494),
            .in1(N__26451),
            .in2(_gnd_net_),
            .in3(N__26437),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_8_20_0_),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_24 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_8_20_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_8_20_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_25_LC_8_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_25_LC_8_20_1  (
            .in0(N__32507),
            .in1(N__26421),
            .in2(_gnd_net_),
            .in3(N__26407),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_25 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_8_20_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_8_20_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_26_LC_8_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_26_LC_8_20_2  (
            .in0(N__32495),
            .in1(N__26391),
            .in2(_gnd_net_),
            .in3(N__26377),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_26 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_8_20_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_8_20_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_27_LC_8_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_27_LC_8_20_3  (
            .in0(N__32508),
            .in1(N__26367),
            .in2(_gnd_net_),
            .in3(N__26353),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_27 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_8_20_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_8_20_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_28_LC_8_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_28_LC_8_20_4  (
            .in0(N__32496),
            .in1(N__26350),
            .in2(_gnd_net_),
            .in3(N__26332),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_28 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_8_20_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_8_20_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_29_LC_8_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_29_LC_8_20_5  (
            .in0(N__32509),
            .in1(N__26329),
            .in2(_gnd_net_),
            .in3(N__26314),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_29 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_8_20_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_8_20_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_30_LC_8_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_30_LC_8_20_6  (
            .in0(N__32497),
            .in1(N__26311),
            .in2(_gnd_net_),
            .in3(N__26296),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_tr.counter_cry_29 ),
            .carryout(\phase_controller_inst2.stoper_tr.counter_cry_30 ),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_8_20_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_8_20_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.counter_31_LC_8_20_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_tr.counter_31_LC_8_20_7  (
            .in0(N__26290),
            .in1(N__32498),
            .in2(_gnd_net_),
            .in3(N__26293),
            .lcout(\phase_controller_inst2.stoper_tr.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52567),
            .ce(N__26272),
            .sr(N__52262));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_8_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_8_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_8_21_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_15_LC_8_21_0  (
            .in0(_gnd_net_),
            .in1(N__26701),
            .in2(N__26683),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_16 ),
            .ltout(),
            .carryin(bfn_8_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_8_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_8_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15_c_RNIDMOM_LC_8_21_1  (
            .in0(_gnd_net_),
            .in1(N__26662),
            .in2(N__26647),
            .in3(N__26629),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_8_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_8_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_8_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16_c_RNIEOPM_LC_8_21_2  (
            .in0(_gnd_net_),
            .in1(N__26626),
            .in2(N__26611),
            .in3(N__26584),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_8_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_8_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17_c_RNIFQQM_LC_8_21_3  (
            .in0(_gnd_net_),
            .in1(N__26581),
            .in2(N__26563),
            .in3(N__26545),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_8_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_8_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_8_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18_c_RNIGSRM_LC_8_21_4  (
            .in0(_gnd_net_),
            .in1(N__26542),
            .in2(N__30764),
            .in3(N__26524),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_8_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_8_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19_c_RNIHUSM_LC_8_21_5  (
            .in0(_gnd_net_),
            .in1(N__26521),
            .in2(N__30766),
            .in3(N__26503),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_8_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_8_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20_c_RNI9FMN_LC_8_21_6  (
            .in0(_gnd_net_),
            .in1(N__26500),
            .in2(N__30765),
            .in3(N__26482),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_8_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_8_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_8_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21_c_RNIAHNN_LC_8_21_7  (
            .in0(_gnd_net_),
            .in1(N__26479),
            .in2(N__30767),
            .in3(N__26461),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_8_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_8_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_22_c_RNIBJON_LC_8_22_0  (
            .in0(_gnd_net_),
            .in1(N__26848),
            .in2(N__30768),
            .in3(N__26830),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_24 ),
            .ltout(),
            .carryin(bfn_8_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_8_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_8_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_8_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23_c_RNICLPN_LC_8_22_1  (
            .in0(_gnd_net_),
            .in1(N__26827),
            .in2(N__30772),
            .in3(N__26812),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_8_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_8_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_8_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24_c_RNIDNQN_LC_8_22_2  (
            .in0(_gnd_net_),
            .in1(N__26809),
            .in2(N__30769),
            .in3(N__26791),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_8_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_8_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_8_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25_c_RNIEPRN_LC_8_22_3  (
            .in0(_gnd_net_),
            .in1(N__26788),
            .in2(N__30773),
            .in3(N__26770),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_8_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_8_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_8_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26_c_RNIFRSN_LC_8_22_4  (
            .in0(_gnd_net_),
            .in1(N__26767),
            .in2(N__30770),
            .in3(N__26749),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_8_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_8_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27_c_RNIGTTN_LC_8_22_5  (
            .in0(_gnd_net_),
            .in1(N__26746),
            .in2(N__30774),
            .in3(N__26728),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_8_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_8_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_8_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28_c_RNIHVUN_LC_8_22_6  (
            .in0(_gnd_net_),
            .in1(N__26725),
            .in2(N__30771),
            .in3(N__26707),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_8_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_8_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_8_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_LUT4_0_LC_8_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26704),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNIO57L_LC_9_5_7  (
            .in0(N__52290),
            .in1(N__34440),
            .in2(_gnd_net_),
            .in3(N__34395),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_LC_9_7_1  (
            .in0(N__34436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52646),
            .ce(),
            .sr(N__52195));
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_3 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_LC_9_7_3  (
            .in0(N__26870),
            .in1(N__34351),
            .in2(N__30955),
            .in3(N__29467),
            .lcout(\phase_controller_inst2.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52646),
            .ce(),
            .sr(N__52195));
    defparam \phase_controller_inst2.start_timer_tr_LC_9_7_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_LC_9_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_tr_LC_9_7_4 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \phase_controller_inst2.start_timer_tr_LC_9_7_4  (
            .in0(N__29441),
            .in1(N__26854),
            .in2(N__29409),
            .in3(N__29268),
            .lcout(\phase_controller_inst2.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52646),
            .ce(),
            .sr(N__52195));
    defparam \phase_controller_inst2.state_1_LC_9_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_1_LC_9_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_1_LC_9_7_5 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \phase_controller_inst2.state_1_LC_9_7_5  (
            .in0(N__26895),
            .in1(N__29442),
            .in2(N__26878),
            .in3(N__29404),
            .lcout(\phase_controller_inst2.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52646),
            .ce(),
            .sr(N__52195));
    defparam \phase_controller_inst2.start_timer_hc_LC_9_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_timer_hc_LC_9_7_6 .LUT_INIT=16'b1111001111100000;
    LogicCell40 \phase_controller_inst2.start_timer_hc_LC_9_7_6  (
            .in0(N__29375),
            .in1(N__26894),
            .in2(N__29331),
            .in3(N__34435),
            .lcout(\phase_controller_inst2.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52646),
            .ce(),
            .sr(N__52195));
    defparam \phase_controller_inst2.state_2_LC_9_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_2_LC_9_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_2_LC_9_7_7 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst2.state_2_LC_9_7_7  (
            .in0(N__26896),
            .in1(N__29376),
            .in2(N__26877),
            .in3(N__29327),
            .lcout(\phase_controller_inst2.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52646),
            .ce(),
            .sr(N__52195));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_9_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_9_8_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNIEPKV_LC_9_8_0  (
            .in0(N__52292),
            .in1(N__29267),
            .in2(_gnd_net_),
            .in3(N__32537),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_8_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.start_timer_tr_RNO_0_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__26893),
            .in2(_gnd_net_),
            .in3(N__26869),
            .lcout(\phase_controller_inst2.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_9_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_9_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIL9L7_5_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__29697),
            .in2(_gnd_net_),
            .in3(N__27054),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_9_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_9_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_18_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26967),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_8_4 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_RNIODFQ_LC_9_8_4  (
            .in0(N__29466),
            .in1(_gnd_net_),
            .in2(N__34396),
            .in3(N__34430),
            .lcout(\phase_controller_inst2.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU6AF_1_LC_9_8_6  (
            .in0(N__29850),
            .in1(N__29715),
            .in2(N__29812),
            .in3(N__29767),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6HPBB_28_LC_9_9_0  (
            .in0(N__33767),
            .in1(N__27744),
            .in2(_gnd_net_),
            .in3(N__27079),
            .lcout(elapsed_time_ns_1_RNI6HPBB_0_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV8OBB_12_LC_9_9_1  (
            .in0(N__33709),
            .in1(N__27136),
            .in2(_gnd_net_),
            .in3(N__26923),
            .lcout(elapsed_time_ns_1_RNIV8OBB_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_9_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_9_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNII56P1_15_LC_9_9_2  (
            .in0(N__26976),
            .in1(N__27126),
            .in2(N__26997),
            .in3(N__29535),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_9_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_9_9_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNISL457_15_LC_9_9_3  (
            .in0(N__27292),
            .in1(N__27004),
            .in2(N__26980),
            .in3(N__27064),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI5FOBB_18_LC_9_9_4  (
            .in0(N__26977),
            .in1(N__33710),
            .in2(_gnd_net_),
            .in3(N__26968),
            .lcout(elapsed_time_ns_1_RNI5FOBB_0_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIJRME1_9_LC_9_9_5  (
            .in0(N__29511),
            .in1(N__26952),
            .in2(N__26940),
            .in3(N__26922),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_9_9_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_9_9_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI6O9B2_13_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__26910),
            .in2(N__26899),
            .in3(N__33843),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_9_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_9_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_12_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27135),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_9_10_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_9_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3DOBB_16_LC_9_10_0  (
            .in0(N__33693),
            .in1(N__27115),
            .in2(_gnd_net_),
            .in3(N__27127),
            .lcout(elapsed_time_ns_1_RNI3DOBB_0_16),
            .ltout(elapsed_time_ns_1_RNI3DOBB_0_16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_9_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_9_10_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_16_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27109),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_9_10_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_9_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIMDAP1_25_LC_9_10_2  (
            .in0(N__27105),
            .in1(N__27090),
            .in2(N__29988),
            .in3(N__27075),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_10_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIHG91B_5_LC_9_10_3  (
            .in0(N__27043),
            .in1(N__33691),
            .in2(_gnd_net_),
            .in3(N__27058),
            .lcout(elapsed_time_ns_1_RNIHG91B_0_5),
            .ltout(elapsed_time_ns_1_RNIHG91B_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_9_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_9_10_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_5_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27034),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_9_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_9_10_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0CQBB_31_LC_9_10_5  (
            .in0(N__29598),
            .in1(N__36690),
            .in2(_gnd_net_),
            .in3(N__33692),
            .lcout(elapsed_time_ns_1_RNI0CQBB_0_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_9_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_9_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNID5BP1_23_LC_9_10_6  (
            .in0(N__27030),
            .in1(N__30003),
            .in2(N__27019),
            .in3(N__33603),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_9_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_9_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7T8P1_19_LC_9_10_7  (
            .in0(N__29664),
            .in1(N__27303),
            .in2(N__29880),
            .in3(N__33807),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1_c_inv_LC_9_11_0  (
            .in0(N__29566),
            .in1(N__36677),
            .in2(N__27286),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_1 ),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_inv_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(N__27277),
            .in2(_gnd_net_),
            .in3(N__29751),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axb_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2_c_RNIPD1B_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__29728),
            .in2(_gnd_net_),
            .in3(N__27271),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2B_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(N__29959),
            .in2(_gnd_net_),
            .in3(N__27247),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3_c_RNIQF2BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3B_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__27244),
            .in2(_gnd_net_),
            .in3(N__27217),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4_c_RNIRH3BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4B_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(N__29677),
            .in2(_gnd_net_),
            .in3(N__27193),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5_c_RNISJ4BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5B_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(N__27190),
            .in2(_gnd_net_),
            .in3(N__27160),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6_c_RNITL5BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6B_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__29908),
            .in2(_gnd_net_),
            .in3(N__27139),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7_c_RNIUN6BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7B_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__27523),
            .in2(_gnd_net_),
            .in3(N__27499),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_8_c_RNIVP7BZ0 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8B_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__27496),
            .in2(_gnd_net_),
            .in3(N__27478),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9_c_RNI0S8BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83Q9_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__29491),
            .in2(_gnd_net_),
            .in3(N__27457),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10_c_RNI83QZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95R9_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__27454),
            .in2(_gnd_net_),
            .in3(N__27424),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11_c_RNI95RZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7S9_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__33823),
            .in2(_gnd_net_),
            .in3(N__27400),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12_c_RNIA7SZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9T9_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__27397),
            .in2(_gnd_net_),
            .in3(N__27373),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13_c_RNIB9TZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBU9_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__27370),
            .in2(_gnd_net_),
            .in3(N__27343),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14_c_RNICBUZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_12_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDV9_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__27340),
            .in2(_gnd_net_),
            .in3(N__27313),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15_c_RNIDDVZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0A_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__29551),
            .in2(_gnd_net_),
            .in3(N__27712),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_16_c_RNIEF0AZ0 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1A_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__27709),
            .in2(_gnd_net_),
            .in3(N__27688),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17_c_RNIFH1AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2A_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__27685),
            .in2(_gnd_net_),
            .in3(N__27658),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18_c_RNIGJ2AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3A_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__30148),
            .in2(_gnd_net_),
            .in3(N__27634),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19_c_RNIHL3AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TA_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__27631),
            .in2(_gnd_net_),
            .in3(N__27604),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20_c_RNI96TAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UA_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__29890),
            .in2(_gnd_net_),
            .in3(N__27580),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21_c_RNIA8UAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVA_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__27577),
            .in2(_gnd_net_),
            .in3(N__27547),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22_c_RNIBAVAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0B_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__29941),
            .in2(_gnd_net_),
            .in3(N__27526),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23_c_RNICC0BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_23 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1B_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__30130),
            .in2(_gnd_net_),
            .in3(N__27898),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_24_c_RNIDE1BZ0 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2B_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__27895),
            .in2(_gnd_net_),
            .in3(N__27874),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25_c_RNIEG2BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3B_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__27871),
            .in2(_gnd_net_),
            .in3(N__27841),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26_c_RNIFI3BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4B_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__27730),
            .in2(_gnd_net_),
            .in3(N__27817),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27_c_RNIGK4BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5B_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__27814),
            .in2(_gnd_net_),
            .in3(N__27781),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28_c_RNIHM5BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6B_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__33583),
            .in2(_gnd_net_),
            .in3(N__27760),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29_c_RNIIO6BZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_tr.un3_target_ticks_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_14_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_14_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_cry_27_c_RNIL68G_LC_9_14_6  (
            .in0(N__36692),
            .in1(N__27757),
            .in2(_gnd_net_),
            .in3(N__27748),
            .lcout(phase_controller_inst1_stoper_tr_target_ticks_1_i_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_9_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_9_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_28_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27745),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_axb_8_LC_9_15_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un3_threshold_axb_8_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_axb_8_LC_9_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \pwm_generator_inst.un3_threshold_axb_8_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__28249),
            .in2(N__28237),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_9_15_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_1_s_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__28195),
            .in2(N__28180),
            .in3(N__28144),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_1_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_0 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_9_15_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_2_s_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__28141),
            .in2(N__28123),
            .in3(N__28087),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_2_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_1 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_9_15_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_3_s_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__28084),
            .in2(N__28066),
            .in3(N__28036),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_3_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_2 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_9_15_4 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_4_s_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__28388),
            .in2(N__28033),
            .in3(N__28003),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_4_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_3 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_9_15_5 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_9_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_5_s_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__28000),
            .in2(N__28409),
            .in3(N__27973),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_5_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_4 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_9_15_6 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_9_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_6_s_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__27970),
            .in2(N__28411),
            .in3(N__27943),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_6_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_5 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_9_15_7 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_9_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_7_s_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(N__27940),
            .in2(N__28410),
            .in3(N__28516),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_7_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_6 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_9_16_0 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_9_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_8_s_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__28513),
            .in2(N__28412),
            .in3(N__28483),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_8_sZ0 ),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_9_16_1 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_9_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_9_s_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__28401),
            .in2(N__28480),
            .in3(N__28450),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_9_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_8 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_9_16_2 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_9_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_10_s_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__28447),
            .in2(N__28413),
            .in3(N__28417),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_10_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_9 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_9_16_3 .C_ON=1'b1;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_9_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_s_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__28405),
            .in2(N__28330),
            .in3(N__28297),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_sZ0 ),
            .ltout(),
            .carryin(\pwm_generator_inst.un2_threshold_add_1_cry_10 ),
            .carryout(\pwm_generator_inst.un2_threshold_add_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_9_16_4 .C_ON=1'b0;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_LUT4_0_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28294),
            .lcout(\pwm_generator_inst.un2_threshold_add_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_17_0 .LUT_INIT=16'b0111010100010000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_24_LC_9_17_0  (
            .in0(N__31990),
            .in1(N__32014),
            .in2(N__28264),
            .in3(N__28669),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_24_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28275),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52579),
            .ce(N__36624),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_17_2 .LUT_INIT=16'b1111011101010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_24_LC_9_17_2  (
            .in0(N__31989),
            .in1(N__32013),
            .in2(N__28263),
            .in3(N__28668),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_25_LC_9_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28680),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52579),
            .ce(N__36624),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_17_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_26_LC_9_17_4  (
            .in0(N__28645),
            .in1(N__32368),
            .in2(N__31965),
            .in3(N__28621),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_26_LC_9_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28656),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52579),
            .ce(N__36624),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_17_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_26_LC_9_17_6  (
            .in0(N__28644),
            .in1(N__32367),
            .in2(N__31966),
            .in3(N__28620),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_9_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_27_LC_9_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_27_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28632),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52579),
            .ce(N__36624),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_1_LC_9_18_0 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_1_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(N__34693),
            .in2(N__28612),
            .in3(N__32878),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_1 ),
            .ltout(),
            .carryin(bfn_9_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .clk(N__52574),
            .ce(),
            .sr(N__52252));
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_2_LC_9_18_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_2_LC_9_18_1  (
            .in0(N__32877),
            .in1(N__34655),
            .in2(N__28588),
            .in3(N__28567),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .clk(N__52574),
            .ce(),
            .sr(N__52252));
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_3_LC_9_18_2 .LUT_INIT=16'b1101011101111101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_3_LC_9_18_2  (
            .in0(N__32880),
            .in1(N__34628),
            .in2(N__28564),
            .in3(N__28543),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .clk(N__52574),
            .ce(),
            .sr(N__52252));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_4_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(N__35089),
            .in2(N__28540),
            .in3(N__28519),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_5_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(N__35052),
            .in2(N__28876),
            .in3(N__28852),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_6_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(N__34998),
            .in2(N__28849),
            .in3(N__28828),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_7_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(N__34945),
            .in2(N__28825),
            .in3(N__28804),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_8_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(N__34909),
            .in2(N__28801),
            .in3(N__28783),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_9_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__28780),
            .in2(N__34860),
            .in3(N__28759),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_9 ),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_10_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__34822),
            .in2(N__28756),
            .in3(N__28738),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_11_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__34770),
            .in2(N__28735),
            .in3(N__28714),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_12_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__35424),
            .in2(N__28711),
            .in3(N__28687),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_13_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(N__35362),
            .in2(N__29014),
            .in3(N__28990),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_14_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__35299),
            .in2(N__28987),
            .in3(N__28963),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_15_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(N__35265),
            .in2(N__28960),
            .in3(N__28939),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_16_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__35202),
            .in2(N__28936),
            .in3(N__28921),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_17_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__28918),
            .in2(N__37619),
            .in3(N__28909),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_17 ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_18_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__28906),
            .in2(N__35157),
            .in3(N__28900),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_19_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__37667),
            .in2(N__28897),
            .in3(N__28888),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_20_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(N__28885),
            .in2(N__37704),
            .in3(N__28879),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_21_LC_9_20_4  (
            .in0(_gnd_net_),
            .in1(N__35685),
            .in2(N__29131),
            .in3(N__29119),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_22_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__29116),
            .in2(N__37580),
            .in3(N__29110),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_23_LC_9_20_6  (
            .in0(_gnd_net_),
            .in1(N__35652),
            .in2(N__29107),
            .in3(N__29098),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_24_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__35612),
            .in2(N__29095),
            .in3(N__29080),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_25_LC_9_21_0  (
            .in0(_gnd_net_),
            .in1(N__35577),
            .in2(N__29077),
            .in3(N__29068),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_25 ),
            .ltout(),
            .carryin(bfn_9_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_26_LC_9_21_1  (
            .in0(_gnd_net_),
            .in1(N__35547),
            .in2(N__29065),
            .in3(N__29056),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_27_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__35504),
            .in2(N__29053),
            .in3(N__29044),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_28_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__35462),
            .in2(N__29041),
            .in3(N__29029),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_29_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__35932),
            .in2(N__29026),
            .in3(N__29017),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNO_0_30_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__35898),
            .in2(N__29209),
            .in3(N__29200),
            .lcout(\current_shift_inst.PI_CTRL.integrator_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.un1_integrator_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.un1_integrator_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_9_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_er_31_LC_9_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_er_31_LC_9_21_6  (
            .in0(N__35829),
            .in1(N__29197),
            .in2(N__30670),
            .in3(N__29191),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52557),
            .ce(N__32924),
            .sr(N__52263));
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_27_LC_9_22_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_27_LC_9_22_0  (
            .in0(N__35817),
            .in1(N__32917),
            .in2(_gnd_net_),
            .in3(N__29188),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52553),
            .ce(),
            .sr(N__52264));
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_9_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_28_LC_9_22_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_28_LC_9_22_1  (
            .in0(N__32916),
            .in1(N__35820),
            .in2(_gnd_net_),
            .in3(N__29182),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52553),
            .ce(),
            .sr(N__52264));
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_9_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_29_LC_9_22_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_29_LC_9_22_2  (
            .in0(N__35818),
            .in1(N__32918),
            .in2(_gnd_net_),
            .in3(N__29176),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52553),
            .ce(),
            .sr(N__52264));
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_13_LC_9_22_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_13_LC_9_22_7  (
            .in0(N__32915),
            .in1(N__35819),
            .in2(_gnd_net_),
            .in3(N__29170),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52553),
            .ce(),
            .sr(N__52264));
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_9_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_9_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_15_LC_9_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_15_LC_9_23_1  (
            .in0(N__32925),
            .in1(N__35856),
            .in2(_gnd_net_),
            .in3(N__29161),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52548),
            .ce(),
            .sr(N__52267));
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_12_LC_9_23_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_12_LC_9_23_6  (
            .in0(N__35855),
            .in1(N__29152),
            .in2(_gnd_net_),
            .in3(N__32926),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52548),
            .ce(),
            .sr(N__52267));
    defparam \phase_controller_inst2.S1_LC_9_24_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.S1_LC_9_24_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S1_LC_9_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S1_LC_9_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29335),
            .lcout(s3_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52545),
            .ce(),
            .sr(N__52270));
    defparam \phase_controller_inst2.S2_LC_9_26_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.S2_LC_9_26_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.S2_LC_9_26_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.S2_LC_9_26_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29419),
            .lcout(s4_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52540),
            .ce(),
            .sr(N__52271));
    defparam \phase_controller_inst2.stoper_hc.running_LC_10_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.running_LC_10_6_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.running_LC_10_6_0 .LUT_INIT=16'b1100010011101110;
    LogicCell40 \phase_controller_inst2.stoper_hc.running_LC_10_6_0  (
            .in0(N__34434),
            .in1(N__29465),
            .in2(N__30954),
            .in3(N__34386),
            .lcout(\phase_controller_inst2.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52641),
            .ce(),
            .sr(N__52178));
    defparam \phase_controller_inst2.state_0_LC_10_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_0_LC_10_6_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_0_LC_10_6_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst2.state_0_LC_10_6_3  (
            .in0(N__29298),
            .in1(N__29446),
            .in2(N__29353),
            .in3(N__29405),
            .lcout(\phase_controller_inst2.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52641),
            .ce(),
            .sr(N__52178));
    defparam \phase_controller_inst2.state_RNO_0_3_LC_10_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.state_RNO_0_3_LC_10_7_0 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \phase_controller_inst2.state_RNO_0_3_LC_10_7_0  (
            .in0(N__29380),
            .in1(N__29323),
            .in2(N__29299),
            .in3(N__29349),
            .lcout(),
            .ltout(\phase_controller_inst2.state_ns_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.state_3_LC_10_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_3_LC_10_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.state_3_LC_10_7_1 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \phase_controller_inst2.state_3_LC_10_7_1  (
            .in0(N__34008),
            .in1(N__34063),
            .in2(N__29338),
            .in3(N__34084),
            .lcout(\phase_controller_inst2.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52635),
            .ce(),
            .sr(N__52187));
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_10_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_10_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_RNO_0_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__29265),
            .in2(_gnd_net_),
            .in3(N__32545),
            .lcout(),
            .ltout(\phase_controller_inst2.stoper_tr.un4_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_10_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_10_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.time_passed_LC_10_7_3 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \phase_controller_inst2.stoper_tr.time_passed_LC_10_7_3  (
            .in0(N__29653),
            .in1(N__29297),
            .in2(N__29302),
            .in3(N__29238),
            .lcout(\phase_controller_inst2.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52635),
            .ce(),
            .sr(N__52187));
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_10_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_10_7_6 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_RNI96ON_LC_10_7_6  (
            .in0(N__29651),
            .in1(N__29264),
            .in2(_gnd_net_),
            .in3(N__32544),
            .lcout(\phase_controller_inst2.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.running_LC_10_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.running_LC_10_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_tr.running_LC_10_7_7 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst2.stoper_tr.running_LC_10_7_7  (
            .in0(N__29266),
            .in1(N__29652),
            .in2(N__32555),
            .in3(N__29239),
            .lcout(\phase_controller_inst2.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52635),
            .ce(),
            .sr(N__52187));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_10_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_25_LC_10_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_25_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41143),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52629),
            .ce(N__41915),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_9_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_9_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNICUKU_7_LC_10_9_0  (
            .in0(N__29934),
            .in1(N__29638),
            .in2(N__29632),
            .in3(N__29608),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3lto30_i_a2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_9_1 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI7SETA_31_LC_10_9_1  (
            .in0(N__29602),
            .in1(N__29584),
            .in2(N__29578),
            .in3(N__29575),
            .lcout(\delay_measurement_inst.delay_tr_timer.delay_tr3 ),
            .ltout(\delay_measurement_inst.delay_tr_timer.delay_tr3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_10_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_10_9_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIDC91B_1_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__29808),
            .in2(N__29569),
            .in3(N__29565),
            .lcout(elapsed_time_ns_1_RNIDC91B_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_17_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29523),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI4EOBB_17_LC_10_9_4  (
            .in0(N__29524),
            .in1(_gnd_net_),
            .in2(N__33727),
            .in3(N__29539),
            .lcout(elapsed_time_ns_1_RNI4EOBB_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_9_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU7OBB_11_LC_10_9_5  (
            .in0(N__29500),
            .in1(N__29515),
            .in2(_gnd_net_),
            .in3(N__33682),
            .lcout(elapsed_time_ns_1_RNIU7OBB_0_11),
            .ltout(elapsed_time_ns_1_RNIU7OBB_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_9_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_11_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29494),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_10_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_10_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIFE91B_3_LC_10_9_7  (
            .in0(N__29740),
            .in1(N__29857),
            .in2(_gnd_net_),
            .in3(N__33681),
            .lcout(elapsed_time_ns_1_RNIFE91B_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_10_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_10_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_1_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__29839),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52613),
            .ce(N__36462),
            .sr(N__52206));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_10_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_2_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29794),
            .lcout(\delay_measurement_inst.delay_tr_timer.elapsed_time_tr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52613),
            .ce(N__36462),
            .sr(N__52206));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_10_10_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_10_10_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIED91B_2_LC_10_10_4  (
            .in0(N__29752),
            .in1(N__33694),
            .in2(_gnd_net_),
            .in3(N__29766),
            .lcout(elapsed_time_ns_1_RNIED91B_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_10_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_10_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_3_LC_10_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29739),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_10_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_10_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIGF91B_4_LC_10_10_7  (
            .in0(N__33695),
            .in1(N__29971),
            .in2(_gnd_net_),
            .in3(N__29722),
            .lcout(elapsed_time_ns_1_RNIGF91B_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIIH91B_6_LC_10_11_0  (
            .in0(N__29704),
            .in1(N__29686),
            .in2(_gnd_net_),
            .in3(N__33723),
            .lcout(elapsed_time_ns_1_RNIIH91B_0_6),
            .ltout(elapsed_time_ns_1_RNIIH91B_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_11_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_6_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29680),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0BPBB_22_LC_10_11_2  (
            .in0(N__29902),
            .in1(N__29671),
            .in2(_gnd_net_),
            .in3(N__33724),
            .lcout(elapsed_time_ns_1_RNI0BPBB_0_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI2DPBB_24_LC_10_11_3  (
            .in0(N__33725),
            .in1(N__29953),
            .in2(_gnd_net_),
            .in3(N__30010),
            .lcout(elapsed_time_ns_1_RNI2DPBB_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_11_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI3EPBB_25_LC_10_11_4  (
            .in0(N__30142),
            .in1(N__33726),
            .in2(_gnd_net_),
            .in3(N__29992),
            .lcout(elapsed_time_ns_1_RNI3EPBB_0_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_4_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29970),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_12_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_12_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_24_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29952),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_12_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIKJ91B_8_LC_10_12_1  (
            .in0(N__29935),
            .in1(N__29917),
            .in2(_gnd_net_),
            .in3(N__33728),
            .lcout(elapsed_time_ns_1_RNIKJ91B_0_8),
            .ltout(elapsed_time_ns_1_RNIKJ91B_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_12_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_8_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29911),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_10_12_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_10_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_22_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29901),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIU8PBB_20_LC_10_12_5  (
            .in0(N__29863),
            .in1(N__29884),
            .in2(_gnd_net_),
            .in3(N__33729),
            .lcout(elapsed_time_ns_1_RNIU8PBB_0_20),
            .ltout(elapsed_time_ns_1_RNIU8PBB_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_12_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_20_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30151),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_25_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30141),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_10_13_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_10_13_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_1_LC_10_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_1_LC_10_13_0  (
            .in0(N__30121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_10_13_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_6_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_6_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30106),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_10_13_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_5_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_5_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30091),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_10_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_13_LC_10_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_13_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30076),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_10_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_7_LC_10_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_7_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30058),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_10_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_4_LC_10_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_4_LC_10_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30043),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_10_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_2_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_2_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30024),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_10_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_3_LC_10_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_3_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30265),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52590),
            .ce(N__36617),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_10_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_10_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_0_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__36649),
            .in2(N__30250),
            .in3(N__31425),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_0 ),
            .ltout(),
            .carryin(bfn_10_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_10_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_1_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(N__30241),
            .in2(N__30235),
            .in3(N__31785),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_10_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_10_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_2_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__30217),
            .in2(N__30226),
            .in3(N__31770),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_10_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_10_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_3_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(N__30211),
            .in2(N__30205),
            .in3(N__31755),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_10_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_10_14_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_4_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__30196),
            .in2(N__30190),
            .in3(N__31740),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_10_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_10_14_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_5_LC_10_14_5  (
            .in0(N__31726),
            .in1(N__30181),
            .in2(N__30175),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_10_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_10_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_6_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(N__30166),
            .in2(N__30160),
            .in3(N__31707),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_10_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_10_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_7_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__30358),
            .in2(N__30352),
            .in3(N__31693),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_10_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_10_15_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_8_LC_10_15_0  (
            .in0(N__31674),
            .in1(N__30340),
            .in2(N__34156),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_8 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_10_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_10_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_9_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__34123),
            .in2(N__30334),
            .in3(N__31659),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_10_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_10_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_10_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__30325),
            .in2(N__34096),
            .in3(N__31936),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_10_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_10_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_11_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__34183),
            .in2(N__30319),
            .in3(N__31914),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_10_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_10_15_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_12_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__34243),
            .in2(N__30310),
            .in3(N__31899),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_10_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_10_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_13_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__30301),
            .in2(N__30292),
            .in3(N__31884),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_10_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_10_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_14_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__34270),
            .in2(N__30283),
            .in3(N__31869),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_10_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_10_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_inv_15_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__34213),
            .in2(N__30274),
            .in3(N__31854),
            .lcout(\phase_controller_inst1.stoper_tr.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_10_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_10_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_16_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__30454),
            .in2(N__30439),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_10_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_10_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_18_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__30421),
            .in2(N__30406),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_10_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_10_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_10_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_20_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__32080),
            .in2(N__32173),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_10_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_10_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_10_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_22_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__32692),
            .in2(N__32770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_10_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_10_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_10_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_24_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(N__30388),
            .in2(N__30382),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_10_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_10_16_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_10_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_26_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__30373),
            .in2(N__30367),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_10_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_10_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_28_LC_10_16_6  (
            .in0(_gnd_net_),
            .in1(N__34591),
            .in2(N__34528),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_10_16_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_10_16_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_10_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_30_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__34456),
            .in2(N__34516),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.un6_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_10_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_LUT4_0_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30502),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_17_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNI207E_LC_10_17_3  (
            .in0(N__36817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_10_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_10_17_4 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_RNI6D081_LC_10_17_4  (
            .in0(N__34315),
            .in1(N__36781),
            .in2(_gnd_net_),
            .in3(N__36816),
            .lcout(\phase_controller_inst1.stoper_tr.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_10_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_10_17_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNI5GRG_30_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(N__36815),
            .in2(_gnd_net_),
            .in3(N__34326),
            .lcout(\phase_controller_inst1.stoper_tr.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_4_LC_10_18_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_4_LC_10_18_0  (
            .in0(N__35863),
            .in1(N__30478),
            .in2(_gnd_net_),
            .in3(N__32898),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52563),
            .ce(),
            .sr(N__52245));
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_8_LC_10_18_2 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_8_LC_10_18_2  (
            .in0(N__35864),
            .in1(N__30472),
            .in2(_gnd_net_),
            .in3(N__32899),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52563),
            .ce(),
            .sr(N__52245));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_18_5 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI5DRS2_3_LC_10_18_5  (
            .in0(N__30550),
            .in1(N__35094),
            .in2(N__34920),
            .in3(N__34629),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_10_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_10_18_6 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNID5COE_18_LC_10_18_6  (
            .in0(N__33040),
            .in1(N__30526),
            .in2(N__30466),
            .in3(N__32962),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0 ),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_10_LC_10_18_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_10_LC_10_18_7  (
            .in0(N__30463),
            .in1(_gnd_net_),
            .in2(N__30457),
            .in3(N__35865),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52563),
            .ce(),
            .sr(N__52245));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_10_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_10_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIF12L1_5_LC_10_19_0  (
            .in0(N__34950),
            .in1(N__34997),
            .in2(N__35051),
            .in3(N__34859),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_6_LC_10_19_2 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_6_LC_10_19_2  (
            .in0(N__30544),
            .in1(N__35860),
            .in2(_gnd_net_),
            .in3(N__32881),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52559),
            .ce(),
            .sr(N__52247));
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_10_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_10_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_7_LC_10_19_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_7_LC_10_19_3  (
            .in0(N__35859),
            .in1(N__32879),
            .in2(_gnd_net_),
            .in3(N__30538),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52559),
            .ce(),
            .sr(N__52247));
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_9_LC_10_19_4 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_9_LC_10_19_4  (
            .in0(N__30532),
            .in1(N__35861),
            .in2(_gnd_net_),
            .in3(N__32882),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52559),
            .ce(),
            .sr(N__52247));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_10_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_10_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI95V81_18_LC_10_19_5  (
            .in0(N__35858),
            .in1(N__35150),
            .in2(_gnd_net_),
            .in3(N__32932),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_10_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_10_19_6 .LUT_INIT=16'b0000000001010111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIUF1L1_1_LC_10_19_6  (
            .in0(N__34627),
            .in1(N__34656),
            .in2(N__34701),
            .in3(N__35090),
            .lcout(\current_shift_inst.PI_CTRL.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_10_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_10_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_LC_10_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__34697),
            .in2(_gnd_net_),
            .in3(N__34729),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52559),
            .ce(),
            .sr(N__52247));
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_14_LC_10_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_14_LC_10_20_0  (
            .in0(N__35822),
            .in1(N__30520),
            .in2(_gnd_net_),
            .in3(N__32905),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_18_LC_10_20_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_18_LC_10_20_1  (
            .in0(N__32902),
            .in1(N__35826),
            .in2(_gnd_net_),
            .in3(N__30514),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_10_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_10_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_16_LC_10_20_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_16_LC_10_20_3  (
            .in0(N__32900),
            .in1(N__35825),
            .in2(_gnd_net_),
            .in3(N__30508),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_10_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_10_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_5_LC_10_20_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_5_LC_10_20_4  (
            .in0(N__35824),
            .in1(N__30607),
            .in2(_gnd_net_),
            .in3(N__32906),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_10_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_10_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_17_LC_10_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_17_LC_10_20_5  (
            .in0(N__32901),
            .in1(N__30598),
            .in2(_gnd_net_),
            .in3(N__35828),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_10_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_10_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_23_LC_10_20_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_23_LC_10_20_6  (
            .in0(N__35823),
            .in1(N__32904),
            .in2(_gnd_net_),
            .in3(N__30592),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_10_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_10_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_22_LC_10_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_22_LC_10_20_7  (
            .in0(N__32903),
            .in1(N__35827),
            .in2(_gnd_net_),
            .in3(N__30586),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52555),
            .ce(),
            .sr(N__52253));
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_10_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_24_LC_10_21_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_24_LC_10_21_1  (
            .in0(N__32907),
            .in1(N__35814),
            .in2(_gnd_net_),
            .in3(N__30580),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52550),
            .ce(),
            .sr(N__52257));
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_10_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_10_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_20_LC_10_21_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_20_LC_10_21_2  (
            .in0(N__35811),
            .in1(N__32910),
            .in2(_gnd_net_),
            .in3(N__30574),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52550),
            .ce(),
            .sr(N__52257));
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_30_LC_10_21_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_30_LC_10_21_3  (
            .in0(N__32909),
            .in1(N__35816),
            .in2(_gnd_net_),
            .in3(N__30568),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52550),
            .ce(),
            .sr(N__52257));
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_10_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_10_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_25_LC_10_21_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_25_LC_10_21_4  (
            .in0(N__35813),
            .in1(N__32912),
            .in2(_gnd_net_),
            .in3(N__30562),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52550),
            .ce(),
            .sr(N__52257));
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_26_LC_10_21_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_26_LC_10_21_5  (
            .in0(N__32908),
            .in1(N__35815),
            .in2(_gnd_net_),
            .in3(N__30556),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52550),
            .ce(),
            .sr(N__52257));
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_10_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_21_LC_10_21_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_21_LC_10_21_6  (
            .in0(N__35812),
            .in1(N__32911),
            .in2(_gnd_net_),
            .in3(N__30808),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52550),
            .ce(),
            .sr(N__52257));
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_11_LC_10_22_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_11_LC_10_22_2  (
            .in0(N__35821),
            .in1(N__30802),
            .in2(_gnd_net_),
            .in3(N__32914),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52547),
            .ce(),
            .sr(N__52261));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_10_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_10_23_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_0_12_LC_10_23_0  (
            .in0(N__35461),
            .in1(N__35503),
            .in2(N__35413),
            .in3(N__35897),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_23_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_er_RNO_0_31_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__30793),
            .in2(_gnd_net_),
            .in3(N__30775),
            .lcout(\current_shift_inst.PI_CTRL.integrator_1_0_add_1_axb_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_5_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_0_LC_11_5_0  (
            .in0(N__31102),
            .in1(N__41965),
            .in2(N__30658),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_0 ),
            .ltout(),
            .carryin(bfn_11_5_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_1_LC_11_5_1  (
            .in0(_gnd_net_),
            .in1(N__33298),
            .in2(N__30649),
            .in3(N__31087),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_2_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__33004),
            .in2(N__30640),
            .in3(N__31066),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_3_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__32998),
            .in2(N__30628),
            .in3(N__31048),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_4_LC_11_5_4  (
            .in0(_gnd_net_),
            .in1(N__33088),
            .in2(N__30619),
            .in3(N__31024),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_5_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_5_LC_11_5_5  (
            .in0(N__31006),
            .in1(N__32992),
            .in2(N__30877),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_5_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_6_LC_11_5_6  (
            .in0(N__30988),
            .in1(N__33094),
            .in2(N__30868),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_5_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_7_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__33100),
            .in2(N__30859),
            .in3(N__31300),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_8_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(N__30850),
            .in2(N__32986),
            .in3(N__31279),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_8 ),
            .ltout(),
            .carryin(bfn_11_6_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_9_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__33010),
            .in2(N__30844),
            .in3(N__31258),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_10_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(N__33292),
            .in2(N__30835),
            .in3(N__31240),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_11_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__30826),
            .in2(N__33076),
            .in3(N__31222),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_12_LC_11_6_4  (
            .in0(_gnd_net_),
            .in1(N__33055),
            .in2(N__30820),
            .in3(N__31204),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_13_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__33082),
            .in2(N__30907),
            .in3(N__31186),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_14_LC_11_6_6  (
            .in0(N__31165),
            .in1(N__33067),
            .in2(N__30898),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_inv_15_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__33061),
            .in2(N__30886),
            .in3(N__31147),
            .lcout(\phase_controller_inst2.stoper_hc.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_16_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__33286),
            .in2(N__33223),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_18_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__30961),
            .in2(N__33130),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_20_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__30967),
            .in2(N__31126),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_22_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__30913),
            .in2(N__30922),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_24_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__33307),
            .in2(N__33505),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_26_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__33493),
            .in2(N__33430),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_28_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__33406),
            .in2(N__33364),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_30_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__33925),
            .in2(N__33865),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.un6_running_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30970),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_8_1 .LUT_INIT=16'b0010101100001010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_20_LC_11_8_1  (
            .in0(N__33349),
            .in1(N__31402),
            .in2(N__31381),
            .in3(N__33109),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_11_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_11_8_2 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_18_LC_11_8_2  (
            .in0(N__33189),
            .in1(N__33205),
            .in2(N__33166),
            .in3(N__33121),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_8_3 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNIH2SA_30_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__34397),
            .in2(_gnd_net_),
            .in3(N__30938),
            .lcout(\phase_controller_inst2.stoper_hc.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_8_4 .LUT_INIT=16'b0000101010001110;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_22_LC_11_8_4  (
            .in0(N__33331),
            .in1(N__33340),
            .in2(N__31327),
            .in3(N__31353),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_11_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_11_8_5 .LUT_INIT=16'b1000110011101111;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_22_LC_11_8_5  (
            .in0(N__33339),
            .in1(N__33330),
            .in2(N__31354),
            .in3(N__31326),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_11_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_11_8_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst2.stoper_hc.start_latched_RNI8HE4_LC_11_8_6  (
            .in0(N__34398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_11_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_11_8_7 .LUT_INIT=16'b1010111100101011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_20_LC_11_8_7  (
            .in0(N__33348),
            .in1(N__31401),
            .in2(N__31380),
            .in3(N__33108),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_11_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_11_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_0_LC_11_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_0_LC_11_9_0  (
            .in0(N__31575),
            .in1(N__31101),
            .in2(N__31117),
            .in3(N__31116),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_0 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_11_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_11_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_1_LC_11_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_1_LC_11_9_1  (
            .in0(N__31613),
            .in1(N__31083),
            .in2(_gnd_net_),
            .in3(N__31069),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_0 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_1 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_11_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_11_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_2_LC_11_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_2_LC_11_9_2  (
            .in0(N__31576),
            .in1(N__31065),
            .in2(_gnd_net_),
            .in3(N__31051),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_1 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_2 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_11_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_11_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_3_LC_11_9_3 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_3_LC_11_9_3  (
            .in0(N__31614),
            .in1(_gnd_net_),
            .in2(N__31047),
            .in3(N__31027),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_2 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_3 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_11_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_11_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_4_LC_11_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_4_LC_11_9_4  (
            .in0(N__31577),
            .in1(N__31023),
            .in2(_gnd_net_),
            .in3(N__31009),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_3 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_4 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_11_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_11_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_5_LC_11_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_5_LC_11_9_5  (
            .in0(N__31615),
            .in1(N__31005),
            .in2(_gnd_net_),
            .in3(N__30991),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_4 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_5 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_11_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_11_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_6_LC_11_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_6_LC_11_9_6  (
            .in0(N__31578),
            .in1(N__30987),
            .in2(_gnd_net_),
            .in3(N__30973),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_5 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_6 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_11_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_7_LC_11_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_7_LC_11_9_7  (
            .in0(N__31616),
            .in1(N__31296),
            .in2(_gnd_net_),
            .in3(N__31282),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_6 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_7 ),
            .clk(N__52614),
            .ce(N__31490),
            .sr(N__52191));
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_11_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_11_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_8_LC_11_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_8_LC_11_10_0  (
            .in0(N__31600),
            .in1(N__31275),
            .in2(_gnd_net_),
            .in3(N__31261),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_8 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_11_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_9_LC_11_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_9_LC_11_10_1  (
            .in0(N__31612),
            .in1(N__31257),
            .in2(_gnd_net_),
            .in3(N__31243),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_8 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_9 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_11_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_11_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_10_LC_11_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_10_LC_11_10_2  (
            .in0(N__31597),
            .in1(N__31239),
            .in2(_gnd_net_),
            .in3(N__31225),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_9 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_10 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_11_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_11_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_11_LC_11_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_11_LC_11_10_3  (
            .in0(N__31609),
            .in1(N__31221),
            .in2(_gnd_net_),
            .in3(N__31207),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_10 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_11 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_11_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_11_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_12_LC_11_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_12_LC_11_10_4  (
            .in0(N__31598),
            .in1(N__31203),
            .in2(_gnd_net_),
            .in3(N__31189),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_11 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_12 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_11_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_11_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_13_LC_11_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_13_LC_11_10_5  (
            .in0(N__31610),
            .in1(N__31182),
            .in2(_gnd_net_),
            .in3(N__31168),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_12 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_13 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_11_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_11_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_14_LC_11_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_14_LC_11_10_6  (
            .in0(N__31599),
            .in1(N__31164),
            .in2(_gnd_net_),
            .in3(N__31150),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_13 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_14 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_11_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_11_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_15_LC_11_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_15_LC_11_10_7  (
            .in0(N__31611),
            .in1(N__31143),
            .in2(_gnd_net_),
            .in3(N__31129),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_14 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_15 ),
            .clk(N__52605),
            .ce(N__31489),
            .sr(N__52196));
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_11_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_11_11_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_16_LC_11_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_16_LC_11_11_0  (
            .in0(N__31601),
            .in1(N__33237),
            .in2(_gnd_net_),
            .in3(N__31414),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_16 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_11_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_11_11_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_17_LC_11_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_17_LC_11_11_1  (
            .in0(N__31605),
            .in1(N__33264),
            .in2(_gnd_net_),
            .in3(N__31411),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_16 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_17 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_11_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_11_11_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_18_LC_11_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_18_LC_11_11_2  (
            .in0(N__31602),
            .in1(N__33152),
            .in2(_gnd_net_),
            .in3(N__31408),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_17 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_18 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_11_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_19_LC_11_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_19_LC_11_11_3  (
            .in0(N__31606),
            .in1(N__33185),
            .in2(_gnd_net_),
            .in3(N__31405),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_18 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_19 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_11_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_11_11_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_20_LC_11_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_20_LC_11_11_4  (
            .in0(N__31603),
            .in1(N__31400),
            .in2(_gnd_net_),
            .in3(N__31384),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_19 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_20 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_11_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_11_11_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_21_LC_11_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_21_LC_11_11_5  (
            .in0(N__31607),
            .in1(N__31373),
            .in2(_gnd_net_),
            .in3(N__31357),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_20 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_21 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_11_11_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_11_11_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_22_LC_11_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_22_LC_11_11_6  (
            .in0(N__31604),
            .in1(N__31344),
            .in2(_gnd_net_),
            .in3(N__31330),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_21 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_22 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_11_11_7 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_11_11_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_23_LC_11_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_23_LC_11_11_7  (
            .in0(N__31608),
            .in1(N__31317),
            .in2(_gnd_net_),
            .in3(N__31303),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_22 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_23 ),
            .clk(N__52598),
            .ce(N__31491),
            .sr(N__52207));
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_11_12_0 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_11_12_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_24_LC_11_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_24_LC_11_12_0  (
            .in0(N__31617),
            .in1(N__33521),
            .in2(_gnd_net_),
            .in3(N__31645),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_24 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_11_12_1 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_11_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_25_LC_11_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_25_LC_11_12_1  (
            .in0(N__31622),
            .in1(N__33560),
            .in2(_gnd_net_),
            .in3(N__31642),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_24 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_25 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_11_12_2 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_11_12_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_26_LC_11_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_26_LC_11_12_2  (
            .in0(N__31618),
            .in1(N__33444),
            .in2(_gnd_net_),
            .in3(N__31639),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_25 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_26 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_11_12_3 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_11_12_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_27_LC_11_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_27_LC_11_12_3  (
            .in0(N__31623),
            .in1(N__33473),
            .in2(_gnd_net_),
            .in3(N__31636),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_26 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_27 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_11_12_4 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_28_LC_11_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_28_LC_11_12_4  (
            .in0(N__31619),
            .in1(N__33379),
            .in2(_gnd_net_),
            .in3(N__31633),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_27 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_28 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_11_12_5 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_11_12_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_29_LC_11_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_29_LC_11_12_5  (
            .in0(N__31624),
            .in1(N__33394),
            .in2(_gnd_net_),
            .in3(N__31630),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_28 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_29 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_11_12_6 .C_ON=1'b1;
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_11_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_30_LC_11_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_30_LC_11_12_6  (
            .in0(N__31620),
            .in1(N__33883),
            .in2(_gnd_net_),
            .in3(N__31627),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst2.stoper_hc.counter_cry_29 ),
            .carryout(\phase_controller_inst2.stoper_hc.counter_cry_30 ),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_11_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_11_12_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.stoper_hc.counter_31_LC_11_12_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst2.stoper_hc.counter_31_LC_11_12_7  (
            .in0(N__33898),
            .in1(N__31621),
            .in2(_gnd_net_),
            .in3(N__31495),
            .lcout(\phase_controller_inst2.stoper_hc.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52591),
            .ce(N__31492),
            .sr(N__52213));
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_11_13_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_11_13_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_0_LC_11_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_0_LC_11_13_0  (
            .in0(N__32320),
            .in1(N__31426),
            .in2(N__31447),
            .in3(N__31446),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_0 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_11_13_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_11_13_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_1_LC_11_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_1_LC_11_13_1  (
            .in0(N__32324),
            .in1(N__31786),
            .in2(_gnd_net_),
            .in3(N__31774),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_1 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_11_13_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_11_13_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_2_LC_11_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_2_LC_11_13_2  (
            .in0(N__32321),
            .in1(N__31771),
            .in2(_gnd_net_),
            .in3(N__31759),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_2 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_11_13_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_11_13_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_3_LC_11_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_3_LC_11_13_3  (
            .in0(N__32325),
            .in1(N__31756),
            .in2(_gnd_net_),
            .in3(N__31744),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_3 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_11_13_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_11_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_4_LC_11_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_4_LC_11_13_4  (
            .in0(N__32322),
            .in1(N__31741),
            .in2(_gnd_net_),
            .in3(N__31729),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_4 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_11_13_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_11_13_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_5_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_5_LC_11_13_5  (
            .in0(N__32326),
            .in1(N__31725),
            .in2(_gnd_net_),
            .in3(N__31711),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_5 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_11_13_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_11_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_6_LC_11_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_6_LC_11_13_6  (
            .in0(N__32323),
            .in1(N__31708),
            .in2(_gnd_net_),
            .in3(N__31696),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_6 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_11_13_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_11_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_7_LC_11_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_7_LC_11_13_7  (
            .in0(N__32327),
            .in1(N__31692),
            .in2(_gnd_net_),
            .in3(N__31678),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_7 ),
            .clk(N__52586),
            .ce(N__32191),
            .sr(N__52220));
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_11_14_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_11_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_8_LC_11_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_8_LC_11_14_0  (
            .in0(N__32331),
            .in1(N__31675),
            .in2(_gnd_net_),
            .in3(N__31663),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_8 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_11_14_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_11_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_9_LC_11_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_9_LC_11_14_1  (
            .in0(N__32335),
            .in1(N__31660),
            .in2(_gnd_net_),
            .in3(N__31648),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_9 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_11_14_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_11_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_10_LC_11_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_10_LC_11_14_2  (
            .in0(N__32328),
            .in1(N__31932),
            .in2(_gnd_net_),
            .in3(N__31918),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_10 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_11_14_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_11_LC_11_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_11_LC_11_14_3  (
            .in0(N__32332),
            .in1(N__31915),
            .in2(_gnd_net_),
            .in3(N__31903),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_11 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_11_14_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_11_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_12_LC_11_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_12_LC_11_14_4  (
            .in0(N__32329),
            .in1(N__31900),
            .in2(_gnd_net_),
            .in3(N__31888),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_12 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_11_14_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_11_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_13_LC_11_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_13_LC_11_14_5  (
            .in0(N__32333),
            .in1(N__31885),
            .in2(_gnd_net_),
            .in3(N__31873),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_13 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_11_14_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_11_14_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_14_LC_11_14_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_14_LC_11_14_6  (
            .in0(N__32330),
            .in1(N__31870),
            .in2(_gnd_net_),
            .in3(N__31858),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_14 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_11_14_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_11_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_15_LC_11_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_15_LC_11_14_7  (
            .in0(N__32334),
            .in1(N__31855),
            .in2(_gnd_net_),
            .in3(N__31843),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_15 ),
            .clk(N__52581),
            .ce(N__32190),
            .sr(N__52229));
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_11_15_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_11_15_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_16_LC_11_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_16_LC_11_15_0  (
            .in0(N__32312),
            .in1(N__31827),
            .in2(_gnd_net_),
            .in3(N__31813),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_16 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_11_15_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_17_LC_11_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_17_LC_11_15_1  (
            .in0(N__32316),
            .in1(N__31803),
            .in2(_gnd_net_),
            .in3(N__31789),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_17 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_11_15_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_18_LC_11_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_18_LC_11_15_2  (
            .in0(N__32313),
            .in1(N__32066),
            .in2(_gnd_net_),
            .in3(N__32050),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_18 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_11_15_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_19_LC_11_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_19_LC_11_15_3  (
            .in0(N__32317),
            .in1(N__32045),
            .in2(_gnd_net_),
            .in3(N__32029),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_19 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_11_15_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_20_LC_11_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_20_LC_11_15_4  (
            .in0(N__32314),
            .in1(N__32096),
            .in2(_gnd_net_),
            .in3(N__32026),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_20 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_11_15_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_11_15_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_21_LC_11_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_21_LC_11_15_5  (
            .in0(N__32318),
            .in1(N__32114),
            .in2(_gnd_net_),
            .in3(N__32023),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_21 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_11_15_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_11_15_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_22_LC_11_15_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_22_LC_11_15_6  (
            .in0(N__32315),
            .in1(N__32708),
            .in2(_gnd_net_),
            .in3(N__32020),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_22 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_11_15_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_11_15_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_23_LC_11_15_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_23_LC_11_15_7  (
            .in0(N__32319),
            .in1(N__32741),
            .in2(_gnd_net_),
            .in3(N__32017),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_23 ),
            .clk(N__52576),
            .ce(N__32189),
            .sr(N__52235));
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_11_16_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_11_16_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_24_LC_11_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_24_LC_11_16_0  (
            .in0(N__32268),
            .in1(N__32007),
            .in2(_gnd_net_),
            .in3(N__31993),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_11_16_0_),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_24 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_11_16_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_11_16_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_25_LC_11_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_25_LC_11_16_1  (
            .in0(N__32272),
            .in1(N__31983),
            .in2(_gnd_net_),
            .in3(N__31969),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_25 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_11_16_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_11_16_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_26_LC_11_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_26_LC_11_16_2  (
            .in0(N__32269),
            .in1(N__31953),
            .in2(_gnd_net_),
            .in3(N__31939),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_26 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_11_16_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_11_16_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_27_LC_11_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_27_LC_11_16_3  (
            .in0(N__32273),
            .in1(N__32361),
            .in2(_gnd_net_),
            .in3(N__32347),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_27 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_11_16_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_28_LC_11_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_28_LC_11_16_4  (
            .in0(N__32270),
            .in1(N__34543),
            .in2(_gnd_net_),
            .in3(N__32344),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_28 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_11_16_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_11_16_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_29_LC_11_16_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_29_LC_11_16_5  (
            .in0(N__32274),
            .in1(N__34558),
            .in2(_gnd_net_),
            .in3(N__32341),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_29 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_11_16_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_11_16_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_30_LC_11_16_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_30_LC_11_16_6  (
            .in0(N__32271),
            .in1(N__34504),
            .in2(_gnd_net_),
            .in3(N__32338),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_tr.counter_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_tr.counter_cry_30 ),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_11_16_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_11_16_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.counter_31_LC_11_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.counter_31_LC_11_16_7  (
            .in0(N__32275),
            .in1(N__34471),
            .in2(_gnd_net_),
            .in3(N__32194),
            .lcout(\phase_controller_inst1.stoper_tr.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52569),
            .ce(N__32188),
            .sr(N__52238));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_17_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_17_0 .LUT_INIT=16'b0000110010001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_20_LC_11_17_0  (
            .in0(N__32143),
            .in1(N__32134),
            .in2(N__32122),
            .in3(N__32098),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_11_17_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_20_LC_11_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_20_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32161),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52564),
            .ce(N__36616),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_17_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_17_2 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_20_LC_11_17_2  (
            .in0(N__32142),
            .in1(N__32133),
            .in2(N__32121),
            .in3(N__32097),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_17_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_17_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_22_LC_11_17_4  (
            .in0(N__32743),
            .in1(N__32725),
            .in2(N__32716),
            .in3(N__32668),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_11_17_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_22_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_22_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32761),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52564),
            .ce(N__36616),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_17_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_17_6 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_22_LC_11_17_6  (
            .in0(N__32742),
            .in1(N__32724),
            .in2(N__32715),
            .in3(N__32667),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_11_17_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_23_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_23_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32686),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52564),
            .ce(N__36616),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_11_18_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_tr.target_ticks_28_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_tr.target_ticks_28_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34582),
            .lcout(\phase_controller_inst2.stoper_tr.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52560),
            .ce(N__32638),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_11_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_inv_LC_11_18_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_inv_LC_11_18_7  (
            .in0(N__42556),
            .in1(N__51142),
            .in2(_gnd_net_),
            .in3(N__40039),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_11_19_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_11_19_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst2.stoper_tr.start_latched_RNI3ORE_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32560),
            .lcout(\phase_controller_inst2.stoper_tr.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_11_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_11_19_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_0_11_LC_11_19_2  (
            .in0(N__35200),
            .in1(N__35363),
            .in2(N__35307),
            .in3(N__34766),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_11_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_11_19_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIQGDL2_18_LC_11_19_3  (
            .in0(N__35857),
            .in1(N__35149),
            .in2(N__32371),
            .in3(N__32938),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_11_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_11_19_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNILDEP7_12_LC_11_19_4  (
            .in0(N__32977),
            .in1(N__33031),
            .in2(N__32965),
            .in3(N__32947),
            .lcout(\current_shift_inst.PI_CTRL.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_11_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_11_19_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIPEP71_5_LC_11_19_6  (
            .in0(N__34946),
            .in1(N__34990),
            .in2(_gnd_net_),
            .in3(N__35041),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_o2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_11_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_11_19_7 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI23CN3_8_LC_11_19_7  (
            .in0(N__34855),
            .in1(N__34913),
            .in2(N__32956),
            .in3(N__32953),
            .lcout(\current_shift_inst.PI_CTRL.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_11_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_11_20_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIAA5B_23_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__35942),
            .in2(_gnd_net_),
            .in3(N__35644),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_11_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_11_20_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNINJGC1_10_LC_11_20_1  (
            .in0(N__35260),
            .in1(N__34823),
            .in2(N__32941),
            .in3(N__37543),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_11_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_11_20_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_17_LC_11_20_3  (
            .in0(N__37696),
            .in1(N__37657),
            .in2(N__37579),
            .in3(N__37609),
            .lcout(\current_shift_inst.PI_CTRL.N_46_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_11_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_11_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.integrator_19_LC_11_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_19_LC_11_20_7  (
            .in0(N__32913),
            .in1(N__35866),
            .in2(_gnd_net_),
            .in3(N__32779),
            .lcout(\current_shift_inst.PI_CTRL.integratorZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52551),
            .ce(),
            .sr(N__52248));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_11_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_11_21_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_21_LC_11_21_0  (
            .in0(N__35683),
            .in1(N__35536),
            .in2(N__35616),
            .in3(N__35576),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_10_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_11_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_11_21_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNI626M_11_LC_11_21_1  (
            .in0(N__35300),
            .in1(N__34759),
            .in2(N__35370),
            .in3(N__35201),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_8_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_11_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_11_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIA53P2_10_LC_11_21_2  (
            .in0(N__33022),
            .in1(N__33049),
            .in2(N__33043),
            .in3(N__33016),
            .lcout(\current_shift_inst.PI_CTRL.N_46_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_11_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_11_21_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICCAM_0_21_LC_11_21_3  (
            .in0(N__35575),
            .in1(N__35611),
            .in2(N__35546),
            .in3(N__35684),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_11_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_11_21_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIDDAM_12_LC_11_21_5  (
            .in0(N__35472),
            .in1(N__35514),
            .in2(N__35423),
            .in3(N__35893),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_11_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_11_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_11_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNIB98M_10_LC_11_21_6  (
            .in0(N__34824),
            .in1(N__35261),
            .in2(N__35953),
            .in3(N__35645),
            .lcout(\current_shift_inst.PI_CTRL.integrator_4_iv_0_a3_0_20_9_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_9_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40792),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_5_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_2_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40633),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_3_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40609),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_5_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_5_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40885),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_8_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40813),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_7_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40837),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_6_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40861),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_4_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40909),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52634),
            .ce(N__41932),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_13_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41083),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_11_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40744),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_14_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41059),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_15_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41563),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_12_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_18_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_18_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40978),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_12_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40720),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_6_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_1_LC_12_6_6  (
            .in0(N__40657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_10_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40768),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52628),
            .ce(N__41933),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_7_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_16_LC_12_7_0  (
            .in0(N__33280),
            .in1(N__33271),
            .in2(N__33250),
            .in3(N__33214),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_12_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_16_LC_12_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_16_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41032),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52622),
            .ce(N__41934),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_12_7_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_12_7_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_16_LC_12_7_2  (
            .in0(N__33279),
            .in1(N__33270),
            .in2(N__33249),
            .in3(N__33213),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_12_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_17_LC_12_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_17_LC_12_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41005),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52622),
            .ce(N__41934),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_12_7_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_12_7_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_18_LC_12_7_6  (
            .in0(N__33204),
            .in1(N__33190),
            .in2(N__33165),
            .in3(N__33120),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_12_7_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_19_LC_12_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_19_LC_12_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40956),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52622),
            .ce(N__41934),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_12_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_20_LC_12_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_20_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40930),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52612),
            .ce(N__41947),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_21_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41224),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52612),
            .ce(N__41947),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_12_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_22_LC_12_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_22_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41203),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52612),
            .ce(N__41947),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_12_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_12_8_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_23_LC_12_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_23_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41182),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52612),
            .ce(N__41947),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_9_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_9_0  (
            .in0(N__33320),
            .in1(N__36147),
            .in2(_gnd_net_),
            .in3(N__36165),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_12_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_28_LC_12_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_28_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42601),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52604),
            .ce(N__42032),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_12_9_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_12_9_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_28_LC_12_9_2  (
            .in0(N__33319),
            .in1(N__36146),
            .in2(_gnd_net_),
            .in3(N__36164),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_12_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_12_9_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_30_LC_12_9_3  (
            .in0(N__36104),
            .in1(N__36128),
            .in2(_gnd_net_),
            .in3(N__33321),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_9_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_9_4  (
            .in0(N__33322),
            .in1(N__36105),
            .in2(_gnd_net_),
            .in3(N__36129),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_12_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_12_10_0 .LUT_INIT=16'b0011000010110010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_24_LC_12_10_0  (
            .in0(N__33571),
            .in1(N__33562),
            .in2(N__33543),
            .in3(N__33523),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_12_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_24_LC_12_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_24_LC_12_10_1  (
            .in0(N__41161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52597),
            .ce(N__41948),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_12_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_12_10_2 .LUT_INIT=16'b1011001011110011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_24_LC_12_10_2  (
            .in0(N__33570),
            .in1(N__33561),
            .in2(N__33544),
            .in3(N__33522),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_12_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_12_10_4 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_26_LC_12_10_4  (
            .in0(N__33484),
            .in1(N__33475),
            .in2(N__33457),
            .in3(N__33415),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_12_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_26_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_26_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41122),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52597),
            .ce(N__41948),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_12_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_12_10_6 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_26_LC_12_10_6  (
            .in0(N__33483),
            .in1(N__33474),
            .in2(N__33456),
            .in3(N__33414),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_12_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_27_LC_12_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_27_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41104),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52597),
            .ce(N__41948),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_11_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_28_LC_12_11_0  (
            .in0(N__33911),
            .in1(N__33393),
            .in2(_gnd_net_),
            .in3(N__33378),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_12_11_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_12_11_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_28_LC_12_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_28_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42597),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52589),
            .ce(N__41953),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_12_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_12_11_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_28_LC_12_11_2  (
            .in0(N__33910),
            .in1(N__33392),
            .in2(_gnd_net_),
            .in3(N__33377),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_11_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_30_LC_12_11_3  (
            .in0(N__33896),
            .in1(N__33881),
            .in2(_gnd_net_),
            .in3(N__33912),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_1_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_11_4 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_11_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst2.stoper_hc.un6_running_cry_c_RNO_0_30_LC_12_11_4  (
            .in0(N__33913),
            .in1(N__33897),
            .in2(_gnd_net_),
            .in3(N__33882),
            .lcout(\phase_controller_inst2.stoper_hc.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_12_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIM3UN_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__47524),
            .in2(_gnd_net_),
            .in3(N__47501),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_165_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.running_LC_12_12_3 .LUT_INIT=16'b0101111101010000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_LC_12_12_3  (
            .in0(N__47502),
            .in1(_gnd_net_),
            .in2(N__47534),
            .in3(N__47580),
            .lcout(\delay_measurement_inst.delay_hc_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52585),
            .ce(),
            .sr(N__52208));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_12_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNI0AOBB_13_LC_12_12_5  (
            .in0(N__33768),
            .in1(N__33850),
            .in2(_gnd_net_),
            .in3(N__33832),
            .lcout(elapsed_time_ns_1_RNI0AOBB_0_13),
            .ltout(elapsed_time_ns_1_RNI0AOBB_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_12_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_12_12_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_13_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33826),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIV9PBB_21_LC_12_13_0  (
            .in0(N__33769),
            .in1(N__33792),
            .in2(_gnd_net_),
            .in3(N__33814),
            .lcout(elapsed_time_ns_1_RNIV9PBB_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_12_13_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_12_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.elapsed_time_ns_1_RNIVAQBB_30_LC_12_13_2  (
            .in0(N__33770),
            .in1(N__33592),
            .in2(_gnd_net_),
            .in3(N__33610),
            .lcout(elapsed_time_ns_1_RNIVAQBB_0_30),
            .ltout(elapsed_time_ns_1_RNIVAQBB_0_30_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_12_13_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_12_13_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_tr.un3_target_ticks_axb_30_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33586),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_tr.un3_target_ticks_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_flag_LC_12_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_flag_LC_12_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_flag_LC_12_13_4 .LUT_INIT=16'b1111100011111000;
    LogicCell40 \phase_controller_inst1.start_flag_LC_12_13_4  (
            .in0(N__34032),
            .in1(N__33989),
            .in2(N__33973),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52580),
            .ce(),
            .sr(N__52214));
    defparam \phase_controller_inst1.state_4_LC_12_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_4_LC_12_13_5 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst1.state_4_LC_12_13_5 .LUT_INIT=16'b1000100010101010;
    LogicCell40 \phase_controller_inst1.state_4_LC_12_13_5  (
            .in0(N__33990),
            .in1(N__33968),
            .in2(_gnd_net_),
            .in3(N__34033),
            .lcout(\phase_controller_inst1.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52580),
            .ce(),
            .sr(N__52214));
    defparam \phase_controller_inst2.start_flag_LC_12_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.start_flag_LC_12_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst2.start_flag_LC_12_13_6 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \phase_controller_inst2.start_flag_LC_12_13_6  (
            .in0(N__34034),
            .in1(_gnd_net_),
            .in2(N__34062),
            .in3(N__34076),
            .lcout(\phase_controller_inst2.start_flagZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52580),
            .ce(),
            .sr(N__52214));
    defparam \phase_controller_inst2.state_4_LC_12_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst2.state_4_LC_12_13_7 .SEQ_MODE=4'b1011;
    defparam \phase_controller_inst2.state_4_LC_12_13_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst2.state_4_LC_12_13_7  (
            .in0(N__34077),
            .in1(N__34055),
            .in2(_gnd_net_),
            .in3(N__34035),
            .lcout(\phase_controller_inst2.stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52580),
            .ce(),
            .sr(N__52214));
    defparam \phase_controller_inst1.state_RNO_0_3_LC_12_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.state_RNO_0_3_LC_12_14_0 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \phase_controller_inst1.state_RNO_0_3_LC_12_14_0  (
            .in0(N__36409),
            .in1(N__50328),
            .in2(N__33951),
            .in3(N__33933),
            .lcout(),
            .ltout(\phase_controller_inst1.state_ns_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_3_LC_12_14_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_3_LC_12_14_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_3_LC_12_14_1 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \phase_controller_inst1.state_3_LC_12_14_1  (
            .in0(N__34036),
            .in1(N__33991),
            .in2(N__33976),
            .in3(N__33972),
            .lcout(state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52575),
            .ce(),
            .sr(N__52221));
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_RNO_0_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__36771),
            .in2(_gnd_net_),
            .in3(N__36803),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_tr.un4_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_3 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \phase_controller_inst1.stoper_tr.time_passed_LC_12_14_3  (
            .in0(N__34310),
            .in1(N__33950),
            .in2(N__33955),
            .in3(N__34335),
            .lcout(\phase_controller_inst1.tr_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52575),
            .ce(),
            .sr(N__52221));
    defparam \phase_controller_inst1.state_0_LC_12_14_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_0_LC_12_14_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_0_LC_12_14_4 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \phase_controller_inst1.state_0_LC_12_14_4  (
            .in0(N__36333),
            .in1(N__38096),
            .in2(N__33952),
            .in3(N__33934),
            .lcout(\phase_controller_inst1.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52575),
            .ce(),
            .sr(N__52221));
    defparam \phase_controller_inst1.start_timer_tr_LC_12_14_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_LC_12_14_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_tr_LC_12_14_5 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_LC_12_14_5  (
            .in0(N__38095),
            .in1(N__36332),
            .in2(N__36780),
            .in3(N__36223),
            .lcout(\phase_controller_inst1.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52575),
            .ce(),
            .sr(N__52221));
    defparam \phase_controller_inst1.stoper_tr.running_LC_12_14_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.running_LC_12_14_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.running_LC_12_14_7 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst1.stoper_tr.running_LC_12_14_7  (
            .in0(N__36772),
            .in1(N__34311),
            .in2(N__36814),
            .in3(N__34336),
            .lcout(\phase_controller_inst1.stoper_tr.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52575),
            .ce(),
            .sr(N__52221));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_15_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_14_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34291),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_12_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34261),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_15_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34234),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_15_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_11_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34201),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_15_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_8_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34174),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_15_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_9_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34141),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_15_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_10_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34114),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52568),
            .ce(N__36593),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_12_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_12_16_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_28_LC_12_16_0  (
            .in0(N__34485),
            .in1(N__34557),
            .in2(_gnd_net_),
            .in3(N__34542),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_16_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_28_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34581),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52562),
            .ce(N__36595),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_12_16_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_12_16_2 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_28_LC_12_16_2  (
            .in0(N__34484),
            .in1(N__34556),
            .in2(_gnd_net_),
            .in3(N__34541),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_12_16_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_12_16_3 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_30_LC_12_16_3  (
            .in0(N__34469),
            .in1(N__34502),
            .in2(_gnd_net_),
            .in3(N__34483),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0Z0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_12_16_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_12_16_4 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \phase_controller_inst1.stoper_tr.un6_running_cry_c_RNO_0_30_LC_12_16_4  (
            .in0(N__34503),
            .in1(_gnd_net_),
            .in2(N__34489),
            .in3(N__34470),
            .lcout(\phase_controller_inst1.stoper_tr.un6_running_lt30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_12_16_6 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_12_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst2.stoper_hc.time_passed_RNO_0_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__34447),
            .in2(_gnd_net_),
            .in3(N__34399),
            .lcout(\phase_controller_inst2.stoper_hc.un4_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_12_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_12_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_13_LC_12_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_13_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37404),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52558),
            .ce(),
            .sr(N__52239));
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_2_LC_12_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36984),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52558),
            .ce(),
            .sr(N__52239));
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_12_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_12_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_1_LC_12_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_1_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37008),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52558),
            .ce(),
            .sr(N__52239));
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_12_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_12_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_4_LC_12_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_4_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37233),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52558),
            .ce(),
            .sr(N__52239));
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_12_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_12_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_10_LC_12_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_10_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37068),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52554),
            .ce(),
            .sr(N__52241));
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_12_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_12_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_5_LC_12_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_5_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37206),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52554),
            .ce(),
            .sr(N__52241));
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_12_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_6_LC_12_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_6_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37179),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52554),
            .ce(),
            .sr(N__52241));
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_12_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_12_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_9_LC_12_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_9_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37095),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52554),
            .ce(),
            .sr(N__52241));
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_12_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_12_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_12_LC_12_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_12_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37434),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52554),
            .ce(),
            .sr(N__52241));
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_3_LC_12_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_3_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36957),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52554),
            .ce(),
            .sr(N__52241));
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_12_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_12_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_14_LC_12_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_14_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37374),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_12_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_12_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_11_LC_12_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_11_LC_12_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37041),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_12_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_12_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_15_LC_12_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_15_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37350),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_12_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_12_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_16_LC_12_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_16_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37323),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_12_19_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_12_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_17_LC_12_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_17_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37296),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_19_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_7_LC_12_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_7_LC_12_19_5  (
            .in0(N__37152),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_12_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_12_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_19_LC_12_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_19_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37263),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_12_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_12_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_8_LC_12_19_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_8_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(N__37119),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52549),
            .ce(),
            .sr(N__52243));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_12_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_12_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_1_cry_1_c_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__34725),
            .in2(N__34708),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_12_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_2_LC_12_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_2_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__34675),
            .in2(N__34666),
            .in3(N__34639),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_12_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_3_LC_12_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_3_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(N__34636),
            .in2(N__34606),
            .in3(N__34594),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_12_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_4_LC_12_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_4_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__35110),
            .in2(N__35101),
            .in3(N__35068),
            .lcout(\current_shift_inst.PI_CTRL.un7_enablelto4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_12_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_5_LC_12_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_5_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(N__35065),
            .in2(N__35056),
            .in3(N__35014),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_12_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_12_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_6_LC_12_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_6_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(N__35011),
            .in2(N__35002),
            .in3(N__34966),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_12_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_12_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_7_LC_12_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_7_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(N__34963),
            .in2(N__34957),
            .in3(N__34924),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_12_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_12_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_8_LC_12_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_8_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(N__34921),
            .in2(N__34888),
            .in3(N__34879),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_8 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_7 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_8 ),
            .clk(N__52546),
            .ce(),
            .sr(N__52246));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_12_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_12_21_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_9_LC_12_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_9_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(N__34876),
            .in2(N__34867),
            .in3(N__34831),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_9 ),
            .ltout(),
            .carryin(bfn_12_21_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_12_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_12_21_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_10_LC_12_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_10_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__34828),
            .in2(N__34798),
            .in3(N__34786),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_12_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_12_21_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_11_LC_12_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_11_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(N__34783),
            .in2(N__34774),
            .in3(N__34732),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_12_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_12_21_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_12_LC_12_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_12_LC_12_21_3  (
            .in0(_gnd_net_),
            .in1(N__35434),
            .in2(N__35425),
            .in3(N__35383),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_12_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_12_21_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_13_LC_12_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_13_LC_12_21_4  (
            .in0(_gnd_net_),
            .in1(N__35380),
            .in2(N__35371),
            .in3(N__35326),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_12_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_12_21_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_14_LC_12_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_14_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(N__35323),
            .in2(N__35314),
            .in3(N__35278),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_12_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_12_21_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_15_LC_12_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_15_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__35275),
            .in2(N__35266),
            .in3(N__35224),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_12_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_12_21_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_16_LC_12_21_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_16_LC_12_21_7  (
            .in0(_gnd_net_),
            .in1(N__35221),
            .in2(N__35212),
            .in3(N__35179),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_16 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_15 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_16 ),
            .clk(N__52543),
            .ce(),
            .sr(N__52249));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_12_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_12_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_17_LC_12_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_17_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__35176),
            .in2(N__37632),
            .in3(N__35167),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_17 ),
            .ltout(),
            .carryin(bfn_12_22_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_12_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_12_22_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_18_LC_12_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_18_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(N__37510),
            .in2(N__35164),
            .in3(N__35128),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_12_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_19_LC_12_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_19_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(N__35125),
            .in2(N__37672),
            .in3(N__35113),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_12_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_12_22_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_20_LC_12_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_20_LC_12_22_3  (
            .in0(_gnd_net_),
            .in1(N__37918),
            .in2(N__37711),
            .in3(N__35698),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_12_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_12_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_21_LC_12_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_21_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__37888),
            .in2(N__35695),
            .in3(N__35665),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_12_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_12_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_22_LC_12_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_22_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(N__37585),
            .in2(N__37978),
            .in3(N__35662),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_12_22_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_12_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_23_LC_12_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_23_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(N__37945),
            .in2(N__35659),
            .in3(N__35626),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_12_22_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_12_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_24_LC_12_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_24_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(N__37477),
            .in2(N__35623),
            .in3(N__35590),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_24 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_23 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_24 ),
            .clk(N__52541),
            .ce(),
            .sr(N__52254));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_12_23_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_12_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_25_LC_12_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_25_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(N__38188),
            .in2(N__35587),
            .in3(N__35557),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_25 ),
            .ltout(),
            .carryin(bfn_12_23_0_),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_12_23_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_12_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_26_LC_12_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_26_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(N__37771),
            .in2(N__35554),
            .in3(N__35521),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_12_23_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_12_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_27_LC_12_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_27_LC_12_23_2  (
            .in0(_gnd_net_),
            .in1(N__37801),
            .in2(N__35518),
            .in3(N__35479),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_12_23_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_12_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_28_LC_12_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_28_LC_12_23_3  (
            .in0(_gnd_net_),
            .in1(N__38161),
            .in2(N__35476),
            .in3(N__35437),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_12_23_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_12_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_29_LC_12_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_29_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(N__37828),
            .in2(N__35952),
            .in3(N__35908),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_12_23_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_12_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_30_LC_12_23_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_30_LC_12_23_5  (
            .in0(_gnd_net_),
            .in1(N__37861),
            .in2(N__35905),
            .in3(N__35869),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.output_unclamped_1_cry_30 ),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_12_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_12_23_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_31_LC_12_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_31_LC_12_23_6  (
            .in0(N__35862),
            .in1(N__38215),
            .in2(_gnd_net_),
            .in3(N__35722),
            .lcout(\current_shift_inst.PI_CTRL.un8_enablelto31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52539),
            .ce(),
            .sr(N__52258));
    defparam GB_BUFFER_reset_c_g_THRU_LUT4_0_LC_12_30_1.C_ON=1'b0;
    defparam GB_BUFFER_reset_c_g_THRU_LUT4_0_LC_12_30_1.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_reset_c_g_THRU_LUT4_0_LC_12_30_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_reset_c_g_THRU_LUT4_0_LC_12_30_1 (
            .in0(N__52294),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_reset_c_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_13_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_16_LC_13_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_16_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41031),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52636),
            .ce(N__42037),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_13_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_17_LC_13_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_17_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41004),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52636),
            .ce(N__42037),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_13_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_13_6_4 .LUT_INIT=16'b0010111100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_18_LC_13_6_4  (
            .in0(N__35707),
            .in1(N__36079),
            .in2(N__36057),
            .in3(N__35983),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_13_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_18_LC_13_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_18_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40977),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52636),
            .ce(N__42037),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_13_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_13_6_6 .LUT_INIT=16'b1011111100001011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_18_LC_13_6_6  (
            .in0(N__35706),
            .in1(N__36078),
            .in2(N__36058),
            .in3(N__35982),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_13_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_19_LC_13_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_19_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40957),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52636),
            .ce(N__42037),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_13_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_13_7_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_0_LC_13_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_0_LC_13_7_0  (
            .in0(N__36922),
            .in1(N__38058),
            .in2(N__38752),
            .in3(N__38751),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_0 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_13_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_1_LC_13_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_1_LC_13_7_1  (
            .in0(N__36933),
            .in1(N__38031),
            .in2(_gnd_net_),
            .in3(N__35974),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_1 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_13_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_13_7_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_2_LC_13_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_2_LC_13_7_2  (
            .in0(N__36923),
            .in1(N__38421),
            .in2(_gnd_net_),
            .in3(N__35971),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_2 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_13_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_13_7_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_3_LC_13_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_3_LC_13_7_3  (
            .in0(N__36934),
            .in1(N__38397),
            .in2(_gnd_net_),
            .in3(N__35968),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_3 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_13_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_13_7_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_4_LC_13_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_4_LC_13_7_4  (
            .in0(N__36924),
            .in1(N__38373),
            .in2(_gnd_net_),
            .in3(N__35965),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_4 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_13_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_13_7_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_5_LC_13_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_5_LC_13_7_5  (
            .in0(N__36935),
            .in1(N__38349),
            .in2(_gnd_net_),
            .in3(N__35962),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_5 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_13_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_13_7_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_6_LC_13_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_6_LC_13_7_6  (
            .in0(N__36925),
            .in1(N__38322),
            .in2(_gnd_net_),
            .in3(N__35959),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_6 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_13_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_13_7_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_7_LC_13_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_7_LC_13_7_7  (
            .in0(N__36936),
            .in1(N__38301),
            .in2(_gnd_net_),
            .in3(N__35956),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_7 ),
            .clk(N__52630),
            .ce(N__36214),
            .sr(N__52174));
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_13_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_13_8_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_8_LC_13_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_8_LC_13_8_0  (
            .in0(N__36921),
            .in1(N__38271),
            .in2(_gnd_net_),
            .in3(N__36010),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_8 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_13_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_13_8_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_9_LC_13_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_9_LC_13_8_1  (
            .in0(N__36940),
            .in1(N__38247),
            .in2(_gnd_net_),
            .in3(N__36007),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_9 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_13_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_13_8_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_10_LC_13_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_10_LC_13_8_2  (
            .in0(N__36918),
            .in1(N__38586),
            .in2(_gnd_net_),
            .in3(N__36004),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_10 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_13_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_13_8_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_11_LC_13_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_11_LC_13_8_3  (
            .in0(N__36937),
            .in1(N__38562),
            .in2(_gnd_net_),
            .in3(N__36001),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_11 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_13_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_13_8_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_12_LC_13_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_12_LC_13_8_4  (
            .in0(N__36919),
            .in1(N__38538),
            .in2(_gnd_net_),
            .in3(N__35998),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_12 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_13_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_13_8_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_13_LC_13_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_13_LC_13_8_5  (
            .in0(N__36938),
            .in1(N__38514),
            .in2(_gnd_net_),
            .in3(N__35995),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_13 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_13_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_13_8_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_14_LC_13_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_14_LC_13_8_6  (
            .in0(N__36920),
            .in1(N__38487),
            .in2(_gnd_net_),
            .in3(N__35992),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_14 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_13_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_13_8_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_15_LC_13_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_15_LC_13_8_7  (
            .in0(N__36939),
            .in1(N__38460),
            .in2(_gnd_net_),
            .in3(N__35989),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_15 ),
            .clk(N__52623),
            .ce(N__36209),
            .sr(N__52176));
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_13_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_13_9_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_16_LC_13_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_16_LC_13_9_0  (
            .in0(N__36914),
            .in1(N__38854),
            .in2(_gnd_net_),
            .in3(N__35986),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_16 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_13_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_13_9_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_17_LC_13_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_17_LC_13_9_1  (
            .in0(N__36929),
            .in1(N__38871),
            .in2(_gnd_net_),
            .in3(N__36082),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_17 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_17 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_13_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_18_LC_13_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_18_LC_13_9_2  (
            .in0(N__36915),
            .in1(N__36077),
            .in2(_gnd_net_),
            .in3(N__36061),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_18 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_18 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_13_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_19_LC_13_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_19_LC_13_9_3  (
            .in0(N__36930),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__36031),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_19 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_19 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_13_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_13_9_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_20_LC_13_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_20_LC_13_9_4  (
            .in0(N__36916),
            .in1(N__38720),
            .in2(_gnd_net_),
            .in3(N__36028),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_20 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_20 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_13_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_13_9_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_21_LC_13_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_21_LC_13_9_5  (
            .in0(N__36931),
            .in1(N__38737),
            .in2(_gnd_net_),
            .in3(N__36025),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_21 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_21 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_13_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_22_LC_13_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_22_LC_13_9_6  (
            .in0(N__36917),
            .in1(N__39023),
            .in2(_gnd_net_),
            .in3(N__36022),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_22 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_22 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_13_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_23_LC_13_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_23_LC_13_9_7  (
            .in0(N__36932),
            .in1(N__39049),
            .in2(_gnd_net_),
            .in3(N__36019),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_23 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_23 ),
            .clk(N__52615),
            .ce(N__36213),
            .sr(N__52179));
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_13_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_13_10_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_24_LC_13_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_24_LC_13_10_0  (
            .in0(N__36909),
            .in1(N__38951),
            .in2(_gnd_net_),
            .in3(N__36016),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_24 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_13_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_13_10_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_25_LC_13_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_25_LC_13_10_1  (
            .in0(N__36926),
            .in1(N__38968),
            .in2(_gnd_net_),
            .in3(N__36013),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_25 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_25 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_13_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_13_10_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_26_LC_13_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_26_LC_13_10_2  (
            .in0(N__36910),
            .in1(N__39112),
            .in2(_gnd_net_),
            .in3(N__36172),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_26 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_13_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_13_10_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_27_LC_13_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_27_LC_13_10_3  (
            .in0(N__36927),
            .in1(N__39136),
            .in2(_gnd_net_),
            .in3(N__36169),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_27 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_27 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_13_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_28_LC_13_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_28_LC_13_10_4  (
            .in0(N__36911),
            .in1(N__36166),
            .in2(_gnd_net_),
            .in3(N__36151),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_28 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_28 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_13_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_13_10_5 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_29_LC_13_10_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_29_LC_13_10_5  (
            .in0(N__36928),
            .in1(N__36148),
            .in2(_gnd_net_),
            .in3(N__36133),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_29 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_29 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_13_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_13_10_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_30_LC_13_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_30_LC_13_10_6  (
            .in0(N__36912),
            .in1(N__36130),
            .in2(_gnd_net_),
            .in3(N__36112),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_30 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.counter_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_hc.counter_cry_30 ),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_13_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_13_10_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.counter_31_LC_13_10_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \phase_controller_inst1.stoper_hc.counter_31_LC_13_10_7  (
            .in0(N__36106),
            .in1(N__36913),
            .in2(_gnd_net_),
            .in3(N__36109),
            .lcout(\phase_controller_inst1.stoper_hc.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52606),
            .ce(N__36205),
            .sr(N__52188));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_30_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36249),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_11_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI36DN9_25_LC_13_11_1  (
            .in0(N__50485),
            .in1(N__36091),
            .in2(_gnd_net_),
            .in3(N__46576),
            .lcout(elapsed_time_ns_1_RNI36DN9_0_25),
            .ltout(elapsed_time_ns_1_RNI36DN9_0_25_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_13_11_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_13_11_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_25_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36085),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_11_3 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV2EN9_30_LC_13_11_3  (
            .in0(N__36250),
            .in1(_gnd_net_),
            .in2(N__50528),
            .in3(N__46960),
            .lcout(elapsed_time_ns_1_RNIV2EN9_0_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_13_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_13_11_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI03DN9_22_LC_13_11_4  (
            .in0(N__46927),
            .in1(N__36241),
            .in2(_gnd_net_),
            .in3(N__50484),
            .lcout(elapsed_time_ns_1_RNI03DN9_0_22),
            .ltout(elapsed_time_ns_1_RNI03DN9_0_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_11_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_11_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_22_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36235),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_13_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_13_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7ADN9_29_LC_13_11_6  (
            .in0(N__36232),
            .in1(N__46996),
            .in2(_gnd_net_),
            .in3(N__50486),
            .lcout(elapsed_time_ns_1_RNI7ADN9_0_29),
            .ltout(elapsed_time_ns_1_RNI7ADN9_0_29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_13_11_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_13_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_29_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36226),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.state_2_LC_13_12_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_2_LC_13_12_1 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_2_LC_13_12_1 .LUT_INIT=16'b1100111000001010;
    LogicCell40 \phase_controller_inst1.state_2_LC_13_12_1  (
            .in0(N__36293),
            .in1(N__36404),
            .in2(N__36274),
            .in3(N__50341),
            .lcout(\phase_controller_inst1.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52592),
            .ce(),
            .sr(N__52197));
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_12_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.start_timer_tr_RNO_0_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__36292),
            .in2(_gnd_net_),
            .in3(N__36268),
            .lcout(\phase_controller_inst1.start_timer_tr_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_12_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_12_5 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_RNILKNQ_LC_13_12_5  (
            .in0(N__36374),
            .in1(N__36356),
            .in2(_gnd_net_),
            .in3(N__38808),
            .lcout(\phase_controller_inst1.stoper_hc.un2_start_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_12_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_12_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.running_LC_13_12_6 .LUT_INIT=16'b1100111001001110;
    LogicCell40 \phase_controller_inst1.stoper_hc.running_LC_13_12_6  (
            .in0(N__36358),
            .in1(N__36375),
            .in2(N__38817),
            .in3(N__38775),
            .lcout(\phase_controller_inst1.stoper_hc.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52592),
            .ce(),
            .sr(N__52197));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_13_12_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_13_12_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNIMU8Q_LC_13_12_7  (
            .in0(N__52291),
            .in1(N__36357),
            .in2(_gnd_net_),
            .in3(N__38807),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_0 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNIUNOR_LC_13_13_0  (
            .in0(N__36497),
            .in1(_gnd_net_),
            .in2(N__38155),
            .in3(N__38136),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_168_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_13_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_tr_timer.running_LC_13_13_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_LC_13_13_1  (
            .in0(N__38137),
            .in1(N__36498),
            .in2(_gnd_net_),
            .in3(N__38154),
            .lcout(\delay_measurement_inst.delay_tr_timer.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52587),
            .ce(),
            .sr(N__52209));
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_13_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \delay_measurement_inst.delay_tr_timer.running_RNICNBI_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__36496),
            .in2(_gnd_net_),
            .in3(N__38150),
            .lcout(\delay_measurement_inst.delay_tr_timer.N_167_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.start_timer_hc_LC_13_13_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_13_4 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.start_timer_hc_LC_13_13_4 .LUT_INIT=16'b1100111011001010;
    LogicCell40 \phase_controller_inst1.start_timer_hc_LC_13_13_4  (
            .in0(N__36354),
            .in1(N__50332),
            .in2(N__36301),
            .in3(N__36405),
            .lcout(\phase_controller_inst1.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52587),
            .ce(),
            .sr(N__52209));
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_RNO_0_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(N__36353),
            .in2(_gnd_net_),
            .in3(N__38812),
            .lcout(),
            .ltout(\phase_controller_inst1.stoper_hc.un4_start_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_13_6 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.time_passed_LC_13_13_6 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \phase_controller_inst1.stoper_hc.time_passed_LC_13_13_6  (
            .in0(N__36376),
            .in1(N__36272),
            .in2(N__36361),
            .in3(N__38779),
            .lcout(\phase_controller_inst1.hc_time_passed ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52587),
            .ce(),
            .sr(N__52209));
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_13_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_13_7 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_hc.start_latched_LC_13_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36355),
            .lcout(\phase_controller_inst1.stoper_hc.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52587),
            .ce(),
            .sr(N__52209));
    defparam \phase_controller_inst1.state_1_LC_13_14_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.state_1_LC_13_14_2 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.state_1_LC_13_14_2 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \phase_controller_inst1.state_1_LC_13_14_2  (
            .in0(N__36334),
            .in1(N__36300),
            .in2(N__38100),
            .in3(N__36273),
            .lcout(\phase_controller_inst1.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52582),
            .ce(),
            .sr(N__52215));
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_14_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_14_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.stoper_tr.start_latched_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36776),
            .lcout(\phase_controller_inst1.stoper_tr.start_latchedZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52582),
            .ce(),
            .sr(N__52215));
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_15_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_15_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.start_latched_RNI7PP3_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38816),
            .lcout(\phase_controller_inst1.stoper_hc.start_latched_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_15_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_15_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \phase_controller_inst1.stoper_tr.start_latched_RNICIM41_LC_13_15_2  (
            .in0(N__36802),
            .in1(N__52293),
            .in2(_gnd_net_),
            .in3(N__36770),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticks_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_15_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_0_9_LC_13_15_4  (
            .in0(N__48116),
            .in1(N__49494),
            .in2(N__50113),
            .in3(N__48097),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIAC37_9_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48115),
            .lcout(\current_shift_inst.un4_control_input_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ26A_18_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47887),
            .lcout(\current_shift_inst.un4_control_input_1_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJS6A_20_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47758),
            .lcout(\current_shift_inst.un4_control_input_1_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_13_16_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_tr.target_ticks_0_LC_13_16_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.stoper_tr.target_ticks_0_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__36741),
            .in2(_gnd_net_),
            .in3(N__36703),
            .lcout(\phase_controller_inst1.stoper_tr.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52570),
            .ce(N__36594),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKS5A_12_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47275),
            .lcout(\current_shift_inst.un4_control_input_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKT6A_21_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44669),
            .lcout(\current_shift_inst.un4_control_input_1_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILT5A_13_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44044),
            .lcout(\current_shift_inst.un4_control_input_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILU6A_22_LC_13_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44561),
            .lcout(\current_shift_inst.un4_control_input_1_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV6A_23_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48050),
            .lcout(\current_shift_inst.un4_control_input_1_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIN07A_24_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47986),
            .lcout(\current_shift_inst.un4_control_input_1_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_16_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO06A_16_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44443),
            .lcout(\current_shift_inst.un4_control_input_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_cry_0_c_inv_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__37024),
            .in2(_gnd_net_),
            .in3(N__40030),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axb_0 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_13_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_13_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_1_LC_13_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_1_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__40021),
            .in2(_gnd_net_),
            .in3(N__36994),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_1 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_0 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_13_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_13_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_2_LC_13_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__40009),
            .in2(_gnd_net_),
            .in3(N__36970),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_2 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_1 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_13_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_13_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_3_LC_13_17_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_3_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(N__39997),
            .in2(_gnd_net_),
            .in3(N__36943),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_2 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_13_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_13_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_4_LC_13_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_4_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__39985),
            .in2(_gnd_net_),
            .in3(N__37219),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_3 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_13_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_13_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_5_LC_13_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_5_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(N__39970),
            .in2(_gnd_net_),
            .in3(N__37192),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_4 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_13_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_13_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_6_LC_13_17_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_6_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40153),
            .in3(N__37165),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_5 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_13_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_13_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_7_LC_13_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_7_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(N__40138),
            .in2(_gnd_net_),
            .in3(N__37132),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_6 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_7 ),
            .clk(N__52565),
            .ce(),
            .sr(N__52236));
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_13_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_13_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_8_LC_13_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_8_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__40126),
            .in2(_gnd_net_),
            .in3(N__37105),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_8 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_13_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_13_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_9_LC_13_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_9_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__40114),
            .in2(_gnd_net_),
            .in3(N__37081),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_8 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_13_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_13_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_10_LC_13_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_10_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__40102),
            .in2(_gnd_net_),
            .in3(N__37054),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_9 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_13_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_13_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_11_LC_13_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_11_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(N__40090),
            .in2(_gnd_net_),
            .in3(N__37027),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_10 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_13_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_13_18_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_12_LC_13_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_12_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__40078),
            .in2(_gnd_net_),
            .in3(N__37420),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_11 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_13_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_13_18_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_13_LC_13_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_13_LC_13_18_5  (
            .in0(_gnd_net_),
            .in1(N__40066),
            .in2(_gnd_net_),
            .in3(N__37390),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_12 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_13_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_13_18_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_14_LC_13_18_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_14_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40054),
            .in3(N__37360),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_13 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_13_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_15_LC_13_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_15_LC_13_18_7  (
            .in0(_gnd_net_),
            .in1(N__40252),
            .in2(_gnd_net_),
            .in3(N__37336),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_14 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_15 ),
            .clk(N__52561),
            .ce(),
            .sr(N__52240));
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_13_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_13_19_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_16_LC_13_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_16_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(N__40240),
            .in2(_gnd_net_),
            .in3(N__37309),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_16 ),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_13_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_17_LC_13_19_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_17_LC_13_19_1  (
            .in0(_gnd_net_),
            .in1(N__40228),
            .in2(_gnd_net_),
            .in3(N__37282),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_16 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_13_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_13_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_18_LC_13_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_18_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__40216),
            .in2(_gnd_net_),
            .in3(N__37279),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_17 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_13_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_13_19_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_19_LC_13_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_19_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(N__40204),
            .in2(_gnd_net_),
            .in3(N__37249),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_18 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_13_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_20_LC_13_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_20_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__40192),
            .in2(_gnd_net_),
            .in3(N__37246),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_19 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_13_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_21_LC_13_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_21_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(N__40180),
            .in2(_gnd_net_),
            .in3(N__37471),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_20 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_13_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_22_LC_13_19_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_22_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40168),
            .in3(N__37468),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_21 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_13_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_13_19_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_23_LC_13_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_23_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__40348),
            .in2(_gnd_net_),
            .in3(N__37465),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_22 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_23 ),
            .clk(N__52556),
            .ce(),
            .sr(N__52242));
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_13_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_13_20_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_24_LC_13_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_24_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__40336),
            .in2(_gnd_net_),
            .in3(N__37462),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_24 ),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_13_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_13_20_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_25_LC_13_20_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_25_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(N__40324),
            .in2(_gnd_net_),
            .in3(N__37459),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_24 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_13_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_13_20_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_26_LC_13_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_26_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(N__40312),
            .in2(_gnd_net_),
            .in3(N__37456),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_25 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_13_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_13_20_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_27_LC_13_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_27_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(N__40300),
            .in2(_gnd_net_),
            .in3(N__37453),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_26 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_13_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_13_20_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_28_LC_13_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_28_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(N__40288),
            .in2(_gnd_net_),
            .in3(N__37450),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_27 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_13_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_13_20_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_29_LC_13_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_29_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(N__40276),
            .in2(_gnd_net_),
            .in3(N__37447),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_28 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_13_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_13_20_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_30_LC_13_20_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_30_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40522),
            .in3(N__37765),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.PI_CTRL.error_control_2_cry_29 ),
            .carryout(\current_shift_inst.PI_CTRL.error_control_2_cry_30 ),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_13_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_13_20_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_31_LC_13_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_31_LC_13_20_7  (
            .in0(_gnd_net_),
            .in1(N__40261),
            .in2(_gnd_net_),
            .in3(N__37762),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52552),
            .ce(),
            .sr(N__52244));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_13_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_13_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_13_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIF9C4_12_LC_13_21_3  (
            .in0(N__37750),
            .in1(N__37759),
            .in2(N__37732),
            .in3(N__37740),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_11_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_13_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_13_21_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA4C4_10_LC_13_21_4  (
            .in0(N__37758),
            .in1(N__40440),
            .in2(N__40468),
            .in3(N__37749),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_13_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_13_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPL52_13_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(N__40503),
            .in2(_gnd_net_),
            .in3(N__40482),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_13_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_13_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_13_21_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIPCN8_12_LC_13_21_6  (
            .in0(N__37741),
            .in1(N__37731),
            .in2(N__37720),
            .in3(N__37717),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_13_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_13_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_13_21_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \current_shift_inst.PI_CTRL.integrator_RNICA8M_0_17_LC_13_21_7  (
            .in0(N__37703),
            .in1(N__37671),
            .in2(N__37633),
            .in3(N__37584),
            .lcout(\current_shift_inst.PI_CTRL.un3_enable_0_a3_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_13_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_13_22_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_18_LC_13_22_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_18_LC_13_22_0  (
            .in0(N__37527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52544),
            .ce(),
            .sr(N__52250));
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_13_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_13_22_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_24_LC_13_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_24_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37497),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52544),
            .ce(),
            .sr(N__52250));
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_13_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_13_22_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_22_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_22_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38004),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52544),
            .ce(),
            .sr(N__52250));
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_13_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_13_22_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_23_LC_13_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_23_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37962),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52544),
            .ce(),
            .sr(N__52250));
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_13_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_13_22_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_20_LC_13_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_20_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37938),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52544),
            .ce(),
            .sr(N__52250));
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_13_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_13_22_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_21_LC_13_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_21_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37908),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52544),
            .ce(),
            .sr(N__52250));
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_13_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_13_23_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_30_LC_13_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_30_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37878),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_13_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_13_23_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_29_LC_13_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_29_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37848),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_13_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_13_23_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_27_LC_13_23_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_27_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__37821),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_13_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_13_23_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_26_LC_13_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_26_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37788),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_13_23_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_13_23_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_31_LC_13_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_31_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38224),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_13_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_13_23_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_25_LC_13_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_25_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38205),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_13_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_13_23_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_28_LC_13_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_28_LC_13_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38181),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52542),
            .ce(),
            .sr(N__52255));
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_24_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_24_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_tr_LC_13_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_tr_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38127),
            .lcout(\delay_measurement_inst.stop_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38110),
            .ce(),
            .sr(N__52259));
    defparam \delay_measurement_inst.start_timer_tr_LC_13_24_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_tr_LC_13_24_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_tr_LC_13_24_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_tr_LC_13_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38126),
            .lcout(\delay_measurement_inst.start_timer_trZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38110),
            .ce(),
            .sr(N__52259));
    defparam \phase_controller_inst1.S2_LC_13_27_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.S2_LC_13_27_3 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S2_LC_13_27_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S2_LC_13_27_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38101),
            .lcout(s2_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52538),
            .ce(),
            .sr(N__52265));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_5_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_5_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_0_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(N__40696),
            .in2(N__38044),
            .in3(N__38062),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_0 ),
            .ltout(),
            .carryin(bfn_14_5_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_5_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_1_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(N__40555),
            .in2(N__38017),
            .in3(N__38035),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_5_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_5_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_2_LC_14_5_2  (
            .in0(_gnd_net_),
            .in1(N__38407),
            .in2(N__40357),
            .in3(N__38422),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_5_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_5_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_3_LC_14_5_3  (
            .in0(N__38401),
            .in1(N__40576),
            .in2(N__38383),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_5_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_5_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_4_LC_14_5_4  (
            .in0(_gnd_net_),
            .in1(N__38359),
            .in2(N__40564),
            .in3(N__38374),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_4 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_5_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_5_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_5_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__40549),
            .in2(N__38335),
            .in3(N__38353),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_5 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_5_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_5_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_5_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_6_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__38308),
            .in2(N__40585),
            .in3(N__38326),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_6 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_5_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_5_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_7_LC_14_5_7  (
            .in0(N__38302),
            .in1(N__40570),
            .in2(N__38287),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_7 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_6_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_6_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_8_LC_14_6_0  (
            .in0(_gnd_net_),
            .in1(N__40669),
            .in2(N__38257),
            .in3(N__38275),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_8 ),
            .ltout(),
            .carryin(bfn_14_6_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_6_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_9_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__40675),
            .in2(N__38233),
            .in3(N__38248),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_6_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_6_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_10_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(N__40681),
            .in2(N__38572),
            .in3(N__38590),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_10 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_6_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_6_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_11_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__40537),
            .in2(N__38548),
            .in3(N__38563),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_11 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_6_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_12_LC_14_6_4  (
            .in0(_gnd_net_),
            .in1(N__38524),
            .in2(N__40690),
            .in3(N__38539),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_12 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_6_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_13_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__40543),
            .in2(N__38500),
            .in3(N__38518),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_13 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_6_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_6_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_14_LC_14_6_6  (
            .in0(N__38488),
            .in1(N__40531),
            .in2(N__38473),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_14 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_6_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_6_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_inv_15_LC_14_6_7  (
            .in0(N__38464),
            .in1(N__41542),
            .in2(N__38446),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.counter_i_15 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_16_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(N__38596),
            .in2(N__38839),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_7_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_18_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(N__38437),
            .in2(N__38431),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_7_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_20_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(N__38602),
            .in2(N__38701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_7_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_22_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(N__39004),
            .in2(N__38674),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_7_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_24_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(N__38986),
            .in2(N__38932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_7_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_26_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(N__38911),
            .in2(N__39097),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_7_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_28_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(N__38662),
            .in2(N__38650),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_30_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(N__38635),
            .in2(N__38620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un6_running_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un6_running_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_8_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_LUT4_0_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38605),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_30_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_14_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_14_8_1 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_20_LC_14_8_1  (
            .in0(N__38691),
            .in1(N__38735),
            .in2(N__38721),
            .in3(N__38682),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_14_8_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_14_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_14_8_2 .LUT_INIT=16'b0111000100110000;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_16_LC_14_8_2  (
            .in0(N__38853),
            .in1(N__38870),
            .in2(N__38887),
            .in3(N__38902),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_14_8_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_14_8_3 .LUT_INIT=16'b1000111011001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_16_LC_14_8_3  (
            .in0(N__38901),
            .in1(N__38886),
            .in2(N__38872),
            .in3(N__38852),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_8_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIG23T9_4_LC_14_8_4  (
            .in0(N__43711),
            .in1(N__50529),
            .in2(_gnd_net_),
            .in3(N__38827),
            .lcout(elapsed_time_ns_1_RNIG23T9_0_4),
            .ltout(elapsed_time_ns_1_RNIG23T9_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_14_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_14_8_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_4_LC_14_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38821),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_8_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_8_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNIFAMA_30_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(N__38818),
            .in2(_gnd_net_),
            .in3(N__38763),
            .lcout(\phase_controller_inst1.stoper_hc.counter ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_14_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_14_8_7 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_20_LC_14_8_7  (
            .in0(N__38692),
            .in1(N__38736),
            .in2(N__38722),
            .in3(N__38683),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_14_9_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_20_LC_14_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_20_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40923),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52624),
            .ce(N__42033),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_14_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_21_LC_14_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_21_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41217),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52624),
            .ce(N__42033),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_14_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_14_9_4 .LUT_INIT=16'b0101110100000100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_22_LC_14_9_4  (
            .in0(N__39048),
            .in1(N__39034),
            .in2(N__39025),
            .in3(N__38995),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_14_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_22_LC_14_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_22_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41196),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52624),
            .ce(N__42033),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_14_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_14_9_6 .LUT_INIT=16'b1101111101000101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_22_LC_14_9_6  (
            .in0(N__39047),
            .in1(N__39033),
            .in2(N__39024),
            .in3(N__38994),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_14_9_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_23_LC_14_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_23_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41175),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52624),
            .ce(N__42033),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_14_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_14_10_0 .LUT_INIT=16'b0011101100000010;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_24_LC_14_10_0  (
            .in0(N__38977),
            .in1(N__38967),
            .in2(N__38953),
            .in3(N__38920),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_14_10_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_24_LC_14_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_24_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41157),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52616),
            .ce(N__42022),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_10_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_10_2 .LUT_INIT=16'b1011111100100011;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_24_LC_14_10_2  (
            .in0(N__38976),
            .in1(N__38966),
            .in2(N__38952),
            .in3(N__38919),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_14_10_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_25_LC_14_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_25_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41136),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52616),
            .ce(N__42022),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_10_4 .LUT_INIT=16'b0101000011010100;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_0_26_LC_14_10_4  (
            .in0(N__39135),
            .in1(N__39121),
            .in2(N__39085),
            .in3(N__39111),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_lt26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_14_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_26_LC_14_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_26_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41118),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52616),
            .ce(N__42022),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_10_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_10_6 .LUT_INIT=16'b1101010011110101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un6_running_cry_c_RNO_26_LC_14_10_6  (
            .in0(N__39134),
            .in1(N__39120),
            .in2(N__39084),
            .in3(N__39110),
            .lcout(\phase_controller_inst1.stoper_hc.un6_running_cry_c_RNOZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_14_10_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_14_10_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_27_LC_14_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_27_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41100),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52616),
            .ce(N__42022),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_11_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_11_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_0_LC_14_11_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_0_LC_14_11_0  (
            .in0(N__47246),
            .in1(N__42521),
            .in2(_gnd_net_),
            .in3(N__39070),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_0 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_11_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_11_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_1_LC_14_11_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_1_LC_14_11_1  (
            .in0(N__47238),
            .in1(N__41243),
            .in2(_gnd_net_),
            .in3(N__39067),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_0 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_1 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_11_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_11_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_2_LC_14_11_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_2_LC_14_11_2  (
            .in0(N__47247),
            .in1(N__39237),
            .in2(_gnd_net_),
            .in3(N__39064),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_1 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_2 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_11_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_11_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_3_LC_14_11_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_3_LC_14_11_3  (
            .in0(N__47239),
            .in1(N__39209),
            .in2(_gnd_net_),
            .in3(N__39061),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_3 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_11_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_11_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_4_LC_14_11_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_4_LC_14_11_4  (
            .in0(N__47248),
            .in1(N__39507),
            .in2(_gnd_net_),
            .in3(N__39058),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_4 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_11_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_11_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_5_LC_14_11_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_5_LC_14_11_5  (
            .in0(N__47240),
            .in1(N__39482),
            .in2(_gnd_net_),
            .in3(N__39055),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_5 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_11_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_11_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_6_LC_14_11_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_6_LC_14_11_6  (
            .in0(N__47249),
            .in1(N__39450),
            .in2(_gnd_net_),
            .in3(N__39052),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_6 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_11_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_11_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_7_LC_14_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_7_LC_14_11_7  (
            .in0(N__47241),
            .in1(N__39422),
            .in2(_gnd_net_),
            .in3(N__39163),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_7 ),
            .clk(N__52607),
            .ce(N__47367),
            .sr(N__52189));
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_12_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_12_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_8_LC_14_12_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_8_LC_14_12_0  (
            .in0(N__47237),
            .in1(N__39398),
            .in2(_gnd_net_),
            .in3(N__39160),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_12_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_8 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_12_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_9_LC_14_12_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_9_LC_14_12_1  (
            .in0(N__47245),
            .in1(N__39368),
            .in2(_gnd_net_),
            .in3(N__39157),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_9 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_12_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_10_LC_14_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_10_LC_14_12_2  (
            .in0(N__47234),
            .in1(N__39335),
            .in2(_gnd_net_),
            .in3(N__39154),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_9 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_10 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_12_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_12_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_11_LC_14_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_11_LC_14_12_3  (
            .in0(N__47242),
            .in1(N__39309),
            .in2(_gnd_net_),
            .in3(N__39151),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_11 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_12_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_12_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_12_LC_14_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_12_LC_14_12_4  (
            .in0(N__47235),
            .in1(N__39285),
            .in2(_gnd_net_),
            .in3(N__39148),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_12 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_12_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_12_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_13_LC_14_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_13_LC_14_12_5  (
            .in0(N__47243),
            .in1(N__39719),
            .in2(_gnd_net_),
            .in3(N__39145),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_13 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_12_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_14_LC_14_12_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_14_LC_14_12_6  (
            .in0(N__47236),
            .in1(N__39687),
            .in2(_gnd_net_),
            .in3(N__39142),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_14 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_12_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_15_LC_14_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_15_LC_14_12_7  (
            .in0(N__47244),
            .in1(N__39665),
            .in2(_gnd_net_),
            .in3(N__39139),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_15 ),
            .clk(N__52599),
            .ce(N__47360),
            .sr(N__52192));
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_13_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_16_LC_14_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_16_LC_14_13_0  (
            .in0(N__47254),
            .in1(N__39635),
            .in2(_gnd_net_),
            .in3(N__39190),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_16 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_13_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_17_LC_14_13_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_17_LC_14_13_1  (
            .in0(N__47250),
            .in1(N__39605),
            .in2(_gnd_net_),
            .in3(N__39187),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_17 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_13_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_18_LC_14_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_18_LC_14_13_2  (
            .in0(N__47255),
            .in1(N__39581),
            .in2(_gnd_net_),
            .in3(N__39184),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_17 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_18 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_19_LC_14_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_19_LC_14_13_3  (
            .in0(N__47251),
            .in1(N__39560),
            .in2(_gnd_net_),
            .in3(N__39181),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_19 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_13_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_20_LC_14_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_20_LC_14_13_4  (
            .in0(N__47256),
            .in1(N__39533),
            .in2(_gnd_net_),
            .in3(N__39178),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_20 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_21_LC_14_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_21_LC_14_13_5  (
            .in0(N__47252),
            .in1(N__39950),
            .in2(_gnd_net_),
            .in3(N__39175),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_21 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_13_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_22_LC_14_13_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_22_LC_14_13_6  (
            .in0(N__47257),
            .in1(N__39924),
            .in2(_gnd_net_),
            .in3(N__39172),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_22 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_13_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_23_LC_14_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_23_LC_14_13_7  (
            .in0(N__47253),
            .in1(N__39896),
            .in2(_gnd_net_),
            .in3(N__39169),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_23 ),
            .clk(N__52593),
            .ce(N__47371),
            .sr(N__52198));
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_14_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_24_LC_14_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_24_LC_14_14_0  (
            .in0(N__47228),
            .in1(N__39869),
            .in2(_gnd_net_),
            .in3(N__39166),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\current_shift_inst.timer_s1.counter_cry_24 ),
            .clk(N__52588),
            .ce(N__47353),
            .sr(N__52210));
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_25_LC_14_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_25_LC_14_14_1  (
            .in0(N__47232),
            .in1(N__39839),
            .in2(_gnd_net_),
            .in3(N__39268),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_25 ),
            .clk(N__52588),
            .ce(N__47353),
            .sr(N__52210));
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_14_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_26_LC_14_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_26_LC_14_14_2  (
            .in0(N__47229),
            .in1(N__39797),
            .in2(_gnd_net_),
            .in3(N__39265),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_25 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_26 ),
            .clk(N__52588),
            .ce(N__47353),
            .sr(N__52210));
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_27_LC_14_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_27_LC_14_14_3  (
            .in0(N__47233),
            .in1(N__39752),
            .in2(_gnd_net_),
            .in3(N__39262),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_27 ),
            .clk(N__52588),
            .ce(N__47353),
            .sr(N__52210));
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_28_LC_14_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \current_shift_inst.timer_s1.counter_28_LC_14_14_4  (
            .in0(N__47230),
            .in1(N__39816),
            .in2(_gnd_net_),
            .in3(N__39259),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.counter_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.counter_cry_28 ),
            .clk(N__52588),
            .ce(N__47353),
            .sr(N__52210));
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.counter_29_LC_14_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \current_shift_inst.timer_s1.counter_29_LC_14_14_5  (
            .in0(N__39771),
            .in1(N__47231),
            .in2(_gnd_net_),
            .in3(N__39256),
            .lcout(\current_shift_inst.timer_s1.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52588),
            .ce(N__47353),
            .sr(N__52210));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_15_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_3_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__42525),
            .in2(N__39249),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_3 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_4_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__41245),
            .in2(N__39220),
            .in3(N__39253),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_2 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_5_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__39513),
            .in2(N__39250),
            .in3(N__39223),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_3 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_6_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__39219),
            .in2(N__39489),
            .in3(N__39193),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_4 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_7_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__39514),
            .in2(N__39462),
            .in3(N__39493),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_5 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_8_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(N__39429),
            .in2(N__39490),
            .in3(N__39466),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_6 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_9_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(N__39399),
            .in2(N__39463),
            .in3(N__39436),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_7 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_10_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__39369),
            .in2(N__39433),
            .in3(N__39406),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_8 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_9 ),
            .clk(N__52583),
            .ce(N__44194),
            .sr(N__52216));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_11_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__39342),
            .in2(N__39403),
            .in3(N__39379),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_11 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_12_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__39315),
            .in2(N__39376),
            .in3(N__39349),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_10 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_13_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__39291),
            .in2(N__39346),
            .in3(N__39319),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_11 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_14_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__39316),
            .in2(N__39726),
            .in3(N__39295),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_12 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_15_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__39292),
            .in2(N__39699),
            .in3(N__39271),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_13 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_16_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_16_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__39666),
            .in2(N__39727),
            .in3(N__39703),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_14 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_17_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__39636),
            .in2(N__39700),
            .in3(N__39673),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_15 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_16_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_18_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__39606),
            .in2(N__39670),
            .in3(N__39646),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_16 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_17 ),
            .clk(N__52577),
            .ce(N__44193),
            .sr(N__52222));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_19_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__39582),
            .in2(N__39643),
            .in3(N__39616),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_19 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_20_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__39561),
            .in2(N__39613),
            .in3(N__39586),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_18 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_17_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_21_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__39583),
            .in2(N__39540),
            .in3(N__39565),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_19 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_17_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_22_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__39562),
            .in2(N__39957),
            .in3(N__39544),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_20 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_17_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_23_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__39930),
            .in2(N__39541),
            .in3(N__39517),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_21 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_17_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_24_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(N__39903),
            .in2(N__39958),
            .in3(N__39934),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_22 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_25_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__39931),
            .in2(N__39876),
            .in3(N__39910),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_23 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_17_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_26_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__39840),
            .in2(N__39907),
            .in3(N__39880),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_24 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_25 ),
            .clk(N__52571),
            .ce(N__44192),
            .sr(N__52230));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_27_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(N__39798),
            .in2(N__39877),
            .in3(N__39850),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_27 ),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .clk(N__52566),
            .ce(N__44191),
            .sr(N__52237));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_18_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_28_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__39753),
            .in2(N__39847),
            .in3(N__39820),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_26 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .clk(N__52566),
            .ce(N__44191),
            .sr(N__52237));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_18_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_29_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(N__39817),
            .in2(N__39802),
            .in3(N__39778),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_27 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .clk(N__52566),
            .ce(N__44191),
            .sr(N__52237));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_30_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(N__39775),
            .in2(N__39757),
            .in3(N__39733),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_28 ),
            .carryout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29 ),
            .clk(N__52566),
            .ce(N__44191),
            .sr(N__52237));
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_LUT4_0_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39730),
            .lcout(\current_shift_inst.timer_s1.un13_elapsed_time_ns_cry_29_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR47A_28_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44371),
            .lcout(\current_shift_inst.un4_control_input_1_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_18_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIS57A_29_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43396),
            .lcout(\current_shift_inst.un4_control_input_1_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_fast_31_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44213),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_fast_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52566),
            .ce(N__44191),
            .sr(N__52237));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_14_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_14_19_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNIT83B4_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__43102),
            .in2(N__43090),
            .in3(N__43089),
            .lcout(\current_shift_inst.control_input_1 ),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\current_shift_inst.control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_19_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_1_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__41461),
            .in2(_gnd_net_),
            .in3(N__40012),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_1 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_0 ),
            .carryout(\current_shift_inst.control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_19_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_2_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__41455),
            .in2(_gnd_net_),
            .in3(N__40000),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_2 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_1 ),
            .carryout(\current_shift_inst.control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_19_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_3_LC_14_19_3  (
            .in0(_gnd_net_),
            .in1(N__41449),
            .in2(_gnd_net_),
            .in3(N__39988),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_3 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_2 ),
            .carryout(\current_shift_inst.control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_14_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_14_19_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_4_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(N__41443),
            .in2(_gnd_net_),
            .in3(N__39973),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_4 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_3 ),
            .carryout(\current_shift_inst.control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_5_LC_14_19_5  (
            .in0(_gnd_net_),
            .in1(N__41437),
            .in2(_gnd_net_),
            .in3(N__39961),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_5 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_4 ),
            .carryout(\current_shift_inst.control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_14_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_14_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_6_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(N__41431),
            .in2(_gnd_net_),
            .in3(N__40141),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_6 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_5 ),
            .carryout(\current_shift_inst.control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_19_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_7_LC_14_19_7  (
            .in0(_gnd_net_),
            .in1(N__41533),
            .in2(_gnd_net_),
            .in3(N__40129),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_7 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_6 ),
            .carryout(\current_shift_inst.control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_20_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_8_LC_14_20_0  (
            .in0(_gnd_net_),
            .in1(N__43300),
            .in2(_gnd_net_),
            .in3(N__40117),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_20_0_),
            .carryout(\current_shift_inst.control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_14_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_14_20_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_9_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__43114),
            .in2(_gnd_net_),
            .in3(N__40105),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_9 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_8 ),
            .carryout(\current_shift_inst.control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_20_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_10_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(N__43066),
            .in2(_gnd_net_),
            .in3(N__40093),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_10 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_9 ),
            .carryout(\current_shift_inst.control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_20_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_11_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(N__43312),
            .in2(_gnd_net_),
            .in3(N__40081),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_11 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_10 ),
            .carryout(\current_shift_inst.control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_20_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_12_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__43273),
            .in2(_gnd_net_),
            .in3(N__40069),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_12 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_11 ),
            .carryout(\current_shift_inst.control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_13_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(N__41527),
            .in2(_gnd_net_),
            .in3(N__40057),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_13 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_12 ),
            .carryout(\current_shift_inst.control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_20_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_14_LC_14_20_6  (
            .in0(_gnd_net_),
            .in1(N__43291),
            .in2(_gnd_net_),
            .in3(N__40042),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_14 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_13 ),
            .carryout(\current_shift_inst.control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_20_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_15_LC_14_20_7  (
            .in0(_gnd_net_),
            .in1(N__43282),
            .in2(_gnd_net_),
            .in3(N__40243),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_15 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_14 ),
            .carryout(\current_shift_inst.control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_21_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_16_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__41497),
            .in2(_gnd_net_),
            .in3(N__40231),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_16 ),
            .ltout(),
            .carryin(bfn_14_21_0_),
            .carryout(\current_shift_inst.control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_21_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_17_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__41503),
            .in2(_gnd_net_),
            .in3(N__40219),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_17 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_16 ),
            .carryout(\current_shift_inst.control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_21_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_18_LC_14_21_2  (
            .in0(_gnd_net_),
            .in1(N__41668),
            .in2(_gnd_net_),
            .in3(N__40207),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_18 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_17 ),
            .carryout(\current_shift_inst.control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_21_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_19_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(N__43510),
            .in2(_gnd_net_),
            .in3(N__40195),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_19 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_18 ),
            .carryout(\current_shift_inst.control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_21_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_20_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(N__43429),
            .in2(_gnd_net_),
            .in3(N__40183),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_20 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_19 ),
            .carryout(\current_shift_inst.control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_14_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_14_21_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_21_LC_14_21_5  (
            .in0(_gnd_net_),
            .in1(N__41521),
            .in2(_gnd_net_),
            .in3(N__40171),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_21 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_20 ),
            .carryout(\current_shift_inst.control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_14_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_14_21_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_22_LC_14_21_6  (
            .in0(_gnd_net_),
            .in1(N__41509),
            .in2(_gnd_net_),
            .in3(N__40156),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_22 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_21 ),
            .carryout(\current_shift_inst.control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_21_7 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_21_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_23_LC_14_21_7  (
            .in0(_gnd_net_),
            .in1(N__49039),
            .in2(_gnd_net_),
            .in3(N__40339),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_23 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_22 ),
            .carryout(\current_shift_inst.control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_14_22_0 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_14_22_0 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_24_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(N__43264),
            .in2(_gnd_net_),
            .in3(N__40327),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_24 ),
            .ltout(),
            .carryin(bfn_14_22_0_),
            .carryout(\current_shift_inst.control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_14_22_1 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_14_22_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_25_LC_14_22_1  (
            .in0(_gnd_net_),
            .in1(N__41491),
            .in2(_gnd_net_),
            .in3(N__40315),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_25 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_24 ),
            .carryout(\current_shift_inst.control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_14_22_2 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_14_22_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_26_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(N__41515),
            .in2(_gnd_net_),
            .in3(N__40303),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_26 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_25 ),
            .carryout(\current_shift_inst.control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_14_22_3 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_14_22_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_27_LC_14_22_3  (
            .in0(_gnd_net_),
            .in1(N__41485),
            .in2(_gnd_net_),
            .in3(N__40291),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_27 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_26 ),
            .carryout(\current_shift_inst.control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_14_22_4 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_14_22_4 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_28_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__45367),
            .in2(_gnd_net_),
            .in3(N__40279),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_28 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_27 ),
            .carryout(\current_shift_inst.control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_14_22_5 .C_ON=1'b1;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_14_22_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_29_LC_14_22_5  (
            .in0(_gnd_net_),
            .in1(N__41767),
            .in2(_gnd_net_),
            .in3(N__40267),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_29 ),
            .ltout(),
            .carryin(\current_shift_inst.control_input_cry_28 ),
            .carryout(\current_shift_inst.control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_14_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_14_22_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \current_shift_inst.control_input_control_input_cry_29_c_RNIMVSI_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(N__49164),
            .in2(_gnd_net_),
            .in3(N__40264),
            .lcout(\current_shift_inst.control_input_31 ),
            .ltout(\current_shift_inst.control_input_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_14_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_14_22_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_2_axb_30_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40525),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.PI_CTRL.error_control_2_axbZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_14_23_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_14_23_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI2182_27_LC_14_23_2  (
            .in0(_gnd_net_),
            .in1(N__41646),
            .in2(_gnd_net_),
            .in3(N__41625),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_14_23_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_14_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNICPJ5_24_LC_14_23_3  (
            .in0(N__40392),
            .in1(N__40377),
            .in2(N__40510),
            .in3(N__40407),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_14_23_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_14_23_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOHB4_13_LC_14_23_5  (
            .in0(N__41761),
            .in1(N__40507),
            .in2(N__40489),
            .in3(N__41740),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_14_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_14_23_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_14_23_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIC8E4_10_LC_14_23_6  (
            .in0(N__40422),
            .in1(N__40467),
            .in2(N__40447),
            .in3(N__41661),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_14_23_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_14_23_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIROF4_24_LC_14_23_7  (
            .in0(N__40426),
            .in1(N__40408),
            .in2(N__40396),
            .in3(N__40378),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_12_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.start_timer_hc_LC_15_4_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_4_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.start_timer_hc_LC_15_4_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.start_timer_hc_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47563),
            .lcout(\delay_measurement_inst.start_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40366),
            .ce(),
            .sr(N__52168));
    defparam \delay_measurement_inst.stop_timer_hc_LC_15_4_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.stop_timer_hc_LC_15_4_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.stop_timer_hc_LC_15_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.stop_timer_hc_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47564),
            .lcout(\delay_measurement_inst.stop_timer_hcZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40366),
            .ce(),
            .sr(N__52168));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_5_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_2_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40629),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_5_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_6_LC_15_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40857),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_15_5_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_3_LC_15_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_3_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40605),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_15_5_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_7_LC_15_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_7_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40833),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_15_5_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_4_LC_15_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_4_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40905),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_5_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_5_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_LC_15_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40653),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_15_5_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_5_LC_15_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_5_LC_15_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40881),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52653),
            .ce(N__42043),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_15_6_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_15_6_0 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_13_LC_15_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_13_LC_15_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41079),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_6_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_11_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40740),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_15_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_14_LC_15_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_14_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41055),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_15_6_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_0_LC_15_6_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_0_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(N__42640),
            .in2(_gnd_net_),
            .in3(N__41833),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_6_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_12_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40716),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_15_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_10_LC_15_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_10_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40764),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_15_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_9_LC_15_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_9_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40788),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_6_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_8_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40812),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52647),
            .ce(N__42039),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_15_7_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_15_7_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_inv_LC_15_7_0  (
            .in0(N__42631),
            .in1(N__40663),
            .in2(N__41832),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.measured_delay_hc_i_31 ),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_15_7_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_15_7_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_0_c_RNIMTQQ_LC_15_7_1  (
            .in0(N__41797),
            .in1(N__41796),
            .in2(N__51646),
            .in3(N__40636),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_1),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_0 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_15_7_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_15_7_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_1_c_RNIO1TQ_LC_15_7_2  (
            .in0(N__41782),
            .in1(N__41781),
            .in2(N__51659),
            .in3(N__40612),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_2),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_15_7_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_15_7_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_2_c_RNIQ5VQ_LC_15_7_3  (
            .in0(N__42175),
            .in1(N__42174),
            .in2(N__51647),
            .in3(N__40588),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_3),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_15_7_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_15_7_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_15_7_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_3_c_RNIS91B_LC_15_7_4  (
            .in0(N__42160),
            .in1(N__42159),
            .in2(N__51660),
            .in3(N__40888),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_4),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_15_7_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_15_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_15_7_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_4_c_RNIUD3B_LC_15_7_5  (
            .in0(N__42145),
            .in1(N__42144),
            .in2(N__51648),
            .in3(N__40864),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_5),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_15_7_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_15_7_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_15_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_5_c_RNI0I5B_LC_15_7_6  (
            .in0(N__42130),
            .in1(N__42129),
            .in2(N__51661),
            .in3(N__40840),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_6),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_15_7_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_15_7_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_15_7_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_6_c_RNI2M7B_LC_15_7_7  (
            .in0(N__42109),
            .in1(N__42108),
            .in2(N__51649),
            .in3(N__40816),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_7),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_15_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_15_8_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_7_c_RNIB4AK_LC_15_8_0  (
            .in0(N__42088),
            .in1(N__42087),
            .in2(N__51590),
            .in3(N__40795),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_8),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_15_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_15_8_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_8_c_RNID8CK_LC_15_8_1  (
            .in0(N__42073),
            .in1(N__42072),
            .in2(N__51587),
            .in3(N__40771),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_9),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_8 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_15_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_15_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_9_c_RNIFCEK_LC_15_8_2  (
            .in0(N__42058),
            .in1(N__42057),
            .in2(N__51591),
            .in3(N__40747),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_10),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_15_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_15_8_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_10_c_RNIOLKH_LC_15_8_3  (
            .in0(N__42340),
            .in1(N__42339),
            .in2(N__51584),
            .in3(N__40723),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_11),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_15_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_15_8_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_11_c_RNIQPMH_LC_15_8_4  (
            .in0(N__42325),
            .in1(N__42324),
            .in2(N__51588),
            .in3(N__40699),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_12),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_15_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_15_8_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_12_c_RNISTOH_LC_15_8_5  (
            .in0(N__42310),
            .in1(N__42309),
            .in2(N__51585),
            .in3(N__41062),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_13),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_15_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_15_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_13_c_RNIU1RH_LC_15_8_6  (
            .in0(N__42295),
            .in1(N__42294),
            .in2(N__51589),
            .in3(N__41038),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_14),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_15_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_15_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_15_8_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_14_c_RNI06TH_LC_15_8_7  (
            .in0(N__42274),
            .in1(N__42273),
            .in2(N__51586),
            .in3(N__41035),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_15),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_15_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_15_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_15_c_RNI2AVH_LC_15_9_0  (
            .in0(N__42256),
            .in1(N__42255),
            .in2(N__51580),
            .in3(N__41008),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_16),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_15_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_15_9_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_16_c_RNI4E1I_LC_15_9_1  (
            .in0(N__42241),
            .in1(N__42240),
            .in2(N__51604),
            .in3(N__40981),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_17),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_16 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_15_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_15_9_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_17_c_RNIT0SI_LC_15_9_2  (
            .in0(N__42219),
            .in1(N__42226),
            .in2(N__51581),
            .in3(N__40960),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_18),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_15_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_15_9_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_18_c_RNIV4UI_LC_15_9_3  (
            .in0(N__42190),
            .in1(N__42189),
            .in2(N__51605),
            .in3(N__40933),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_19),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_15_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_15_9_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_19_c_RNI190J_LC_15_9_4  (
            .in0(N__42502),
            .in1(N__42498),
            .in2(N__51582),
            .in3(N__40912),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_20),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_15_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_15_9_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_20_c_RNIQRQJ_LC_15_9_5  (
            .in0(N__42484),
            .in1(N__42483),
            .in2(N__51606),
            .in3(N__41206),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_21),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_15_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_15_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_21_c_RNISVSJ_LC_15_9_6  (
            .in0(N__42460),
            .in1(N__42459),
            .in2(N__51583),
            .in3(N__41185),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_22),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_15_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_15_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_15_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_22_c_RNIU3VJ_LC_15_9_7  (
            .in0(N__42439),
            .in1(N__42438),
            .in2(N__51607),
            .in3(N__41164),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_23),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_15_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_15_10_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_23_c_RNI081K_LC_15_10_0  (
            .in0(N__42421),
            .in1(N__42420),
            .in2(N__51418),
            .in3(N__41146),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_24),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_15_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_15_10_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_24_c_RNI2C3K_LC_15_10_1  (
            .in0(N__42406),
            .in1(N__42405),
            .in2(N__51420),
            .in3(N__41125),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_25),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_24 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_15_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_15_10_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_25_c_RNI4G5K_LC_15_10_2  (
            .in0(N__42382),
            .in1(N__42381),
            .in2(N__51419),
            .in3(N__41107),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_26),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_15_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_15_10_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_26_c_RNI6K7K_LC_15_10_3  (
            .in0(N__42355),
            .in1(N__42354),
            .in2(N__51421),
            .in3(N__41089),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_27),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_15_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_15_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_LUT4_0_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41086),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_15_10_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_15_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_3_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41256),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_10_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIIF9N1_1_LC_15_10_6  (
            .in0(N__43725),
            .in1(N__41268),
            .in2(N__43710),
            .in3(N__46659),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_11_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIKFJE3_7_LC_15_11_1  (
            .in0(N__43849),
            .in1(N__41275),
            .in2(N__43825),
            .in3(N__42580),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_11_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_1_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45319),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52617),
            .ce(N__43959),
            .sr(N__52180));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_2_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45685),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52617),
            .ce(N__43959),
            .sr(N__52180));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIE03T9_2_LC_15_11_6  (
            .in0(N__41862),
            .in1(N__41269),
            .in2(_gnd_net_),
            .in3(N__50479),
            .lcout(elapsed_time_ns_1_RNIE03T9_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_11_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIF13T9_3_LC_15_11_7  (
            .in0(N__50480),
            .in1(N__41257),
            .in2(_gnd_net_),
            .in3(N__43729),
            .lcout(elapsed_time_ns_1_RNIF13T9_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_12_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITDHV_2_LC_15_12_0  (
            .in0(N__49446),
            .in1(N__48327),
            .in2(N__48223),
            .in3(N__48303),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITDHV_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_12_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_12_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_2_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41244),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52608),
            .ce(N__44196),
            .sr(N__52190));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3537_2_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48301),
            .lcout(\current_shift_inst.un4_control_input_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_12_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_RNO_LC_15_12_4  (
            .in0(N__43177),
            .in1(N__48326),
            .in2(_gnd_net_),
            .in3(N__48302),
            .lcout(\current_shift_inst.un10_control_input_cry_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_12_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNO_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__49447),
            .in2(_gnd_net_),
            .in3(N__44706),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_0_LC_15_12_7  (
            .in0(N__50754),
            .in1(N__49448),
            .in2(N__50112),
            .in3(N__44707),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_13_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_RNO_LC_15_13_0  (
            .in0(N__44149),
            .in1(N__43178),
            .in2(_gnd_net_),
            .in3(N__44160),
            .lcout(\current_shift_inst.un10_control_input_cry_2_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_13_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_13_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_RNO_LC_15_13_1  (
            .in0(N__44513),
            .in1(N__43182),
            .in2(_gnd_net_),
            .in3(N__44477),
            .lcout(\current_shift_inst.un10_control_input_cry_4_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_13_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_RNO_LC_15_13_2  (
            .in0(N__43183),
            .in1(N__47633),
            .in2(_gnd_net_),
            .in3(N__47660),
            .lcout(\current_shift_inst.un10_control_input_cry_5_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_13_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_RNO_LC_15_13_3  (
            .in0(N__48243),
            .in1(N__43184),
            .in2(_gnd_net_),
            .in3(N__48264),
            .lcout(\current_shift_inst.un10_control_input_cry_7_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_13_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_13_4 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_RNO_LC_15_13_4  (
            .in0(N__43181),
            .in1(N__48386),
            .in2(_gnd_net_),
            .in3(N__48350),
            .lcout(\current_shift_inst.un10_control_input_cry_3_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_15_13_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_15_13_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_RNO_LC_15_13_5  (
            .in0(N__43179),
            .in1(N__46794),
            .in2(_gnd_net_),
            .in3(N__46764),
            .lcout(\current_shift_inst.un10_control_input_cry_6_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_13_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_13_6 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_RNO_LC_15_13_6  (
            .in0(N__47315),
            .in1(N__43180),
            .in2(_gnd_net_),
            .in3(N__47285),
            .lcout(\current_shift_inst.un10_control_input_cry_11_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_13_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9B37_8_LC_15_13_7  (
            .in0(N__48242),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_14_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_RNO_LC_15_14_0  (
            .in0(N__44265),
            .in1(N__43219),
            .in2(_gnd_net_),
            .in3(N__44243),
            .lcout(\current_shift_inst.un10_control_input_cry_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_14_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_RNO_LC_15_14_1  (
            .in0(N__43220),
            .in1(N__47063),
            .in2(_gnd_net_),
            .in3(N__47037),
            .lcout(\current_shift_inst.un10_control_input_cry_10_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI6837_5_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44503),
            .lcout(\current_shift_inst.un4_control_input_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI8A37_7_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46787),
            .lcout(\current_shift_inst.un4_control_input_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_14_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_RNO_LC_15_14_4  (
            .in0(N__48117),
            .in1(N__43218),
            .in2(_gnd_net_),
            .in3(N__48083),
            .lcout(\current_shift_inst.un10_control_input_cry_8_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI4637_3_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44135),
            .lcout(\current_shift_inst.un4_control_input_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI7937_6_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47623),
            .lcout(\current_shift_inst.un4_control_input_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5737_4_LC_15_14_7  (
            .in0(N__48372),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un4_control_input_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_15_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_15_15_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_RNO_LC_15_15_0  (
            .in0(N__44045),
            .in1(N__43221),
            .in2(_gnd_net_),
            .in3(N__44021),
            .lcout(\current_shift_inst.un10_control_input_cry_12_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_RNO_LC_15_15_1  (
            .in0(N__43222),
            .in1(N__47720),
            .in2(_gnd_net_),
            .in3(N__47687),
            .lcout(\current_shift_inst.un10_control_input_cry_13_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_15_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP16A_17_LC_15_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47412),
            .lcout(\current_shift_inst.un4_control_input_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJR5A_11_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47054),
            .lcout(\current_shift_inst.un4_control_input_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_15_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_RNO_LC_15_15_4  (
            .in0(N__47088),
            .in1(N__43223),
            .in2(_gnd_net_),
            .in3(N__47123),
            .lcout(\current_shift_inst.un10_control_input_cry_14_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_15_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINV5A_15_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47087),
            .lcout(\current_shift_inst.un4_control_input_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMU5A_14_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47719),
            .lcout(\current_shift_inst.un4_control_input_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIIQ5A_10_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44264),
            .lcout(\current_shift_inst.un4_control_input_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_0_c_LC_15_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_0_c_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__50744),
            .in2(N__42555),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_1_c_LC_15_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_1_c_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__51405),
            .in2(N__41296),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_0 ),
            .carryout(\current_shift_inst.un10_control_input_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_2_c_LC_15_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_2_c_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__41284),
            .in2(N__51502),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_1 ),
            .carryout(\current_shift_inst.un10_control_input_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_3_c_LC_15_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_3_c_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__51409),
            .in2(N__41383),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_2 ),
            .carryout(\current_shift_inst.un10_control_input_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_4_c_LC_15_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_4_c_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(N__41371),
            .in2(N__51503),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_3 ),
            .carryout(\current_shift_inst.un10_control_input_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_16_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_5_c_LC_15_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_5_c_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__51413),
            .in2(N__41362),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_4 ),
            .carryout(\current_shift_inst.un10_control_input_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_16_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_6_c_LC_15_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_6_c_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__41350),
            .in2(N__51504),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_5 ),
            .carryout(\current_shift_inst.un10_control_input_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_16_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_7_c_LC_15_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_7_c_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__51417),
            .in2(N__41341),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_6 ),
            .carryout(\current_shift_inst.un10_control_input_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_8_c_LC_15_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_8_c_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__51401),
            .in2(N__41329),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_9_c_LC_15_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_9_c_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__41317),
            .in2(N__51501),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_8 ),
            .carryout(\current_shift_inst.un10_control_input_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_10_c_LC_15_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_10_c_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__51389),
            .in2(N__41308),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_9 ),
            .carryout(\current_shift_inst.un10_control_input_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_11_c_LC_15_17_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_11_c_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__41425),
            .in2(N__51498),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_10 ),
            .carryout(\current_shift_inst.un10_control_input_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_12_c_LC_15_17_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_12_c_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__51393),
            .in2(N__41416),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_11 ),
            .carryout(\current_shift_inst.un10_control_input_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_13_c_LC_15_17_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_13_c_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__41404),
            .in2(N__51499),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_12 ),
            .carryout(\current_shift_inst.un10_control_input_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_14_c_LC_15_17_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_14_c_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__51397),
            .in2(N__41395),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_13 ),
            .carryout(\current_shift_inst.un10_control_input_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_LC_15_17_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__42931),
            .in2(N__51500),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_14 ),
            .carryout(\current_shift_inst.un10_control_input_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_LC_15_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__51338),
            .in2(N__43027),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_LC_15_18_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(N__51342),
            .in2(N__42925),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_16 ),
            .carryout(\current_shift_inst.un10_control_input_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_LC_15_18_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__51339),
            .in2(N__42574),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_17 ),
            .carryout(\current_shift_inst.un10_control_input_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_LC_15_18_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__51343),
            .in2(N__43018),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_18 ),
            .carryout(\current_shift_inst.un10_control_input_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_LC_15_18_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(N__51340),
            .in2(N__42913),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_19 ),
            .carryout(\current_shift_inst.un10_control_input_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_LC_15_18_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__51344),
            .in2(N__43036),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_20 ),
            .carryout(\current_shift_inst.un10_control_input_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_LC_15_18_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(N__51341),
            .in2(N__43054),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_21 ),
            .carryout(\current_shift_inst.un10_control_input_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_LC_15_18_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_LC_15_18_7  (
            .in0(_gnd_net_),
            .in1(N__51345),
            .in2(N__43003),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_22 ),
            .carryout(\current_shift_inst.un10_control_input_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_LC_15_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(N__51220),
            .in2(N__43126),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_19_0_),
            .carryout(\current_shift_inst.un10_control_input_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_LC_15_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(N__43045),
            .in2(N__51386),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_24 ),
            .carryout(\current_shift_inst.un10_control_input_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_LC_15_19_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(N__51224),
            .in2(N__42994),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_25 ),
            .carryout(\current_shift_inst.un10_control_input_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_LC_15_19_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_LC_15_19_3  (
            .in0(_gnd_net_),
            .in1(N__43252),
            .in2(N__51387),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_26 ),
            .carryout(\current_shift_inst.un10_control_input_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_LC_15_19_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_LC_15_19_4  (
            .in0(_gnd_net_),
            .in1(N__51228),
            .in2(N__42985),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_27 ),
            .carryout(\current_shift_inst.un10_control_input_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_LC_15_19_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(N__42976),
            .in2(N__51388),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_28 ),
            .carryout(\current_shift_inst.un10_control_input_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_LC_15_19_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(N__51232),
            .in2(N__41479),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un10_control_input_cry_29 ),
            .carryout(\current_shift_inst.un10_control_input_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(N__49496),
            .in2(_gnd_net_),
            .in3(N__41464),
            .lcout(\current_shift_inst.un10_control_input_cry_30_c_RNI4B5IZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_20_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNI1GKD3_LC_15_20_0  (
            .in0(N__48136),
            .in1(N__44944),
            .in2(_gnd_net_),
            .in3(N__49109),
            .lcout(\current_shift_inst.control_input_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_15_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_15_20_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNI92B23_LC_15_20_1  (
            .in0(N__49110),
            .in1(N__48577),
            .in2(_gnd_net_),
            .in3(N__44917),
            .lcout(\current_shift_inst.control_input_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_20_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIHK1N3_LC_15_20_2  (
            .in0(N__48553),
            .in1(N__44902),
            .in2(_gnd_net_),
            .in3(N__49111),
            .lcout(\current_shift_inst.control_input_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_20_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIP6OB3_LC_15_20_3  (
            .in0(N__49112),
            .in1(N__44887),
            .in2(_gnd_net_),
            .in3(N__48529),
            .lcout(\current_shift_inst.control_input_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_20_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNI1PE03_LC_15_20_4  (
            .in0(N__44857),
            .in1(N__48499),
            .in2(_gnd_net_),
            .in3(N__49113),
            .lcout(\current_shift_inst.control_input_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_15_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_15_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_15_20_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNI50F14_LC_15_20_5  (
            .in0(N__49114),
            .in1(N__44833),
            .in2(_gnd_net_),
            .in3(N__48472),
            .lcout(\current_shift_inst.control_input_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_20_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIDI5M3_LC_15_20_6  (
            .in0(N__48445),
            .in1(N__44803),
            .in2(_gnd_net_),
            .in3(N__49115),
            .lcout(\current_shift_inst.control_input_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_20_7 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIPCGN2_LC_15_20_7  (
            .in0(N__49116),
            .in1(N__45034),
            .in2(_gnd_net_),
            .in3(N__48685),
            .lcout(\current_shift_inst.control_input_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_21_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIH2CP2_LC_15_21_0  (
            .in0(N__45178),
            .in1(N__48865),
            .in2(_gnd_net_),
            .in3(N__49157),
            .lcout(\current_shift_inst.control_input_axb_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_21_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNILSV03_LC_15_21_1  (
            .in0(N__49160),
            .in1(N__50155),
            .in2(_gnd_net_),
            .in3(N__45430),
            .lcout(\current_shift_inst.control_input_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_21_2 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIPK2E3_LC_15_21_2  (
            .in0(N__45160),
            .in1(N__48841),
            .in2(_gnd_net_),
            .in3(N__49158),
            .lcout(\current_shift_inst.control_input_axb_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_21_3 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNILKDA3_LC_15_21_3  (
            .in0(N__49156),
            .in1(N__48970),
            .in2(_gnd_net_),
            .in3(N__45277),
            .lcout(\current_shift_inst.control_input_axb_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_15_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_15_21_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNID2NL3_LC_15_21_4  (
            .in0(N__44968),
            .in1(N__48604),
            .in2(_gnd_net_),
            .in3(N__49155),
            .lcout(\current_shift_inst.control_input_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_21_5 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNIHB6C3_LC_15_21_5  (
            .in0(N__49159),
            .in1(N__50179),
            .in2(_gnd_net_),
            .in3(N__45451),
            .lcout(\current_shift_inst.control_input_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_15_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_15_21_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIPIEU2_LC_15_21_7  (
            .in0(N__49161),
            .in1(N__50128),
            .in2(_gnd_net_),
            .in3(N__45397),
            .lcout(\current_shift_inst.control_input_axb_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_22_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_22_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_22_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_0_LC_15_22_0  (
            .in0(N__49163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_15_22_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_15_22_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_15_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIOL62_17_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__41688),
            .in2(_gnd_net_),
            .in3(N__41760),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_0_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_15_22_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_15_22_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIT7H5_18_LC_15_22_2  (
            .in0(N__41716),
            .in1(N__41739),
            .in2(N__41719),
            .in3(N__41704),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_15_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_22_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILJ72_21_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(N__41715),
            .in2(_gnd_net_),
            .in3(N__41703),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_15_22_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_15_22_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_15_22_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI7TP8_19_LC_15_22_6  (
            .in0(N__41689),
            .in1(N__41607),
            .in2(N__41677),
            .in3(N__41674),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o3_17_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_22_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_22_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_22_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIPB8R2_LC_15_22_7  (
            .in0(N__45250),
            .in1(N__48943),
            .in2(_gnd_net_),
            .in3(N__49162),
            .lcout(\current_shift_inst.control_input_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_15_23_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_15_23_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_15_23_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNITQF4_19_LC_15_23_0  (
            .in0(N__41662),
            .in1(N__41647),
            .in2(N__41632),
            .in3(N__41611),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_a3_11_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_15_23_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_15_23_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_15_23_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_12_LC_15_23_1  (
            .in0(N__41590),
            .in1(N__41584),
            .in2(N__41572),
            .in3(N__41569),
            .lcout(\current_shift_inst.PI_CTRL.N_160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_6_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_6_5 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_15_LC_16_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41559),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52654),
            .ce(N__42038),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_7_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_7_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI04EN9_31_LC_16_7_0  (
            .in0(N__46702),
            .in1(N__42635),
            .in2(_gnd_net_),
            .in3(N__50547),
            .lcout(elapsed_time_ns_1_RNI04EN9_0_31),
            .ltout(elapsed_time_ns_1_RNI04EN9_0_31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_16_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \phase_controller_inst2.stoper_hc.target_ticks_0_LC_16_7_1 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \phase_controller_inst2.stoper_hc.target_ticks_0_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41968),
            .in3(N__41831),
            .lcout(\phase_controller_inst2.stoper_hc.target_ticksZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52648),
            .ce(N__41952),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI25DN9_24_LC_16_7_2  (
            .in0(N__43579),
            .in1(N__46978),
            .in2(_gnd_net_),
            .in3(N__50548),
            .lcout(elapsed_time_ns_1_RNI25DN9_0_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_16_8_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_16_8_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1_c_inv_LC_16_8_0  (
            .in0(_gnd_net_),
            .in1(N__42630),
            .in2(N__41875),
            .in3(N__46648),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_1 ),
            .ltout(),
            .carryin(bfn_16_8_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_16_8_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_16_8_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_inv_LC_16_8_1  (
            .in0(_gnd_net_),
            .in1(N__41848),
            .in2(_gnd_net_),
            .in3(N__41866),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axb_2 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_1 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_16_8_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_16_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2_c_RNIUTRF_LC_16_8_2  (
            .in0(_gnd_net_),
            .in1(N__41842),
            .in2(_gnd_net_),
            .in3(N__41809),
            .lcout(\phase_controller_inst1.stoper_hc.target_ticksZ0Z_1 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_2 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_16_8_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_16_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSF_LC_16_8_3  (
            .in0(_gnd_net_),
            .in1(N__41806),
            .in2(_gnd_net_),
            .in3(N__41785),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3_c_RNIVVSFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_3 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_16_8_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_16_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UF_LC_16_8_4  (
            .in0(_gnd_net_),
            .in1(N__43516),
            .in2(_gnd_net_),
            .in3(N__41770),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4_c_RNI02UFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_4 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_16_8_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_16_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VF_LC_16_8_5  (
            .in0(_gnd_net_),
            .in1(N__43774),
            .in2(_gnd_net_),
            .in3(N__42163),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5_c_RNI14VFZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_5 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_16_8_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_16_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNI26_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(N__43588),
            .in2(_gnd_net_),
            .in3(N__42148),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6_c_RNIZ0Z26 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_6 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_16_8_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_16_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNI381_LC_16_8_7  (
            .in0(_gnd_net_),
            .in1(N__43663),
            .in2(_gnd_net_),
            .in3(N__42133),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7_c_RNIZ0Z381 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_7 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_16_9_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_16_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4A2_LC_16_9_0  (
            .in0(_gnd_net_),
            .in1(N__43633),
            .in2(_gnd_net_),
            .in3(N__42112),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_8_c_RNI4AZ0Z2 ),
            .ltout(),
            .carryin(bfn_16_9_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_16_9_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_16_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5C3_LC_16_9_1  (
            .in0(_gnd_net_),
            .in1(N__43678),
            .in2(_gnd_net_),
            .in3(N__42091),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9_c_RNI5CZ0Z3 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_9 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_16_9_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_16_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDO49_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__43759),
            .in2(_gnd_net_),
            .in3(N__42076),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10_c_RNIDOZ0Z49 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_10 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_16_9_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_16_9_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQ59_LC_16_9_3  (
            .in0(_gnd_net_),
            .in1(N__43627),
            .in2(_gnd_net_),
            .in3(N__42061),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11_c_RNIEQZ0Z59 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_11 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_16_9_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_16_9_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFS69_LC_16_9_4  (
            .in0(_gnd_net_),
            .in1(N__49003),
            .in2(_gnd_net_),
            .in3(N__42046),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12_c_RNIFSZ0Z69 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_12 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_16_9_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_16_9_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGU79_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__48994),
            .in2(_gnd_net_),
            .in3(N__42328),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13_c_RNIGUZ0Z79 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_13 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_16_9_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_16_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIH099_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__43744),
            .in2(_gnd_net_),
            .in3(N__42313),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14_c_RNIHZ0Z099 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_14 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_16_9_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_16_9_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_16_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2A9_LC_16_9_7  (
            .in0(_gnd_net_),
            .in1(N__43648),
            .in2(_gnd_net_),
            .in3(N__42298),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15_c_RNII2AZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_15 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_16_10_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_16_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4B9_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__43555),
            .in2(_gnd_net_),
            .in3(N__42277),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_16_c_RNIJ4BZ0Z9 ),
            .ltout(),
            .carryin(bfn_16_10_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_16_10_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_16_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6C9_LC_16_10_1  (
            .in0(_gnd_net_),
            .in1(N__46537),
            .in2(_gnd_net_),
            .in3(N__42259),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17_c_RNIK6CZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_17 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_16_10_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_16_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8D9_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__46717),
            .in2(_gnd_net_),
            .in3(N__42244),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18_c_RNIL8DZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_18 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_16_10_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_16_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAE9_LC_16_10_3  (
            .in0(_gnd_net_),
            .in1(N__43534),
            .in2(_gnd_net_),
            .in3(N__42229),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19_c_RNIMAEZ0Z9 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_19 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_16_10_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_16_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7A_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__47593),
            .in2(_gnd_net_),
            .in3(N__42205),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20_c_RNIER7AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_20 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_16_10_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_16_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8A_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__42202),
            .in2(_gnd_net_),
            .in3(N__42178),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21_c_RNIFT8AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_21 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_16_10_6 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_16_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9A_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__50629),
            .in2(_gnd_net_),
            .in3(N__42487),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22_c_RNIGV9AZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_22 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_16_10_7 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_16_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BA_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__43567),
            .in2(_gnd_net_),
            .in3(N__42472),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23_c_RNIH1BAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_23 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_16_11_0 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_16_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CA_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__42469),
            .in2(_gnd_net_),
            .in3(N__42442),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_24_c_RNII3CAZ0 ),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_16_11_1 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_16_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DA_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__50605),
            .in2(_gnd_net_),
            .in3(N__42424),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25_c_RNIJ5DAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_25 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_16_11_2 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_16_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EA_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(N__45346),
            .in2(_gnd_net_),
            .in3(N__42409),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26_c_RNIK7EAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_26 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_16_11_3 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_16_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FA_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(N__46237),
            .in2(_gnd_net_),
            .in3(N__42394),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27_c_RNIL9FAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_27 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_16_11_4 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_16_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGA_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(N__42391),
            .in2(_gnd_net_),
            .in3(N__42370),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28_c_RNIMBGAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_28 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_16_11_5 .C_ON=1'b1;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_16_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHA_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(N__42367),
            .in2(_gnd_net_),
            .in3(N__42343),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29_c_RNINDHAZ0 ),
            .ltout(),
            .carryin(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_29 ),
            .carryout(\phase_controller_inst1.stoper_hc.un3_target_ticks_cry_30 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_16_11_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_16_11_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \phase_controller_inst1.stoper_hc.target_ticks_1_cry_27_c_RNIV62L_LC_16_11_6  (
            .in0(N__42646),
            .in1(N__42639),
            .in2(_gnd_net_),
            .in3(N__42604),
            .lcout(phase_controller_inst1_stoper_hc_target_ticks_1_i_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_11_7 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIVTKR_5_LC_16_11_7  (
            .in0(N__43878),
            .in1(N__43863),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_16_12_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_16_12_0 .LUT_INIT=16'b1011000110110001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_0_19_LC_16_12_0  (
            .in0(N__49497),
            .in1(N__47869),
            .in2(N__47830),
            .in3(N__50077),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_12_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_12_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNILV7A_31_LC_16_12_2  (
            .in0(N__49498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50076),
            .lcout(\current_shift_inst.un38_control_input_axb_31_s0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_12_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_12_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_18_c_RNO_LC_16_12_3  (
            .in0(N__47868),
            .in1(N__43176),
            .in2(_gnd_net_),
            .in3(N__47825),
            .lcout(\current_shift_inst.un10_control_input_cry_18_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_12_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_1_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44077),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_i_1 ),
            .ltout(\current_shift_inst.elapsed_time_ns_s1_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_12_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_12_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNINRRH_1_LC_16_12_5  (
            .in0(N__44078),
            .in1(_gnd_net_),
            .in2(N__42559),
            .in3(N__43175),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNINRRH_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_12_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_12_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_rep1_LC_16_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44230),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52618),
            .ce(N__44197),
            .sr(N__52181));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_12_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_12_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_1_LC_16_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42529),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52618),
            .ce(N__44197),
            .sr(N__52181));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_13_0 .C_ON=1'b1;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI596E_2_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(N__42721),
            .in2(N__44118),
            .in3(N__44114),
            .lcout(\current_shift_inst.un4_control_input1_2 ),
            .ltout(),
            .carryin(bfn_16_13_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_13_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_1_c_RNI4M9L_LC_16_13_1  (
            .in0(_gnd_net_),
            .in1(N__42715),
            .in2(_gnd_net_),
            .in3(N__42709),
            .lcout(\current_shift_inst.un4_control_input1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_1 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_13_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_2_c_RNI6PAL_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__42706),
            .in2(_gnd_net_),
            .in3(N__42700),
            .lcout(\current_shift_inst.un4_control_input1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_2 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_13_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_3_c_RNI8SBL_LC_16_13_3  (
            .in0(_gnd_net_),
            .in1(N__42697),
            .in2(_gnd_net_),
            .in3(N__42691),
            .lcout(\current_shift_inst.un4_control_input1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_3 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_13_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_4_c_RNIAVCL_LC_16_13_4  (
            .in0(_gnd_net_),
            .in1(N__42688),
            .in2(_gnd_net_),
            .in3(N__42682),
            .lcout(\current_shift_inst.un4_control_input1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_4 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_13_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_5_c_RNIC2EL_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__42679),
            .in2(_gnd_net_),
            .in3(N__42673),
            .lcout(\current_shift_inst.un4_control_input1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_5 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_13_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_6_c_RNIE5FL_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__42670),
            .in2(_gnd_net_),
            .in3(N__42664),
            .lcout(\current_shift_inst.un4_control_input1_8 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_6 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_13_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_7_c_RNIG8GL_LC_16_13_7  (
            .in0(_gnd_net_),
            .in1(N__42661),
            .in2(_gnd_net_),
            .in3(N__42649),
            .lcout(\current_shift_inst.un4_control_input1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_7 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_14_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_8_c_RNIPOJO_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__42823),
            .in2(_gnd_net_),
            .in3(N__42817),
            .lcout(\current_shift_inst.un4_control_input1_10 ),
            .ltout(),
            .carryin(bfn_16_14_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_14_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_9_c_RNIRRKO_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(N__42814),
            .in2(_gnd_net_),
            .in3(N__42808),
            .lcout(\current_shift_inst.un4_control_input1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_9 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_14_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_10_c_RNI4CAD_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__42805),
            .in2(_gnd_net_),
            .in3(N__42793),
            .lcout(\current_shift_inst.un4_control_input1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_10 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_14_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_11_c_RNI6FBD_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(N__42790),
            .in2(_gnd_net_),
            .in3(N__42778),
            .lcout(\current_shift_inst.un4_control_input1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_11 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_14_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_12_c_RNI8ICD_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__42775),
            .in2(_gnd_net_),
            .in3(N__42769),
            .lcout(\current_shift_inst.un4_control_input1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_12 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_14_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_13_c_RNIALDD_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(N__42766),
            .in2(_gnd_net_),
            .in3(N__42760),
            .lcout(\current_shift_inst.un4_control_input1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_13 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_14_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_14_c_RNICOED_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__42757),
            .in2(_gnd_net_),
            .in3(N__42745),
            .lcout(\current_shift_inst.un4_control_input1_16 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_14 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_14_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_15_c_RNIERFD_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(N__42742),
            .in2(_gnd_net_),
            .in3(N__42736),
            .lcout(\current_shift_inst.un4_control_input1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_15 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_15_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_16_c_RNIGUGD_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__42733),
            .in2(_gnd_net_),
            .in3(N__42724),
            .lcout(\current_shift_inst.un4_control_input1_18 ),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_17 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_15_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_17_c_RNII1ID_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__44005),
            .in2(_gnd_net_),
            .in3(N__42904),
            .lcout(\current_shift_inst.un4_control_input1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_17 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_18 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_15_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_18_c_RNIBSJD_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__42901),
            .in2(_gnd_net_),
            .in3(N__42892),
            .lcout(\current_shift_inst.un4_control_input1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_18 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_19 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_15_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_15_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_19_c_RNIDVKD_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__42889),
            .in2(_gnd_net_),
            .in3(N__42877),
            .lcout(\current_shift_inst.un4_control_input1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_19 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_20 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_15_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_15_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_20_c_RNI6HEE_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__42874),
            .in2(_gnd_net_),
            .in3(N__42862),
            .lcout(\current_shift_inst.un4_control_input1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_20 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_21 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_15_5 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_15_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_21_c_RNI8KFE_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__42859),
            .in2(_gnd_net_),
            .in3(N__42847),
            .lcout(\current_shift_inst.un4_control_input1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_21 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_22 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_15_6 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_22_c_RNIANGE_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__42844),
            .in2(_gnd_net_),
            .in3(N__42832),
            .lcout(\current_shift_inst.un4_control_input1_24 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_22 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_23 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_15_7 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_23_c_RNICQHE_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__46816),
            .in2(_gnd_net_),
            .in3(N__42829),
            .lcout(\current_shift_inst.un4_control_input1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_23 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_24 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_16_0 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_24_c_RNIETIE_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__43009),
            .in2(_gnd_net_),
            .in3(N__42826),
            .lcout(\current_shift_inst.un4_control_input1_26 ),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\current_shift_inst.un4_control_input_1_cry_25 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_16_1 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_25_c_RNIG0KE_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__43438),
            .in2(_gnd_net_),
            .in3(N__42970),
            .lcout(\current_shift_inst.un4_control_input1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_25 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_26 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_16_2 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_26_c_RNII3LE_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__42967),
            .in2(_gnd_net_),
            .in3(N__42955),
            .lcout(\current_shift_inst.un4_control_input1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_26 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_27 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_16_3 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_27_c_RNIK6ME_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__42952),
            .in2(_gnd_net_),
            .in3(N__42940),
            .lcout(\current_shift_inst.un4_control_input1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_27 ),
            .carryout(\current_shift_inst.un4_control_input_1_cry_28 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_16_4 .C_ON=1'b1;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_28_c_RNID1OE_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__43246),
            .in2(_gnd_net_),
            .in3(N__42937),
            .lcout(\current_shift_inst.un4_control_input1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un4_control_input_1_cry_28 ),
            .carryout(\current_shift_inst.un4_control_input1_31 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.un4_control_input1_31_THRU_LUT4_0_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42934),
            .lcout(\current_shift_inst.un4_control_input1_31_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_15_c_RNO_LC_16_16_6  (
            .in0(N__43229),
            .in1(N__44453),
            .in2(_gnd_net_),
            .in3(N__44414),
            .lcout(\current_shift_inst.un10_control_input_cry_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_16_7 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_17_c_RNO_LC_16_16_7  (
            .in0(N__47897),
            .in1(N__47930),
            .in2(_gnd_net_),
            .in3(N__43230),
            .lcout(\current_shift_inst.un10_control_input_cry_17_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_16_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_16_17_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_0_5_LC_16_17_0  (
            .in0(N__49877),
            .in1(N__49453),
            .in2(N__44526),
            .in3(N__44485),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_20_c_RNO_LC_16_17_1  (
            .in0(N__43233),
            .in1(N__44676),
            .in2(_gnd_net_),
            .in3(N__44654),
            .lcout(\current_shift_inst.un10_control_input_cry_20_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_22_c_RNO_LC_16_17_2  (
            .in0(N__48059),
            .in1(N__43235),
            .in2(_gnd_net_),
            .in3(N__48033),
            .lcout(\current_shift_inst.un10_control_input_cry_22_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_17_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_25_c_RNO_LC_16_17_3  (
            .in0(N__49452),
            .in1(N__44723),
            .in2(_gnd_net_),
            .in3(N__44766),
            .lcout(\current_shift_inst.un10_control_input_cry_25_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_17_4 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_21_c_RNO_LC_16_17_4  (
            .in0(N__44568),
            .in1(N__43234),
            .in2(_gnd_net_),
            .in3(N__44547),
            .lcout(\current_shift_inst.un10_control_input_cry_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_16_c_RNO_LC_16_17_5  (
            .in0(N__43231),
            .in1(N__47426),
            .in2(_gnd_net_),
            .in3(N__47393),
            .lcout(\current_shift_inst.un10_control_input_cry_16_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_19_c_RNO_LC_16_17_6  (
            .in0(N__47768),
            .in1(N__43232),
            .in2(_gnd_net_),
            .in3(N__47801),
            .lcout(\current_shift_inst.un10_control_input_cry_19_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP27A_26_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44765),
            .lcout(\current_shift_inst.un4_control_input_1_axb_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_0 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_23_c_RNO_LC_16_18_0  (
            .in0(N__43236),
            .in1(N__47965),
            .in2(_gnd_net_),
            .in3(N__48005),
            .lcout(\current_shift_inst.un10_control_input_cry_23_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_18_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_26_c_RNO_LC_16_18_1  (
            .in0(N__44320),
            .in1(N__49409),
            .in2(_gnd_net_),
            .in3(N__44292),
            .lcout(\current_shift_inst.un10_control_input_cry_26_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_18_2 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_18_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_28_c_RNO_LC_16_18_2  (
            .in0(N__49411),
            .in1(N__43406),
            .in2(_gnd_net_),
            .in3(N__43379),
            .lcout(\current_shift_inst.un10_control_input_cry_28_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_18_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_18_3 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_29_c_RNO_LC_16_18_3  (
            .in0(N__43490),
            .in1(N__49412),
            .in2(_gnd_net_),
            .in3(N__43460),
            .lcout(\current_shift_inst.un10_control_input_cry_29_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_4 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.un10_control_input_cry_27_c_RNO_LC_16_18_4  (
            .in0(N__49410),
            .in1(_gnd_net_),
            .in2(N__44390),
            .in3(N__44349),
            .lcout(\current_shift_inst.un10_control_input_cry_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIKU7A_30_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43489),
            .lcout(\current_shift_inst.un4_control_input_1_axb_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_16_18_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_16_18_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_0_16_LC_16_18_6  (
            .in0(N__49413),
            .in1(N__44461),
            .in2(N__50004),
            .in3(N__44421),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_7 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_7 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.un10_control_input_cry_24_c_RNO_LC_16_18_7  (
            .in0(N__46861),
            .in1(N__43237),
            .in2(_gnd_net_),
            .in3(N__43619),
            .lcout(\current_shift_inst.un10_control_input_cry_24_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_19_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_19_0 .LUT_INIT=16'b0010011100100111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIP3M43_LC_16_19_0  (
            .in0(N__49106),
            .in1(N__45109),
            .in2(N__48787),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.control_input_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_19_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_19_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIPTTO3_LC_16_19_1  (
            .in0(N__48157),
            .in1(N__44584),
            .in2(_gnd_net_),
            .in3(N__49104),
            .lcout(\current_shift_inst.control_input_axb_0 ),
            .ltout(\current_shift_inst.control_input_axb_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_16_19_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_16_19_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.error_control_0_LC_16_19_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \current_shift_inst.PI_CTRL.error_control_0_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43093),
            .in3(N__43085),
            .lcout(\current_shift_inst.PI_CTRL.prop_term_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52572),
            .ce(),
            .sr(N__52231));
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_19_3 .C_ON=1'b0;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_19_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un10_control_input_cry_30_c_RNI4B5I_1_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49105),
            .lcout(\current_shift_inst.N_1379_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_19_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_19_6 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNI1MCP2_LC_16_19_6  (
            .in0(N__49107),
            .in1(N__45091),
            .in2(_gnd_net_),
            .in3(N__48760),
            .lcout(\current_shift_inst.control_input_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_19_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_19_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNI983E3_LC_16_19_7  (
            .in0(N__45070),
            .in1(N__48730),
            .in2(_gnd_net_),
            .in3(N__49108),
            .lcout(\current_shift_inst.control_input_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_20_0 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_20_0 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNIHHVF3_LC_16_20_0  (
            .in0(N__48421),
            .in1(N__44779),
            .in2(_gnd_net_),
            .in3(N__49117),
            .lcout(\current_shift_inst.control_input_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_30_LC_16_20_1  (
            .in0(N__50054),
            .in1(N__49501),
            .in2(N__43501),
            .in3(N__43468),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_20_2 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_20_2 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNI1V6C3_LC_16_20_2  (
            .in0(N__48658),
            .in1(N__45010),
            .in2(_gnd_net_),
            .in3(N__49119),
            .lcout(\current_shift_inst.control_input_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_20_3 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_20_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI9HT03_LC_16_20_3  (
            .in0(N__49120),
            .in1(N__44986),
            .in2(_gnd_net_),
            .in3(N__48634),
            .lcout(\current_shift_inst.control_input_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_20_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_20_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_25_LC_16_20_4  (
            .in0(N__49499),
            .in1(N__50055),
            .in2(N__46863),
            .in3(N__43620),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_20_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_20_5 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIHQP23_LC_16_20_5  (
            .in0(N__49118),
            .in1(N__45055),
            .in2(_gnd_net_),
            .in3(N__48709),
            .lcout(\current_shift_inst.control_input_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_20_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_20_6 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI9PFN3_LC_16_20_6  (
            .in0(N__48799),
            .in1(N__45130),
            .in2(_gnd_net_),
            .in3(N__49121),
            .lcout(\current_shift_inst.control_input_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_20_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_29_LC_16_20_7  (
            .in0(N__50053),
            .in1(N__49500),
            .in2(N__43419),
            .in3(N__43380),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_21_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_21_0 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_0_26_LC_16_21_0  (
            .in0(N__50061),
            .in1(N__49503),
            .in2(N__44770),
            .in3(N__44731),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_21_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_21_1 .LUT_INIT=16'b0011001101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNI1UUF3_LC_16_21_1  (
            .in0(N__48919),
            .in1(N__45214),
            .in2(_gnd_net_),
            .in3(N__49165),
            .lcout(\current_shift_inst.control_input_axb_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_21_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_21_2 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMV731_0_30_LC_16_21_2  (
            .in0(N__43500),
            .in1(N__49507),
            .in2(N__50100),
            .in3(N__43467),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMV731_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_3 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_0_28_LC_16_21_3  (
            .in0(N__49506),
            .in1(N__50056),
            .in2(N__44395),
            .in3(N__44353),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIQ37A_27_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44324),
            .lcout(\current_shift_inst.un4_control_input_1_axb_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_0_27_LC_16_21_5  (
            .in0(N__49504),
            .in1(N__50062),
            .in2(N__44329),
            .in3(N__44296),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_6 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_6 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNI9GL43_LC_16_21_6  (
            .in0(N__49166),
            .in1(N__48892),
            .in2(_gnd_net_),
            .in3(N__45196),
            .lcout(\current_shift_inst.control_input_axb_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_21_7 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI5C531_0_29_LC_16_21_7  (
            .in0(N__49505),
            .in1(N__50057),
            .in2(N__43420),
            .in3(N__43381),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI5C531_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIE88N_10_LC_16_22_4  (
            .in0(N__43357),
            .in1(N__43345),
            .in2(N__43339),
            .in3(N__43324),
            .lcout(\current_shift_inst.PI_CTRL.output_unclamped_RNIE88NZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_22_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_22_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_22_5 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPR031_0_25_LC_16_22_5  (
            .in0(N__43621),
            .in1(N__50066),
            .in2(N__46867),
            .in3(N__49502),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPR031_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_17_6_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_17_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIJ53T9_7_LC_17_6_5  (
            .in0(N__43848),
            .in1(N__43597),
            .in2(_gnd_net_),
            .in3(N__50536),
            .lcout(elapsed_time_ns_1_RNIJ53T9_0_7),
            .ltout(elapsed_time_ns_1_RNIJ53T9_0_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_17_6_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_17_6_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_7_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43591),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_17_7_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_17_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_24_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43578),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_17_7_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_17_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_17_LC_17_7_1  (
            .in0(N__45330),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_17_7_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_17_7_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIU0DN9_20_LC_17_7_2  (
            .in0(N__43543),
            .in1(N__46942),
            .in2(_gnd_net_),
            .in3(N__50538),
            .lcout(elapsed_time_ns_1_RNIU0DN9_0_20),
            .ltout(elapsed_time_ns_1_RNIU0DN9_0_20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_17_7_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_17_7_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_20_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43537),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_7_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_7_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIH33T9_5_LC_17_7_4  (
            .in0(N__43525),
            .in1(N__43882),
            .in2(_gnd_net_),
            .in3(N__50537),
            .lcout(elapsed_time_ns_1_RNIH33T9_0_5),
            .ltout(elapsed_time_ns_1_RNIH33T9_0_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_17_7_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_17_7_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_5_LC_17_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43519),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_8_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNITUBN9_10_LC_17_8_0  (
            .in0(N__50532),
            .in1(N__43687),
            .in2(_gnd_net_),
            .in3(N__46180),
            .lcout(elapsed_time_ns_1_RNITUBN9_0_10),
            .ltout(elapsed_time_ns_1_RNITUBN9_0_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_17_8_1 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_17_8_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_10_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43681),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_8_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_8_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI35CN9_16_LC_17_8_2  (
            .in0(N__43657),
            .in1(_gnd_net_),
            .in2(N__50546),
            .in3(N__46264),
            .lcout(elapsed_time_ns_1_RNI35CN9_0_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_8_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIK63T9_8_LC_17_8_3  (
            .in0(N__43821),
            .in1(N__43672),
            .in2(_gnd_net_),
            .in3(N__50530),
            .lcout(elapsed_time_ns_1_RNIK63T9_0_8),
            .ltout(elapsed_time_ns_1_RNIK63T9_0_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_17_8_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_17_8_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_17_8_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_8_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43666),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_17_8_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_17_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_16_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43656),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_8_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIL73T9_9_LC_17_8_6  (
            .in0(N__50531),
            .in1(N__43642),
            .in2(_gnd_net_),
            .in3(N__46228),
            .lcout(elapsed_time_ns_1_RNIL73T9_0_9),
            .ltout(elapsed_time_ns_1_RNIL73T9_0_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_17_8_7 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_17_8_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_9_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43636),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_17_9_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_17_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_12_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43737),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_9_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_9_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI24CN9_15_LC_17_9_1  (
            .in0(N__43753),
            .in1(N__46279),
            .in2(_gnd_net_),
            .in3(N__50518),
            .lcout(elapsed_time_ns_1_RNI24CN9_0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_9_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_9_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNII43T9_6_LC_17_9_2  (
            .in0(N__50515),
            .in1(N__43783),
            .in2(_gnd_net_),
            .in3(N__43864),
            .lcout(elapsed_time_ns_1_RNII43T9_0_6),
            .ltout(elapsed_time_ns_1_RNII43T9_0_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_17_9_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_17_9_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_6_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43777),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_9_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIUVBN9_11_LC_17_9_4  (
            .in0(N__50516),
            .in1(N__43768),
            .in2(_gnd_net_),
            .in3(N__46213),
            .lcout(elapsed_time_ns_1_RNIUVBN9_0_11),
            .ltout(elapsed_time_ns_1_RNIUVBN9_0_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_17_9_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_17_9_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_11_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43762),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_17_9_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_17_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_15_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43752),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV0CN9_12_LC_17_9_7  (
            .in0(N__43738),
            .in1(N__46198),
            .in2(_gnd_net_),
            .in3(N__50517),
            .lcout(elapsed_time_ns_1_RNIV0CN9_0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_10_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_3_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__45315),
            .in2(N__45651),
            .in3(_gnd_net_),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_3 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_4_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__45624),
            .in2(N__45684),
            .in3(N__43690),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_5_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__45603),
            .in2(N__45652),
            .in3(N__43867),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_6_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__45625),
            .in2(N__45573),
            .in3(N__43852),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_7_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__45543),
            .in2(N__45604),
            .in3(N__43828),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_10_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_8_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__45519),
            .in2(N__45574),
            .in3(N__43801),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_8 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_10_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_10_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_9_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__45544),
            .in2(N__45492),
            .in3(N__43798),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_7 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_10_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_10_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_10_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__45942),
            .in2(N__45523),
            .in3(N__43795),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_9 ),
            .clk(N__52637),
            .ce(N__43972),
            .sr(N__52173));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_11_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_11_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_11_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__45493),
            .in2(N__45909),
            .in3(N__43792),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_11 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_11_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_11_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_12_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__45882),
            .in2(N__45946),
            .in3(N__43789),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_11_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_11_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_13_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__45855),
            .in2(N__45910),
            .in3(N__43786),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_11_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_11_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_14_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(N__45883),
            .in2(N__45829),
            .in3(N__43909),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_11_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_11_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_15_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(N__45798),
            .in2(N__45859),
            .in3(N__43906),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_11_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_16_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__45825),
            .in2(N__45777),
            .in3(N__43903),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_16 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_11_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_11_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_17_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__45799),
            .in2(N__45747),
            .in3(N__43900),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_15 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_11_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_11_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_18_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(N__45711),
            .in2(N__45778),
            .in3(N__43897),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_17 ),
            .clk(N__52631),
            .ce(N__43970),
            .sr(N__52175));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_12_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_12_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_19_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__46164),
            .in2(N__45751),
            .in3(N__43894),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_19 ),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_12_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_20_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__46140),
            .in2(N__45718),
            .in3(N__43891),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_12_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_12_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_21_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__46165),
            .in2(N__46119),
            .in3(N__43888),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_12_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_22_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__46141),
            .in2(N__46093),
            .in3(N__43885),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_12_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_12_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_23_LC_17_12_4  (
            .in0(_gnd_net_),
            .in1(N__46062),
            .in2(N__46120),
            .in3(N__43999),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_12_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_24_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__46089),
            .in2(N__46041),
            .in3(N__43996),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_24 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_12_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_12_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_25_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__46063),
            .in2(N__46011),
            .in3(N__43993),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_23 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_12_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_26_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__45972),
            .in2(N__46042),
            .in3(N__43990),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_25 ),
            .clk(N__52625),
            .ce(N__43963),
            .sr(N__52177));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_13_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_13_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_27_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__46392),
            .in2(N__46015),
            .in3(N__43987),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_27 ),
            .ltout(),
            .carryin(bfn_17_13_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .clk(N__52619),
            .ce(N__43971),
            .sr(N__52182));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_13_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_13_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_28_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__46362),
            .in2(N__45979),
            .in3(N__43984),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .clk(N__52619),
            .ce(N__43971),
            .sr(N__52182));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_13_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_13_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_29_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(N__46336),
            .in2(N__46396),
            .in3(N__43981),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_29 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .clk(N__52619),
            .ce(N__43971),
            .sr(N__52182));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_13_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_13_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_30_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__46312),
            .in2(N__46366),
            .in3(N__43978),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_30 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_28 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.un13_elapsed_time_ns_cry_29 ),
            .clk(N__52619),
            .ce(N__43971),
            .sr(N__52182));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_13_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_31_LC_17_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43975),
            .lcout(\delay_measurement_inst.delay_hc_timer.elapsed_time_hc_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52619),
            .ce(N__43971),
            .sr(N__52182));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_0_13_LC_17_14_0  (
            .in0(N__49352),
            .in1(N__50082),
            .in2(N__44062),
            .in3(N__44022),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIR36A_19_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47858),
            .lcout(\current_shift_inst.un4_control_input_1_axb_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_17_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_17_14_2 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_0_12_LC_17_14_2  (
            .in0(N__49351),
            .in1(N__50081),
            .in2(N__47299),
            .in3(N__47319),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_17_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_17_14_3 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_0_15_LC_17_14_3  (
            .in0(N__50083),
            .in1(N__49353),
            .in2(N__47107),
            .in3(N__47127),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_17_14_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_17_14_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_0_6_LC_17_14_4  (
            .in0(N__49349),
            .in1(N__50080),
            .in2(N__47644),
            .in3(N__47664),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_17_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_17_14_5 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_0_4_LC_17_14_5  (
            .in0(N__50078),
            .in1(N__49348),
            .in2(N__48360),
            .in3(N__48393),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_17_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_17_14_6 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_0_11_LC_17_14_6  (
            .in0(N__49350),
            .in1(N__47036),
            .in2(N__47074),
            .in3(N__50079),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_0_17_LC_17_14_7  (
            .in0(N__50084),
            .in1(N__49354),
            .in2(N__47401),
            .in3(N__47434),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_0_10_LC_17_15_0  (
            .in0(N__49333),
            .in1(N__44272),
            .in2(N__50085),
            .in3(N__44247),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI0J1D1_10_LC_17_15_1  (
            .in0(N__44271),
            .in1(N__49332),
            .in2(N__44248),
            .in3(N__49997),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI0J1D1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_31_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44226),
            .lcout(\current_shift_inst.elapsed_time_ns_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52600),
            .ce(N__44195),
            .sr(N__52193));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_15_3 .LUT_INIT=16'b1111000001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNITRK61_3_LC_17_15_3  (
            .in0(N__44148),
            .in1(N__49998),
            .in2(N__44170),
            .in3(N__49331),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNITRK61_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_15_4 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNO_LC_17_15_4  (
            .in0(N__49999),
            .in1(N__44166),
            .in2(N__49408),
            .in3(N__44147),
            .lcout(\current_shift_inst.un38_control_input_cry_2_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_15_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_RNO_LC_17_15_5  (
            .in0(N__44086),
            .in1(N__44095),
            .in2(_gnd_net_),
            .in3(N__49327),
            .lcout(\current_shift_inst.un38_control_input_cry_0_s0_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI2437_0_1_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44119),
            .lcout(\current_shift_inst.un4_control_input1_1 ),
            .ltout(\current_shift_inst.un4_control_input1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_15_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_15_7 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIP7EO_1_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(N__49326),
            .in2(N__44089),
            .in3(N__44085),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIP7EO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_17_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_17_16_0 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_0_23_LC_17_16_0  (
            .in0(N__49367),
            .in1(N__50012),
            .in2(N__48070),
            .in3(N__48032),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_16_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGCP11_13_LC_17_16_1  (
            .in0(N__50006),
            .in1(N__49364),
            .in2(N__44061),
            .in3(N__44026),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGCP11_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_16_2 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_0_22_LC_17_16_2  (
            .in0(N__49368),
            .in1(N__50007),
            .in2(N__44548),
            .in3(N__44575),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_16_3 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIGFT21_22_LC_17_16_3  (
            .in0(N__44574),
            .in1(N__44543),
            .in2(N__50086),
            .in3(N__49369),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIGFT21_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_16_4 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_0_24_LC_17_16_4  (
            .in0(N__49370),
            .in1(N__50013),
            .in2(N__48010),
            .in3(N__47960),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_16_5 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_0_18_LC_17_16_5  (
            .in0(N__50014),
            .in1(N__49366),
            .in2(N__47910),
            .in3(N__47934),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_16_6 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI34N61_5_LC_17_16_6  (
            .in0(N__49363),
            .in1(N__50005),
            .in2(N__44527),
            .in3(N__44484),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI34N61_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_17_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_17_16_7 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_0_14_LC_17_16_7  (
            .in0(N__50011),
            .in1(N__49365),
            .in2(N__47731),
            .in3(N__47694),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_17_17_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_17_17_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIPOS11_16_LC_17_17_0  (
            .in0(N__44460),
            .in1(N__49465),
            .in2(N__44425),
            .in3(N__49824),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIPOS11_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_17_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI28431_28_LC_17_17_1  (
            .in0(N__49471),
            .in1(N__44391),
            .in2(N__50000),
            .in3(N__44348),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI28431_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_17_17_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_17_17_2 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_0_20_LC_17_17_2  (
            .in0(N__47806),
            .in1(N__49817),
            .in2(N__47775),
            .in3(N__49468),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_17_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_17_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV3331_27_LC_17_17_3  (
            .in0(N__49470),
            .in1(N__44328),
            .in2(N__50003),
            .in3(N__44291),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV3331_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_17_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_17_4 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISV131_26_LC_17_17_4  (
            .in0(N__44761),
            .in1(N__49469),
            .in2(N__44730),
            .in3(N__49825),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISV131_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_17_17_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_17_17_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_0_21_LC_17_17_5  (
            .in0(N__49467),
            .in1(N__44683),
            .in2(N__50001),
            .in3(N__44655),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_17_6 .LUT_INIT=16'b1111001111110011;
    LogicCell40 \current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LN_LC_17_17_6  (
            .in0(N__50755),
            .in1(N__49472),
            .in2(N__44705),
            .in3(N__49829),
            .lcout(\current_shift_inst.un4_control_input_1_cry_29_c_RNIN5LNZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_17_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_17_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMS321_21_LC_17_17_7  (
            .in0(N__49466),
            .in1(N__44682),
            .in2(N__50002),
            .in3(N__44656),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMS321_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s0_c_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__44635),
            .in2(N__50676),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_18_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s0_c_inv_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(N__48206),
            .in2(N__44626),
            .in3(N__50749),
            .lcout(\current_shift_inst.un38_control_input_5_1 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_18_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_inv_LC_17_18_2  (
            .in0(N__50750),
            .in1(N__49680),
            .in2(N__44608),
            .in3(_gnd_net_),
            .lcout(\current_shift_inst.un38_control_input_5_2 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s0_c_RNIAOBJ1_LC_17_18_3  (
            .in0(_gnd_net_),
            .in1(N__44593),
            .in2(N__49884),
            .in3(N__44578),
            .lcout(\current_shift_inst.un38_control_input_0_s0_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s0_c_RNIE1ND1_LC_17_18_4  (
            .in0(_gnd_net_),
            .in1(N__49684),
            .in2(N__44953),
            .in3(N__44932),
            .lcout(\current_shift_inst.un38_control_input_0_s0_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s0_c_RNIIA281_LC_17_18_5  (
            .in0(_gnd_net_),
            .in1(N__44929),
            .in2(N__49885),
            .in3(N__44905),
            .lcout(\current_shift_inst.un38_control_input_0_s0_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s0_c_RNIMJDI1_LC_17_18_6  (
            .in0(_gnd_net_),
            .in1(N__49688),
            .in2(N__46753),
            .in3(N__44890),
            .lcout(\current_shift_inst.un38_control_input_0_s0_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s0_c_RNIQSOC1_LC_17_18_7  (
            .in0(_gnd_net_),
            .in1(N__49689),
            .in2(N__48286),
            .in3(N__44875),
            .lcout(\current_shift_inst.un38_control_input_0_s0_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s0_c_RNIU5471_LC_17_19_0  (
            .in0(_gnd_net_),
            .in1(N__49706),
            .in2(N__44872),
            .in3(N__44845),
            .lcout(\current_shift_inst.un38_control_input_0_s0_8 ),
            .ltout(),
            .carryin(bfn_17_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s0_c_RNIG9KN1_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__44842),
            .in2(N__49890),
            .in3(N__44821),
            .lcout(\current_shift_inst.un38_control_input_0_s0_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s0_c_RNIKIVH1_LC_17_19_2  (
            .in0(_gnd_net_),
            .in1(N__49710),
            .in2(N__44818),
            .in3(N__44791),
            .lcout(\current_shift_inst.un38_control_input_0_s0_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s0_c_RNI6ISE1_LC_17_19_3  (
            .in0(_gnd_net_),
            .in1(N__44788),
            .in2(N__49891),
            .in3(N__44773),
            .lcout(\current_shift_inst.un38_control_input_0_s0_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s0_c_RNIAR791_LC_17_19_4  (
            .in0(_gnd_net_),
            .in1(N__49714),
            .in2(N__45121),
            .in3(N__45103),
            .lcout(\current_shift_inst.un38_control_input_0_s0_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s0_c_RNIE4J31_LC_17_19_5  (
            .in0(_gnd_net_),
            .in1(N__45100),
            .in2(N__49892),
            .in3(N__45085),
            .lcout(\current_shift_inst.un38_control_input_0_s0_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s0_c_RNIIDUD1_LC_17_19_6  (
            .in0(_gnd_net_),
            .in1(N__49718),
            .in2(N__45082),
            .in3(N__45064),
            .lcout(\current_shift_inst.un38_control_input_0_s0_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s0_c_RNIMM981_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__45061),
            .in2(N__49893),
            .in3(N__45049),
            .lcout(\current_shift_inst.un38_control_input_0_s0_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s0_c_RNIQVK21_LC_17_20_0  (
            .in0(_gnd_net_),
            .in1(N__49894),
            .in2(N__45046),
            .in3(N__45025),
            .lcout(\current_shift_inst.un38_control_input_0_s0_16 ),
            .ltout(),
            .carryin(bfn_17_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s0_c_RNIU80D1_LC_17_20_1  (
            .in0(_gnd_net_),
            .in1(N__45022),
            .in2(N__50046),
            .in3(N__45004),
            .lcout(\current_shift_inst.un38_control_input_0_s0_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s0_c_RNI2IB71_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(N__49898),
            .in2(N__45001),
            .in3(N__44980),
            .lcout(\current_shift_inst.un38_control_input_0_s0_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s0_c_RNIKAOH1_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(N__44977),
            .in2(N__50047),
            .in3(N__44956),
            .lcout(\current_shift_inst.un38_control_input_0_s0_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s0_c_RNIOJ3C1_LC_17_20_4  (
            .in0(_gnd_net_),
            .in1(N__49902),
            .in2(N__45289),
            .in3(N__45262),
            .lcout(\current_shift_inst.un38_control_input_0_s0_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s0_c_RNIAVG41_LC_17_20_5  (
            .in0(_gnd_net_),
            .in1(N__45259),
            .in2(N__50048),
            .in3(N__45235),
            .lcout(\current_shift_inst.un38_control_input_0_s0_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s0_c_RNIE8SE1_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__49906),
            .in2(N__45232),
            .in3(N__45208),
            .lcout(\current_shift_inst.un38_control_input_0_s0_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_20_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_20_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s0_c_RNIIH791_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(N__45205),
            .in2(N__50049),
            .in3(N__45190),
            .lcout(\current_shift_inst.un38_control_input_0_s0_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_21_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_21_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s0_c_RNIMQI31_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(N__49910),
            .in2(N__45187),
            .in3(N__45169),
            .lcout(\current_shift_inst.un38_control_input_0_s0_24 ),
            .ltout(),
            .carryin(bfn_17_21_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_21_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s0_c_RNIQ3UD1_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__45166),
            .in2(N__50050),
            .in3(N__45151),
            .lcout(\current_shift_inst.un38_control_input_0_s0_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_21_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNIUC981_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__49914),
            .in2(N__45148),
            .in3(N__45139),
            .lcout(\current_shift_inst.un38_control_input_0_s0_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_21_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s0_c_RNI2MKI1_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(N__45136),
            .in2(N__50051),
            .in3(N__45124),
            .lcout(\current_shift_inst.un38_control_input_0_s0_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_21_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s0_c_RNI6VVC1_LC_17_21_4  (
            .in0(_gnd_net_),
            .in1(N__49918),
            .in2(N__45463),
            .in3(N__45439),
            .lcout(\current_shift_inst.un38_control_input_0_s0_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_21_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s0_c_RNIONC71_LC_17_21_5  (
            .in0(_gnd_net_),
            .in1(N__45436),
            .in2(N__50052),
            .in3(N__45421),
            .lcout(\current_shift_inst.un38_control_input_0_s0_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_21_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s0_c_RNIQ2461_LC_17_21_6  (
            .in0(_gnd_net_),
            .in1(N__49922),
            .in2(N__45418),
            .in3(N__45388),
            .lcout(\current_shift_inst.un38_control_input_0_s0_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s0 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_21_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_21_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_21_7 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s0_c_RNI5ORI1_LC_17_21_7  (
            .in0(N__45385),
            .in1(N__49195),
            .in2(N__49177),
            .in3(N__45370),
            .lcout(\current_shift_inst.control_input_axb_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_6_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_6_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_6_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI58DN9_27_LC_18_6_1  (
            .in0(N__45355),
            .in1(N__46600),
            .in2(_gnd_net_),
            .in3(N__50540),
            .lcout(elapsed_time_ns_1_RNI58DN9_0_27),
            .ltout(elapsed_time_ns_1_RNI58DN9_0_27_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_6_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_6_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_6_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_27_LC_18_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__45349),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_6_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_6_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_6_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI46CN9_17_LC_18_6_4  (
            .in0(N__50539),
            .in1(N__45331),
            .in2(_gnd_net_),
            .in3(N__46297),
            .lcout(elapsed_time_ns_1_RNI46CN9_0_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_0_LC_18_7_0  (
            .in0(N__46522),
            .in1(N__45303),
            .in2(_gnd_net_),
            .in3(N__45292),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_7_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_1_LC_18_7_1  (
            .in0(N__46461),
            .in1(N__45677),
            .in2(_gnd_net_),
            .in3(N__45655),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_1 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_0 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_2_LC_18_7_2  (
            .in0(N__46523),
            .in1(N__45644),
            .in2(_gnd_net_),
            .in3(N__45628),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_2 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_1 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_3_LC_18_7_3  (
            .in0(N__46462),
            .in1(N__45623),
            .in2(_gnd_net_),
            .in3(N__45607),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_3 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_2 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_4_LC_18_7_4  (
            .in0(N__46524),
            .in1(N__45596),
            .in2(_gnd_net_),
            .in3(N__45577),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_4 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_3 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_5_LC_18_7_5  (
            .in0(N__46463),
            .in1(N__45561),
            .in2(_gnd_net_),
            .in3(N__45547),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_5 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_4 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_6_LC_18_7_6  (
            .in0(N__46525),
            .in1(N__45542),
            .in2(_gnd_net_),
            .in3(N__45526),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_6 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_5 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_7_LC_18_7_7  (
            .in0(N__46464),
            .in1(N__45512),
            .in2(_gnd_net_),
            .in3(N__45496),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_7 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_6 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_7 ),
            .clk(N__52657),
            .ce(N__47469),
            .sr(N__52169));
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_8_LC_18_8_0  (
            .in0(N__46460),
            .in1(N__45485),
            .in2(_gnd_net_),
            .in3(N__45466),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_8_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_9_LC_18_8_1  (
            .in0(N__46508),
            .in1(N__45941),
            .in2(_gnd_net_),
            .in3(N__45913),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_9 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_8 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_10_LC_18_8_2  (
            .in0(N__46457),
            .in1(N__45902),
            .in2(_gnd_net_),
            .in3(N__45886),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_10 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_9 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_11_LC_18_8_3  (
            .in0(N__46505),
            .in1(N__45876),
            .in2(_gnd_net_),
            .in3(N__45862),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_11 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_10 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_12_LC_18_8_4  (
            .in0(N__46458),
            .in1(N__45848),
            .in2(_gnd_net_),
            .in3(N__45832),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_12 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_11 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_13_LC_18_8_5  (
            .in0(N__46506),
            .in1(N__45821),
            .in2(_gnd_net_),
            .in3(N__45802),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_13 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_12 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_14_LC_18_8_6  (
            .in0(N__46459),
            .in1(N__45797),
            .in2(_gnd_net_),
            .in3(N__45781),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_14 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_13 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_15_LC_18_8_7  (
            .in0(N__46507),
            .in1(N__45770),
            .in2(_gnd_net_),
            .in3(N__45754),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_15 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_14 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_15 ),
            .clk(N__52655),
            .ce(N__47470),
            .sr(N__52170));
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_16_LC_18_9_0  (
            .in0(N__46501),
            .in1(N__45740),
            .in2(_gnd_net_),
            .in3(N__45721),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_16 ),
            .ltout(),
            .carryin(bfn_18_9_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_17_LC_18_9_1  (
            .in0(N__46518),
            .in1(N__45710),
            .in2(_gnd_net_),
            .in3(N__45688),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_17 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_16 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_18_LC_18_9_2  (
            .in0(N__46502),
            .in1(N__46158),
            .in2(_gnd_net_),
            .in3(N__46144),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_18 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_17 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_19_LC_18_9_3  (
            .in0(N__46519),
            .in1(N__46139),
            .in2(_gnd_net_),
            .in3(N__46123),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_19 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_18 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_20_LC_18_9_4  (
            .in0(N__46503),
            .in1(N__46112),
            .in2(_gnd_net_),
            .in3(N__46096),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_20 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_19 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_21_LC_18_9_5  (
            .in0(N__46520),
            .in1(N__46085),
            .in2(_gnd_net_),
            .in3(N__46066),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_21 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_20 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_22_LC_18_9_6  (
            .in0(N__46504),
            .in1(N__46061),
            .in2(_gnd_net_),
            .in3(N__46045),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_22 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_21 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_23_LC_18_9_7  (
            .in0(N__46521),
            .in1(N__46034),
            .in2(_gnd_net_),
            .in3(N__46018),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_23 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_22 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_23 ),
            .clk(N__52649),
            .ce(N__47468),
            .sr(N__52171));
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_24_LC_18_10_0  (
            .in0(N__46465),
            .in1(N__46010),
            .in2(_gnd_net_),
            .in3(N__45982),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_24 ),
            .ltout(),
            .carryin(bfn_18_10_0_),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .clk(N__52642),
            .ce(N__47467),
            .sr(N__52172));
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_25_LC_18_10_1  (
            .in0(N__46499),
            .in1(N__45971),
            .in2(_gnd_net_),
            .in3(N__45949),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_25 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_24 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .clk(N__52642),
            .ce(N__47467),
            .sr(N__52172));
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_26_LC_18_10_2  (
            .in0(N__46466),
            .in1(N__46385),
            .in2(_gnd_net_),
            .in3(N__46369),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_26 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_25 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .clk(N__52642),
            .ce(N__47467),
            .sr(N__52172));
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_27_LC_18_10_3  (
            .in0(N__46500),
            .in1(N__46355),
            .in2(_gnd_net_),
            .in3(N__46339),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_27 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_26 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .clk(N__52642),
            .ce(N__47467),
            .sr(N__52172));
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4 .C_ON=1'b1;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_28_LC_18_10_4  (
            .in0(N__46467),
            .in1(N__46332),
            .in2(_gnd_net_),
            .in3(N__46318),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_28 ),
            .ltout(),
            .carryin(\delay_measurement_inst.delay_hc_timer.counter_cry_27 ),
            .carryout(\delay_measurement_inst.delay_hc_timer.counter_cry_28 ),
            .clk(N__52642),
            .ce(N__47467),
            .sr(N__52172));
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5 .SEQ_MODE=4'b1010;
    defparam \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.counter_29_LC_18_10_5  (
            .in0(N__46311),
            .in1(N__46468),
            .in2(_gnd_net_),
            .in3(N__46315),
            .lcout(\delay_measurement_inst.delay_hc_timer.counterZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52642),
            .ce(N__47467),
            .sr(N__52172));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_18_11_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_18_11_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI47DN9_26_LC_18_11_0  (
            .in0(N__46612),
            .in1(N__50619),
            .in2(_gnd_net_),
            .in3(N__50524),
            .lcout(elapsed_time_ns_1_RNI47DN9_0_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_18_11_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_18_11_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI62E01_15_LC_18_11_1  (
            .in0(N__46290),
            .in1(N__46275),
            .in2(N__46263),
            .in3(N__46557),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_18_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_18_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI69DN9_28_LC_18_11_2  (
            .in0(N__46246),
            .in1(N__46627),
            .in2(_gnd_net_),
            .in3(N__50525),
            .lcout(elapsed_time_ns_1_RNI69DN9_0_28),
            .ltout(elapsed_time_ns_1_RNI69DN9_0_28_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_18_11_3 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_18_11_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_28_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46240),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_18_11_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_18_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI7J461_10_LC_18_11_4  (
            .in0(N__46224),
            .in1(N__46209),
            .in2(N__46197),
            .in3(N__46176),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_18_11_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_18_11_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI4EBM1_13_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__50559),
            .in2(N__46705),
            .in3(N__49023),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_18_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_18_11_6 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI2L8F9_31_LC_18_11_6  (
            .in0(N__46698),
            .in1(N__46873),
            .in2(N__46681),
            .in3(N__46678),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3 ),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_7 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIDV2T9_1_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__46647),
            .in2(N__46666),
            .in3(N__46663),
            .lcout(elapsed_time_ns_1_RNIDV2T9_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_18_12_0 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_18_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIAAI01_25_LC_18_12_0  (
            .in0(N__46623),
            .in1(N__46611),
            .in2(N__46599),
            .in3(N__46569),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_12_1 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_12_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI57CN9_18_LC_18_12_1  (
            .in0(N__46546),
            .in1(N__46558),
            .in2(_gnd_net_),
            .in3(N__50477),
            .lcout(elapsed_time_ns_1_RNI57CN9_0_18),
            .ltout(elapsed_time_ns_1_RNI57CN9_0_18_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_18_12_2 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_18_12_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_18_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46540),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_18_12_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_18_12_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIV1DN9_21_LC_18_12_3  (
            .in0(N__46908),
            .in1(N__47605),
            .in2(_gnd_net_),
            .in3(N__50478),
            .lcout(elapsed_time_ns_1_RNIV1DN9_0_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_12_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNI76BE_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47535),
            .lcout(\delay_measurement_inst.delay_hc_timer.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_18_12_5 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_18_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI12J01_23_LC_18_12_5  (
            .in0(N__46989),
            .in1(N__46971),
            .in2(N__50592),
            .in3(N__46953),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_18_12_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_18_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIRPG01_19_LC_18_12_6  (
            .in0(N__46938),
            .in1(N__46920),
            .in2(N__46909),
            .in3(N__46737),
            .lcout(),
            .ltout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_18_12_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_18_12_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_18_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNIC8424_15_LC_18_12_7  (
            .in0(N__46894),
            .in1(N__46888),
            .in2(N__46882),
            .in3(N__46879),
            .lcout(\delay_measurement_inst.delay_hc_timer.delay_hc3lto30_i_a2_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_18_13_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_18_13_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIO17A_25_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46862),
            .lcout(\current_shift_inst.un4_control_input_1_axb_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_13_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_13_2 .LUT_INIT=16'b1000101110001011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_7_LC_18_13_2  (
            .in0(N__46771),
            .in1(N__49415),
            .in2(N__46804),
            .in3(N__50096),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI9CP61_0_7_LC_18_13_3  (
            .in0(N__49414),
            .in1(N__46803),
            .in2(N__50105),
            .in3(N__46770),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI9CP61_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_13_4 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_13_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI68CN9_19_LC_18_13_4  (
            .in0(N__46726),
            .in1(N__46738),
            .in2(_gnd_net_),
            .in3(N__50526),
            .lcout(elapsed_time_ns_1_RNI68CN9_0_19),
            .ltout(elapsed_time_ns_1_RNI68CN9_0_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_18_13_5 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_18_13_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_19_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__46720),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_18_13_6 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_18_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_21_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47604),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_18_13_7 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_18_13_7 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.running_RNIDNA11_LC_18_13_7  (
            .in0(N__47581),
            .in1(N__47539),
            .in2(_gnd_net_),
            .in3(N__47506),
            .lcout(\delay_measurement_inst.delay_hc_timer.N_166_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_18_14_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_18_14_0 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNISST11_17_LC_18_14_0  (
            .in0(N__47433),
            .in1(N__49380),
            .in2(N__47400),
            .in3(N__50075),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNISST11_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_14_1 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIEOIK_LC_18_14_1  (
            .in0(N__50269),
            .in1(N__50244),
            .in2(_gnd_net_),
            .in3(N__50300),
            .lcout(\current_shift_inst.timer_s1.N_164_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_18_14_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_18_14_2 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNID8O11_12_LC_18_14_2  (
            .in0(N__47320),
            .in1(N__50073),
            .in2(N__47298),
            .in3(N__49378),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNID8O11_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \current_shift_inst.timer_s1.running_RNIUKI8_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50243),
            .lcout(\current_shift_inst.timer_s1.running_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_18_14_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_18_14_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMKR11_15_LC_18_14_6  (
            .in0(N__47131),
            .in1(N__50074),
            .in2(N__47106),
            .in3(N__49379),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMKR11_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_14_7 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_14_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI3N2D1_11_LC_18_14_7  (
            .in0(N__49377),
            .in1(N__47070),
            .in2(N__50104),
            .in3(N__47038),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI3N2D1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_18_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.running_RNII51H_LC_18_15_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.timer_s1.running_RNII51H_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__50248),
            .in2(_gnd_net_),
            .in3(N__50302),
            .lcout(\current_shift_inst.timer_s1.N_163_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_18_15_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_18_15_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_18_15_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIFKR61_9_LC_18_15_1  (
            .in0(N__49371),
            .in1(N__48121),
            .in2(N__50091),
            .in3(N__48096),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIFKR61_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_18_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_18_15_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_18_15_2 .LUT_INIT=16'b1101000111010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJJU21_23_LC_18_15_2  (
            .in0(N__48066),
            .in1(N__49375),
            .in2(N__48037),
            .in3(N__50032),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJJU21_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_15_3 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_15_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_15_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIMNV21_24_LC_18_15_3  (
            .in0(N__49376),
            .in1(N__48006),
            .in2(N__50092),
            .in3(N__47964),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIMNV21_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_18_15_4 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_18_15_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_18_15_4 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIV0V11_18_LC_18_15_4  (
            .in0(N__47938),
            .in1(N__50037),
            .in2(N__47914),
            .in3(N__49372),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIV0V11_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_18_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_18_15_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI25021_19_LC_18_15_5  (
            .in0(N__49373),
            .in1(N__47867),
            .in2(N__50090),
            .in3(N__47829),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI25021_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_6 .LUT_INIT=16'b1010101000001111;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJO221_20_LC_18_15_6  (
            .in0(N__47802),
            .in1(N__50033),
            .in2(N__47776),
            .in3(N__49374),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJO221_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_16_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNIJGQ11_14_LC_18_16_0  (
            .in0(N__49347),
            .in1(N__47727),
            .in2(N__50089),
            .in3(N__47698),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNIJGQ11_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_18_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_18_16_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI68O61_6_LC_18_16_1  (
            .in0(N__49360),
            .in1(N__50018),
            .in2(N__47671),
            .in3(N__47640),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI68O61_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_16_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNI00M61_4_LC_18_16_2  (
            .in0(N__49346),
            .in1(N__48394),
            .in2(N__50087),
            .in3(N__48361),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNI00M61_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_4 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_RNO_LC_18_16_4  (
            .in0(N__49345),
            .in1(N__48334),
            .in2(N__48313),
            .in3(N__48213),
            .lcout(\current_shift_inst.un38_control_input_cry_1_s1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_18_16_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_18_16_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_18_16_5 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_0_8_LC_18_16_5  (
            .in0(N__49361),
            .in1(N__50019),
            .in2(N__48253),
            .in3(N__48273),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_6 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \current_shift_inst.timer_s1.elapsed_time_ns_1_RNICGQ61_8_LC_18_16_6  (
            .in0(N__48274),
            .in1(N__48249),
            .in2(N__50088),
            .in3(N__49362),
            .lcout(\current_shift_inst.elapsed_time_ns_1_RNICGQ61_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_17_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_LC_18_17_0  (
            .in0(_gnd_net_),
            .in1(N__50694),
            .in2(N__50677),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_17_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_17_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_1_s1_c_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__48205),
            .in2(N__48184),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_0_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_17_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_LC_18_17_2  (
            .in0(_gnd_net_),
            .in1(N__48175),
            .in2(N__49881),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_1_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_18_17_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_18_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_2_s1_c_RNIBQCJ1_LC_18_17_3  (
            .in0(_gnd_net_),
            .in1(N__49671),
            .in2(N__48166),
            .in3(N__48145),
            .lcout(\current_shift_inst.un38_control_input_0_s1_3 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_2_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_18_17_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_18_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_3_s1_c_RNIF3OD1_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(N__48142),
            .in2(N__49882),
            .in3(N__48124),
            .lcout(\current_shift_inst.un38_control_input_0_s1_4 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_3_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_18_17_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_18_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_4_s1_c_RNIJC381_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(N__49675),
            .in2(N__48589),
            .in3(N__48565),
            .lcout(\current_shift_inst.un38_control_input_0_s1_5 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_4_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_18_17_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_18_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_5_s1_c_RNINLEI1_LC_18_17_6  (
            .in0(_gnd_net_),
            .in1(N__48562),
            .in2(N__49883),
            .in3(N__48541),
            .lcout(\current_shift_inst.un38_control_input_0_s1_6 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_5_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_18_17_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_18_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_6_s1_c_RNIRUPC1_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__49679),
            .in2(N__48538),
            .in3(N__48517),
            .lcout(\current_shift_inst.un38_control_input_0_s1_7 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_6_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_18_18_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_18_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_7_s1_c_RNIV7571_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__49690),
            .in2(N__48514),
            .in3(N__48487),
            .lcout(\current_shift_inst.un38_control_input_0_s1_8 ),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_18_18_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_18_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_8_s1_c_RNIHBLN1_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__48484),
            .in2(N__49886),
            .in3(N__48460),
            .lcout(\current_shift_inst.un38_control_input_0_s1_9 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_8_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_18_18_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_18_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_9_s1_c_RNILK0I1_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__49694),
            .in2(N__48457),
            .in3(N__48433),
            .lcout(\current_shift_inst.un38_control_input_0_s1_10 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_9_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_18_18_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_10_s1_c_RNI7KTE1_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__48430),
            .in2(N__49887),
            .in3(N__48409),
            .lcout(\current_shift_inst.un38_control_input_0_s1_11 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_10_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_18_18_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_11_s1_c_RNIBT891_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__49698),
            .in2(N__48406),
            .in3(N__48772),
            .lcout(\current_shift_inst.un38_control_input_0_s1_12 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_11_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_18_18_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_18_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_12_s1_c_RNIF6K31_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__48769),
            .in2(N__49888),
            .in3(N__48748),
            .lcout(\current_shift_inst.un38_control_input_0_s1_13 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_12_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_18_18_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_18_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_13_s1_c_RNIJFVD1_LC_18_18_6  (
            .in0(_gnd_net_),
            .in1(N__49702),
            .in2(N__48745),
            .in3(N__48718),
            .lcout(\current_shift_inst.un38_control_input_0_s1_14 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_13_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_18_18_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_18_18_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_18_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_14_s1_c_RNINOA81_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__48715),
            .in2(N__49889),
            .in3(N__48697),
            .lcout(\current_shift_inst.un38_control_input_0_s1_15 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_14_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_15_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_18_19_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_18_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_15_s1_c_RNIR1M21_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__48694),
            .in2(N__49947),
            .in3(N__48673),
            .lcout(\current_shift_inst.un38_control_input_0_s1_16 ),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_18_19_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_16_s1_c_RNIVA1D1_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__49767),
            .in2(N__48670),
            .in3(N__48646),
            .lcout(\current_shift_inst.un38_control_input_0_s1_17 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_16_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_18_19_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_17_s1_c_RNI3KC71_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__48643),
            .in2(N__49948),
            .in3(N__48622),
            .lcout(\current_shift_inst.un38_control_input_0_s1_18 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_17_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_18_19_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_18_s1_c_RNILCPH1_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__49771),
            .in2(N__48619),
            .in3(N__48592),
            .lcout(\current_shift_inst.un38_control_input_0_s1_19 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_18_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_19_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_19_s1_c_RNIPL4C1_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__48982),
            .in2(N__49949),
            .in3(N__48958),
            .lcout(\current_shift_inst.un38_control_input_0_s1_20 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_19_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_19_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_19_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_20_s1_c_RNIB1I41_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__49775),
            .in2(N__48955),
            .in3(N__48931),
            .lcout(\current_shift_inst.un38_control_input_0_s1_21 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_20_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_19_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_19_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_21_s1_c_RNIFATE1_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__48928),
            .in2(N__49950),
            .in3(N__48907),
            .lcout(\current_shift_inst.un38_control_input_0_s1_22 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_21_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_19_7 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_19_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_22_s1_c_RNIJJ891_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__49779),
            .in2(N__48904),
            .in3(N__48880),
            .lcout(\current_shift_inst.un38_control_input_0_s1_23 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_22_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_23_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_20_0 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_23_s1_c_RNINSJ31_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__49951),
            .in2(N__48877),
            .in3(N__48853),
            .lcout(\current_shift_inst.un38_control_input_0_s1_24 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_20_1 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_24_s1_c_RNIR5VD1_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__48850),
            .in2(N__50067),
            .in3(N__48829),
            .lcout(\current_shift_inst.un38_control_input_0_s1_25 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_24_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_20_2 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s1_c_RNIVEA81_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__49955),
            .in2(N__48826),
            .in3(N__48814),
            .lcout(\current_shift_inst.un38_control_input_0_s1_26 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_25_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_20_3 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_26_s1_c_RNI3OLI1_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__48811),
            .in2(N__50068),
            .in3(N__48790),
            .lcout(\current_shift_inst.un38_control_input_0_s1_27 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_26_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_20_4 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_20_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_27_s1_c_RNI711D1_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__49959),
            .in2(N__50191),
            .in3(N__50167),
            .lcout(\current_shift_inst.un38_control_input_0_s1_28 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_27_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_20_5 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_20_5 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_20_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_28_s1_c_RNIPPD71_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__50164),
            .in2(N__50069),
            .in3(N__50143),
            .lcout(\current_shift_inst.un38_control_input_0_s1_29 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_28_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_18_20_6 .C_ON=1'b1;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_18_20_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_18_20_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \current_shift_inst.un38_control_input_cry_29_s1_c_RNIR4561_LC_18_20_6  (
            .in0(_gnd_net_),
            .in1(N__49963),
            .in2(N__50140),
            .in3(N__50116),
            .lcout(\current_shift_inst.un38_control_input_0_s1_30 ),
            .ltout(),
            .carryin(\current_shift_inst.un38_control_input_cry_29_s1 ),
            .carryout(\current_shift_inst.un38_control_input_cry_30_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_18_20_7 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_18_20_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_18_20_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \current_shift_inst.un38_control_input_cry_30_s1_c_RNIHNBG_LC_18_20_7  (
            .in0(N__49964),
            .in1(N__49495),
            .in2(_gnd_net_),
            .in3(N__49198),
            .lcout(\current_shift_inst.un38_control_input_0_s1_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_18_21_4 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_18_21_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_18_21_4 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_25_s0_c_RNI17P23_LC_18_21_4  (
            .in0(N__49189),
            .in1(N__49183),
            .in2(_gnd_net_),
            .in3(N__49173),
            .lcout(\current_shift_inst.control_input_axb_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_20_9_3 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_20_9_3 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_20_9_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI02CN9_13_LC_20_9_3  (
            .in0(N__49030),
            .in1(N__49012),
            .in2(_gnd_net_),
            .in3(N__50527),
            .lcout(elapsed_time_ns_1_RNI02CN9_0_13),
            .ltout(elapsed_time_ns_1_RNI02CN9_0_13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_20_9_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_20_9_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_20_9_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_13_LC_20_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__49006),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_20_10_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_20_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_14_LC_20_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50379),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_20_10_4 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_20_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_23_LC_20_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50574),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_20_11_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_20_11_0 .SEQ_MODE=4'b0000;
    defparam \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_20_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \phase_controller_inst1.stoper_hc.un3_target_ticks_axb_26_LC_20_11_0  (
            .in0(N__50620),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\phase_controller_inst1.stoper_hc.un3_target_ticks_axbZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_20_11_2 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_20_11_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI14DN9_23_LC_20_11_2  (
            .in0(N__50575),
            .in1(N__50596),
            .in2(_gnd_net_),
            .in3(N__50523),
            .lcout(elapsed_time_ns_1_RNI14DN9_0_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_11_6 .C_ON=1'b0;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_11_6 .SEQ_MODE=4'b0000;
    defparam \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_11_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \delay_measurement_inst.delay_hc_timer.elapsed_time_ns_1_RNI13CN9_14_LC_20_11_6  (
            .in0(N__50380),
            .in1(N__50563),
            .in2(_gnd_net_),
            .in3(N__50522),
            .lcout(elapsed_time_ns_1_RNI13CN9_0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \phase_controller_inst1.S1_LC_20_14_0 .C_ON=1'b0;
    defparam \phase_controller_inst1.S1_LC_20_14_0 .SEQ_MODE=4'b1010;
    defparam \phase_controller_inst1.S1_LC_20_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \phase_controller_inst1.S1_LC_20_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50342),
            .lcout(s1_phy_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52632),
            .ce(),
            .sr(N__52183));
    defparam \current_shift_inst.start_timer_s1_LC_20_14_1 .C_ON=1'b0;
    defparam \current_shift_inst.start_timer_s1_LC_20_14_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.start_timer_s1_LC_20_14_1 .LUT_INIT=16'b1001100111001100;
    LogicCell40 \current_shift_inst.start_timer_s1_LC_20_14_1  (
            .in0(N__50357),
            .in1(N__50266),
            .in2(_gnd_net_),
            .in3(N__50344),
            .lcout(\current_shift_inst.start_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52632),
            .ce(),
            .sr(N__52183));
    defparam \current_shift_inst.stop_timer_s1_LC_20_14_3 .C_ON=1'b0;
    defparam \current_shift_inst.stop_timer_s1_LC_20_14_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.stop_timer_s1_LC_20_14_3 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \current_shift_inst.stop_timer_s1_LC_20_14_3  (
            .in0(N__50358),
            .in1(N__50343),
            .in2(N__50301),
            .in3(N__50267),
            .lcout(\current_shift_inst.stop_timer_sZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52632),
            .ce(),
            .sr(N__52183));
    defparam \current_shift_inst.timer_s1.running_LC_20_14_5 .C_ON=1'b0;
    defparam \current_shift_inst.timer_s1.running_LC_20_14_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.timer_s1.running_LC_20_14_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \current_shift_inst.timer_s1.running_LC_20_14_5  (
            .in0(N__50296),
            .in1(N__50239),
            .in2(_gnd_net_),
            .in3(N__50268),
            .lcout(\current_shift_inst.timer_s1.runningZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52632),
            .ce(),
            .sr(N__52183));
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_20_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_20_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.prop_term_0_LC_20_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.prop_term_0_LC_20_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50217),
            .lcout(\current_shift_inst.PI_CTRL.prop_termZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52620),
            .ce(),
            .sr(N__52194));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_16_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_0_LC_20_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51667),
            .lcout(\current_shift_inst.PI_CTRL.output_unclampedZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52620),
            .ce(),
            .sr(N__52194));
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_20_18_1 .C_ON=1'b0;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_20_18_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \current_shift_inst.un38_control_input_cry_0_s1_c_inv_LC_20_18_1  (
            .in0(N__51475),
            .in1(N__50748),
            .in2(_gnd_net_),
            .in3(N__50698),
            .lcout(\current_shift_inst.un38_control_input_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_21_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_21_16_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIRUKD_6_LC_21_16_6  (
            .in0(_gnd_net_),
            .in1(N__53051),
            .in2(_gnd_net_),
            .in3(N__51704),
            .lcout(),
            .ltout(\current_shift_inst.PI_CTRL.control_out_2_i_o3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_21_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_21_16_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_5_LC_21_16_7  (
            .in0(N__52757),
            .in1(N__51903),
            .in2(N__50650),
            .in3(N__53175),
            .lcout(\current_shift_inst.PI_CTRL.N_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_22_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_22_16_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIFJHQ1_31_LC_22_16_0  (
            .in0(N__50646),
            .in1(N__52700),
            .in2(_gnd_net_),
            .in3(N__52874),
            .lcout(\current_shift_inst.PI_CTRL.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_16_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIMF421_6_LC_22_16_1  (
            .in0(N__53052),
            .in1(N__50635),
            .in2(N__51711),
            .in3(N__52770),
            .lcout(\current_shift_inst.PI_CTRL.N_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_22_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_22_16_4 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_22_16_4 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_RNO_0_4_LC_22_16_4  (
            .in0(N__50647),
            .in1(N__52876),
            .in2(N__52718),
            .in3(N__53111),
            .lcout(\current_shift_inst.PI_CTRL.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_22_16_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_22_16_7 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_22_16_7 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNIA0C12_4_LC_22_16_7  (
            .in0(N__52875),
            .in1(N__50645),
            .in2(N__53113),
            .in3(N__52701),
            .lcout(\current_shift_inst.PI_CTRL.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_17_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNISVKD_5_LC_22_17_1  (
            .in0(_gnd_net_),
            .in1(N__51890),
            .in2(_gnd_net_),
            .in3(N__53168),
            .lcout(\current_shift_inst.PI_CTRL.control_out_2_iv_i_o2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_16_1 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNI4C682_31_LC_23_16_1  (
            .in0(N__52900),
            .in1(N__53124),
            .in2(N__51958),
            .in3(N__52823),
            .lcout(\current_shift_inst.PI_CTRL.N_96 ),
            .ltout(\current_shift_inst.PI_CTRL.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_16_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_16_2 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNINBUA6_3_LC_23_16_2  (
            .in0(N__52983),
            .in1(N__51967),
            .in2(N__51961),
            .in3(N__52938),
            .lcout(\current_shift_inst.PI_CTRL.N_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_17_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.output_unclamped_RNILOKD_3_LC_23_17_1  (
            .in0(_gnd_net_),
            .in1(N__53104),
            .in2(_gnd_net_),
            .in3(N__52976),
            .lcout(\current_shift_inst.PI_CTRL.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pwm_generator_inst.un3_threshold_i_LC_24_10_5 .C_ON=1'b0;
    defparam \pwm_generator_inst.un3_threshold_i_LC_24_10_5 .SEQ_MODE=4'b0000;
    defparam \pwm_generator_inst.un3_threshold_i_LC_24_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \pwm_generator_inst.un3_threshold_i_LC_24_10_5  (
            .in0(N__51945),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\pwm_generator_inst.un3_threshold_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_15_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_15_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_9_LC_24_15_0 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_9_LC_24_15_0  (
            .in0(N__52834),
            .in1(N__52918),
            .in2(N__52728),
            .in3(N__51904),
            .lcout(pwm_duty_input_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52650),
            .ce(),
            .sr(N__52217));
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_2 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_2 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_10_LC_24_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52916),
            .lcout(pwm_duty_input_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52650),
            .ce(),
            .sr(N__52217));
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_15_5 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_15_5 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_1_LC_24_15_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_1_LC_24_15_5  (
            .in0(_gnd_net_),
            .in1(N__51769),
            .in2(_gnd_net_),
            .in3(N__53004),
            .lcout(pwm_duty_input_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52650),
            .ce(),
            .sr(N__52217));
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_15_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_15_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_2_LC_24_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_2_LC_24_15_6  (
            .in0(N__53005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51742),
            .lcout(pwm_duty_input_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52650),
            .ce(),
            .sr(N__52217));
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_15_7 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_15_7 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_6_LC_24_15_7 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_6_LC_24_15_7  (
            .in0(N__52917),
            .in1(N__52833),
            .in2(N__51715),
            .in3(N__52722),
            .lcout(pwm_duty_input_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52650),
            .ce(),
            .sr(N__52217));
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_0 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_0 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_0 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_5_LC_24_16_0  (
            .in0(N__52920),
            .in1(N__52830),
            .in2(N__53182),
            .in3(N__52726),
            .lcout(pwm_duty_input_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52643),
            .ce(),
            .sr(N__52223));
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_1 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_1 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_1 .LUT_INIT=16'b0011001100010011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_4_LC_24_16_1  (
            .in0(N__52832),
            .in1(N__53140),
            .in2(N__53131),
            .in3(N__53112),
            .lcout(pwm_duty_input_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52643),
            .ce(),
            .sr(N__52223));
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_16_3 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_16_3 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_7_LC_24_16_3 .LUT_INIT=16'b1011101100110000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_7_LC_24_16_3  (
            .in0(N__52831),
            .in1(N__52921),
            .in2(N__52729),
            .in3(N__53056),
            .lcout(pwm_duty_input_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52643),
            .ce(),
            .sr(N__52223));
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_0_LC_24_16_4  (
            .in0(N__53014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53003),
            .lcout(pwm_duty_input_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52643),
            .ce(),
            .sr(N__52223));
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_6 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_3_LC_24_16_6  (
            .in0(N__52984),
            .in1(N__52948),
            .in2(_gnd_net_),
            .in3(N__52942),
            .lcout(pwm_duty_input_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52643),
            .ce(),
            .sr(N__52223));
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_17_6 .C_ON=1'b0;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_17_6 .SEQ_MODE=4'b1010;
    defparam \current_shift_inst.PI_CTRL.control_out_8_LC_24_17_6 .LUT_INIT=16'b1101010111010000;
    LogicCell40 \current_shift_inst.PI_CTRL.control_out_8_LC_24_17_6  (
            .in0(N__52919),
            .in1(N__52829),
            .in2(N__52774),
            .in3(N__52727),
            .lcout(pwm_duty_input_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52638),
            .ce(),
            .sr(N__52232));
endmodule // MAIN
